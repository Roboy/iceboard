// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Feb 17 12:46:46 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(116[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(117[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(126[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(223[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(225[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(226[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(227[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(228[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(229[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(231[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(232[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(233[22:35])
    
    wire n41153;
    wire [12:0]current;   // verilog/TinyFPGA_B.v(235[22:29])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(263[22:33])
    wire [7:0]data;   // verilog/TinyFPGA_B.v(326[14:18])
    
    wire data_ready, sda_out, n7612, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(350[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(358[15:20])
    
    wire pwm_setpoint_23__N_215;
    wire [23:0]pwm_setpoint_23__N_191;
    
    wire n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, 
        n23, n45412;
    wire [7:0]commutation_state_7__N_216;
    
    wire commutation_state_7__N_224, n30270, n30269;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(222[11:28])
    
    wire n30268, n30267, n30266, n30265, n30264, n30263, n40820, 
        GHA_N_367, GLA_N_384, GHB_N_389, GLB_N_398, GHC_N_403, GLC_N_412, 
        dti_N_416, n30262, n30261, n30260, n30259, n30258, n30257, 
        RX_N_10, n1632;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_279;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        n41152, n1195, n40819, n30256, n41151, n1673;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(224[11:28])
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n30255, n40818, n30254, n28383, n731, n40817, n41150, 
        n41149, n41148, n35762, n7607, n15, n41147, n41146, n40816, 
        n4, n40815, n40389, n41145, n41144, n4_adj_5271, n30253, 
        n41143, n30251, n30250, n30249, n41142, n40814, n30248, 
        n30247, n30246, n30245, n41141, n30244, n22, n7608, n47555, 
        n652, n30243, n21, n20, n30242, n41140, n30241, n30240, 
        n30239, n30238, n41139, n30237, n30236, n49998, n30235, 
        n25788, n4_adj_5272, n41138;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n19, n3, n4_adj_5273, n5, n6, n7, n8, n9, n10, n11, 
        n12, n13, n14, n15_adj_5274, n16, n17, n18, n19_adj_5275, 
        n20_adj_5276, n21_adj_5277, n22_adj_5278, n23_adj_5279, n24_adj_5280, 
        n25_adj_5281, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n41137, n41136, n41135;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n122, n41134, n46564, n52665, n41133, n18_adj_5282, n40405, 
        n771, n41132, n41131, n40388, n625, n623, n622, n41130, 
        n36822, n41129, n36820, n36818, n41128, n41127, n35741, 
        n36810, n36808, n41126, n41125, n41124, n36800, n41123, 
        n45649, n41122, n41121, n41120, n41119, n41118, n41117, 
        n40404, n41116, n41115, n40489, n41114, n40488, n41331, 
        n40487, n41113, n41112, n41111, n36758, n36756, n36752, 
        n7_adj_5283, n36750, n40486, n40435, n40434, n40403, n36740, 
        n36832, n40433, n36770, n40402, n40401, n40432, n40400, 
        n40399, n40398, n40431, n36830, n36722, n40430, n40429, 
        n41110, n41109, n15_adj_5284, n14_adj_5285, n40428, n40397, 
        n41108, n41330, n4_adj_5286, n41107, n41106, n35695, n41329, 
        n44714, n41328, n41105, n41104, n41327, n41326, n41103, 
        n41102, n41325, n41324, n41323, tx_transmit_N_3513, n28407, 
        n41101, n2, n621, n28416, n41100, n15_adj_5287, n41322, 
        n41099, n41098, n41321, n41320, n41097, n41319, n41318, 
        n3303, n41317, n41316, n41096, n41315, n41314, n41313, 
        n41312, n41311, n40396, n41310, n42261, n41095, n41094, 
        n36712, n36710, n41093, n40427, n40426, n41092, n40387, 
        n41091, n41090, n41089, n41088, n52631, n41087, n42259, 
        n40425, n40395, n40485, n54, n46, n40484, n4_adj_5288, 
        n25438, n4452, n41086, n41085, n40483, n40555, n47127, 
        n36688, n40554, n40482, n40553, n40552, n40481, n40551, 
        n40775, n40480, n40774, n52596, n10_adj_5289, n25_adj_5290, 
        n24_adj_5291, n46621, n48240, n47264, n36514, n36700, n36694, 
        n405, n30234, n6_adj_5292, n28292, n36486, n40773, n40772, 
        n40771, n23_adj_5293, n22_adj_5294, n21_adj_5295, n20_adj_5296, 
        n19_adj_5297, n18_adj_5298, n17_adj_5299, n16_adj_5300, n15_adj_5301, 
        n14_adj_5302, n13_adj_5303, n12_adj_5304, n11_adj_5305, n10_adj_5306, 
        n9_adj_5307, n8_adj_5308, n7_adj_5309, n6_adj_5310, n5_adj_5311, 
        n4_adj_5312, n3_adj_5313, n7_adj_5314, n5609, n5_adj_5315, 
        n5_adj_5316, n7609, n6_adj_5317, n28264, n30753, n30752, 
        n30751, n40770, n30750, n30749, n53135, n41074, n41073, 
        n52565, n30748, n30747, n30744, n30743, n30742, n30741, 
        n63, n30740, n30739, n30738, n30737, n30736, n30735, n30734, 
        n30733, n30732, n30731, n30730, n30729, n30728, n30727, 
        n30726, n30725, n30724;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n30723, n30722, n30721, n17_adj_5318, n30719, n30718, 
        n30717, n30716, n2025, n30715, n30714, n16_adj_5319, n15_adj_5320, 
        n30713, n30712, n30711, n30710, n30709, direction_N_3907, 
        n30708, n30707, n30706, n30705, n30704, n10_adj_5321, n30703, 
        n30702, n30701, n30700, n30699, n30698, n30697, n30696, 
        n30695, n30694, n30693, n41072, n30692, n30691, n30690, 
        n30689, n30688, n30687, n30686, n30685, n30684, n30683, 
        n41071, n30682, n30681, n30680, n30679, n30678, n30677, 
        n30676, n30675, n30674, n30673, n30671, n30670, n30669, 
        n30668, n30667, n30666;
    wire [1:0]a_new_adj_5469;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5323, n30665, n41070, n41069, n1958, n41068, 
        n30664, n30663, n30662, n30661, n30660, n30659, n41067, 
        n30658, n30657, direction_N_3907_adj_5324, n30656, n30655, 
        n30654, n30653, n30652, n30651, n30650, n30649, n30648, 
        n45294, n30647, n30646, n30645, n30644, n30643, n30642, 
        n30641, n30640, n30639, n30638, n30637, n30636, n15_adj_5325, 
        n30635, n30634, n30633, n30632, n30631, n30630, n5_adj_5326, 
        n30629, n30628, n30627, n30626, n30625, n30624, n30623, 
        n30622, n30621, n30620, n30619, n30618, n30617, n30616, 
        n30615, n30614, n30613, n30612, n30611, n30610, n30609, 
        rw;
    wire [7:0]state_adj_5493;   // verilog/eeprom.v(23[11:16])
    
    wire n30608, n30607, n30606, n30605, n30604, n2956, n30603, 
        n14_adj_5327, n13_adj_5328, n30602, n30601, n30600, n30599, 
        n30598, n12_adj_5329, n11_adj_5330, n30597, n30596, n30595, 
        clk_out;
    wire [15:0]data_adj_5497;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_5499;   // verilog/tli4970.v(29[13:18])
    
    wire n15_adj_5341, n46606, n30594, n30593, n30592, n30591, n10_adj_5342, 
        n9_adj_5343, n9_adj_5344, n10_adj_5345, n11_adj_5346, n30590, 
        n30589, n30233, n30232, n30231, n30230, n30229, n30228, 
        n30227, n30226, n30225, n30224, n30223, n30222, n30221, 
        n30219, n30218, n4_adj_5347, n7610, n30588, n47917, n30587, 
        n30586, n30585, n30584, n30583, n30582, n30581, n30580, 
        n30579, n30578, n30577, n30576, n30575, n30574, n30573, 
        n30572, n30571, n30570, n30569, n30568, n30567, n30566, 
        n40479, n8_adj_5348, n4_adj_5349, n30565, n30564, n30563, 
        state_7__N_4293, n7066, n30562, n30561, n30216, n41066, 
        n30560, n30559, n30558, n30557, n30556, n30555, n30554, 
        n30553, n30552, n30551, n30550, n30549, n30548, n30547, 
        n30546, n30545, n30544, n41065, n30543, n30542, n30541, 
        n30540, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n3807, n4_adj_5350, n30539, n30538, n30537, n30536, n30535, 
        n30534, n30533, n30532, n30531, n30530, n30529, n41064, 
        n41063, n30528, n40394;
    wire [2:0]r_SM_Main_2__N_3542;
    
    wire n30527, n30526, n30525, n41062, n30523, n30522, n30521, 
        n30520, n30519, n30518, n30517, n30516, n30515, n30514, 
        n30513;
    wire [2:0]r_SM_Main_adj_5506;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5508;   // verilog/uart_tx.v(33[16:27])
    
    wire n41061;
    wire [2:0]r_SM_Main_2__N_3613;
    
    wire n30512, n30511, n30510, n30509, n30508, n30507, n41060, 
        n30505, n30504, n30503, n30502, n30500, n30499, n30498, 
        n30497, n30496, n30495, n30494, n30493, n30492;
    wire [7:0]state_adj_5517;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n30491, n30490, enable_slow_N_4190, n7227, n41059, n30489, 
        n40478, scl_enable_N_4177;
    wire [7:0]state_7__N_4087;
    
    wire n30488, n30212, n6686, n30487, n30486, n30485, n30484, 
        n30483;
    wire [7:0]state_7__N_4103;
    
    wire n40477, n40393, n30482, n30481, n30480, n30479, n30478, 
        n30477, n30476, n30475, n30474, n30473, n30472, n40424, 
        n41058, n41057, n40423, n36650, n40476, n30471, n30470, 
        n30469, n30211, n30210, n30209, n30208, n30207, n30206, 
        n30205, n30204, n30468, n7_adj_5357, n7264, n30203, n30467, 
        n30202, n30201, n30466, n6_adj_5358, n5_adj_5359, n4_adj_5360, 
        n3_adj_5361, n2_adj_5362, n30465, n30464, n30200, n30198, 
        n30197, n30189, n30186, n45170, n46559, n30174, n30173, 
        n30171, n30170, n30168, n30166, n6496, n30165, n30463, 
        n30163, n30462, n40422, n30461, n14_adj_5363, n30460, n10_adj_5364, 
        n30459, n30458, n29965, n36762, n30162, n30161, n30160, 
        n7611, n828, n829, n830, n831, n832, n833, n834, n861, 
        n896, n897, n898, n899, n900, n901, n927, n928, n929, 
        n930, n931, n932, n933, n934, n935, n936, n937, n938, 
        n939, n940, n941, n942, n943, n944, n945, n946, n947, 
        n948, n949, n950, n951, n952, n953, n954, n955, n956, 
        n957, n53023, n960, n10_adj_5365, n995, n996, n997, n998, 
        n999, n1000, n1001, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1059, n1093_adj_5366, n1094_adj_5367, 
        n1095_adj_5368, n1096_adj_5369, n1097_adj_5370, n1098_adj_5371, 
        n1099_adj_5372, n1100_adj_5373, n1101_adj_5374, n1125, n1127, 
        n1128, n1129, n1130, n1131, n1132, n1133, n1158, n21929, 
        n1193, n1194, n1195_adj_5375, n1196, n1197, n1198, n1199, 
        n1200, n1201, n1224, n1225, n1226, n1227, n1228, n1229, 
        n1230, n1231, n1232, n1233, n1257, n1292, n1293, n1294, 
        n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1323, 
        n1324, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
        n1333, n1356, n1391, n1392, n1393, n1394, n1395, n1396, 
        n1397, n1398, n1399, n1400, n1401, n1422, n1423, n1424, 
        n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
        n1433, n1455, n1490, n1491, n1492, n1493, n1494, n1495, 
        n1496, n1497, n1498, n1499, n1500, n1501, n1521, n1522, 
        n1523, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
        n1532, n1533, n1554, n1589, n1590, n1591, n1592, n1593, 
        n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631, n1632_adj_5376, n1633, n1653, 
        n40475, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n29783, 
        n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1752, 
        n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
        n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1818, 
        n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1851, 
        n46642, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
        n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
        n1901, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
        n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
        n1932, n1933, n1950, n41056, n1985, n1986, n1987, n1988, 
        n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
        n1997, n1998, n1999, n2000, n2001, n2016, n2017, n2018, 
        n2019, n2020, n2021, n2022, n2023, n2024, n2025_adj_5377, 
        n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
        n29730, n2049, n2084, n2085, n2086, n2087, n2088, n2089, 
        n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
        n2098, n2099, n2100, n2101, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2148, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
        n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
        n2199, n2200, n2201, n2214, n2215, n2216, n2217, n2218, 
        n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
        n2227, n2228, n2229, n2230, n2231, n2232, n2233, n46679, 
        n2247, n41055, n40474, n40473, n2282, n2283, n2284, n2285, 
        n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
        n40421, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
        n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
        n2328, n2329, n2330, n2331, n2332, n2333, n2346, n52531, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n29701, n2445, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n2511, n2512, n2513, n2514, n2515, 
        n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
        n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
        n2532, n2533, n2544, n28432, n2579, n2580, n2581, n2582, 
        n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
        n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
        n2599, n2600, n2601, n2610, n2611, n2612, n2613, n2614, 
        n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2643, n2678, n2679, n2680, n2681, 
        n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
        n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
        n2698, n2699, n2700, n2701, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
        n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
        n2729, n2730, n2731, n2732, n2733, n2742, n29684, n2777, 
        n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
        n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
        n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
        n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
        n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
        n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, 
        n2832, n2833, n2841, n2876, n2877, n2878, n2879, n2880, 
        n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
        n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
        n2897, n2898, n2899, n2900, n2901, n2907, n2908, n2909, 
        n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
        n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
        n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
        n2940, n41054, n2975, n2976, n2977, n2978, n2979, n2980, 
        n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
        n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
        n2997, n2998, n2999, n3000, n3001, n3006, n3007, n3008, 
        n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
        n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
        n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
        n3033, n3039, n3073, n3074, n3075, n3076, n3077, n3078, 
        n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
        n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
        n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3105, 
        n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
        n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
        n3130, n3131, n3132, n3133, n52669, n3138, n3173, n3174, 
        n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
        n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, 
        n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
        n3199, n3200, n3201, n3204, n3205, n3206, n3207, n3208, 
        n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
        n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
        n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
        n3233, n3237, n29660, n3272, n3273, n3274, n3275, n3276, 
        n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
        n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
        n3293, n3294, n3295, n3296, n3298, n3299, n3300, n3301, 
        n28440, n41259, n24_adj_5378, n47854, n62, n28290, n29618, 
        n41258, n29588, n29939, n30159, n52137, n41938, n41937, 
        n41936, n41935, n41934, n41933, n5_adj_5379, n29564, n41932, 
        n40472, n41931, n41930, n41929, n41928, n41927, n41926, 
        n41925, n49949, n41924, n41923, n41922, n41921, n41920, 
        n63_adj_5380, n41053, n41919, n41918, n41917, n52222, n41916, 
        n41915, n41914, n41913, n41912, n41911, n41910, n51120, 
        n49163, n52502, n41909, n41908, n41257, n41256, n41255, 
        n41254, n41253, n41252, n49155, n41052, n40386, n30158, 
        n49149, n49143, n47698, n49137, n45512, n49133, n41051, 
        n41050, n46298, n5_adj_5381, n30157, n30156, n30155, n30154, 
        n30153, n30152, n30151, n49119, n40471, n49115, n49111, 
        n44944, n48, n49, n50, n51, n52, n53, n54_adj_5382, 
        n55, n46297, n49099, n41251, n49093, n41250, n49087, n12_adj_5383, 
        n46644, n45186, n41249, n49081, n49075, n41248, n49071, 
        n49069, n41049, n46667, n46338, n30150, n30148, n46329, 
        n41048, n46312, n46391, n8_adj_5384, n49051, n46310, n46623, 
        n46308, n49045, n40470, n49039, n49037, n41047, n30147, 
        n45162, n30146, n30145, n30144, n30143, n30142, n30141, 
        n30140, n30139, n49031, n30138, n30137, n30136, n30135, 
        n30134, n30133, n30132, n30131, n49027, n49025, n14_adj_5385, 
        n10_adj_5386, n49003, n30282, n30281, n30280, n30279, n30278, 
        n30277, n48997, n30276, n30275, n30274, n30273, n30272, 
        n30271, n41247, n48991, n48985, n48981, n48977, n48971, 
        n48969, n52472, n48963, n28421, n48957, n9_adj_5387, n47283, 
        n2_adj_5388, n3_adj_5389, n4_adj_5390, n5_adj_5391, n6_adj_5392, 
        n7_adj_5393, n8_adj_5394, n9_adj_5395, n10_adj_5396, n11_adj_5397, 
        n12_adj_5398, n13_adj_5399, n14_adj_5400, n15_adj_5401, n16_adj_5402, 
        n17_adj_5403, n18_adj_5404, n19_adj_5405, n20_adj_5406, n21_adj_5407, 
        n22_adj_5408, n23_adj_5409, n24_adj_5410, n25_adj_5411, n26_adj_5412, 
        n27_adj_5413, n28_adj_5414, n29_adj_5415, n30_adj_5416, n31_adj_5417, 
        n32_adj_5418, n33_adj_5419, n48953, n48947, n48945, n41046, 
        n41045, n12_adj_5420, n40469, n41246, n41245, n41244, n41243, 
        n52200, n40468, n41242, n41738, n41241, n41737, n41736, 
        n41735, n41734, n41733, n41732, n41240, n41239, n48927, 
        n35840, n48921, n41715, n41714, n41713, n41712, n48915, 
        n40467, n41711, n41710, n41709, n41708, n41707, n41706, 
        n48911, n41705, n41704, n41703, n41702, n41701, n41700, 
        n41699, n48903, n41228, n40385, n41227, n41226, n41698, 
        n48899, n41697, n41696, n41695, n41694, n41693, n41225, 
        n40392, n41224, n41692, n41223, n41691, n41690, n41689, 
        n41688, n41687, n41686, n41222, n41221, n41685, n41684, 
        n41220, n6_adj_5421, n41219, n41218, n41683, n41682, n48891, 
        n41681, n41680, n41679, n41678, n48885, n41677, n41676, 
        n46291, n41217, n41216, n41675, n41674, n41215, n41673, 
        n48879, n41214, n41672, n41671, n41670, n41669, n41668, 
        n41667, n48875, n41213, n41212, n40420, n41666, n41211, 
        n41210, n41665, n41664, n41663, n41662, n41661, n41660, 
        n41659, n41209, n41658, n41208, n41657, n41656, n41655, 
        n41654, n41653, n41652, n41651, n41207, n41650, n48865, 
        n41649, n41648, n41206, n41647, n41205, n41646, n41645, 
        n41644, n41643, n41642, n41204, n41203, n41641, n41202, 
        n40419, n40727, n41640, n41639, n41638, n41637, n41636, 
        n13_adj_5422, n15_adj_5423, n17_adj_5424, n19_adj_5425, n41201, 
        n31_adj_5426, n40418, n33_adj_5427, n35, n37, n41635, n41, 
        n40417, n47, n40726, n49_adj_5428, n41200, n59, n61, n48857, 
        n48851, n48847, n46707, n48837, n28437, n48831, n52184, 
        n48821, n48815, n28444, n41634, n41633, n41632, n41631, 
        n48805, n41630, n6_adj_5429, n52445, n51113, n51112, n41199, 
        n51111, n51110, n41629, n41628, n41627, n48793, n40725, 
        n41626, n40724, n41625, n41624, n41623, n41622, n41621, 
        n40723, n41011, n41620, n48789, n41619, n41618, n51109, 
        n41617, n51108, n41616, n41615, n51107, n41614, n50109, 
        n48779, n41198, n48771, n45507, n41010, n48765, n41009, 
        n40722, n52417, n41197, n41613, n41612, n41611, n41008, 
        n46300, n51093, n48759, n8_adj_5430, n28429, n48753, n52241, 
        n28265, n10_adj_5431, n48743, n41610, n41609, n41196, n41608, 
        n41607, n41007, n41606, n41605, n41604, n41603, n48737, 
        n41602, n41601, n41006, n41600, n41599, n41598, n41597, 
        n41596, n40721, n40720, n41195, n47822, n52391, n48731, 
        n48729, n48723, n41005, n50107, n48719, n48717, n50105, 
        n41595, n41594, n41593, n41004, n40719, n40416, n52165, 
        n41592, n41591, n48701, n40718, n41590, n41589, n48697, 
        n41588, n41587, n41586, n41585, n41584, n41583, n41582, 
        n41581, n41580, n41579, n41578, n41577, n52967, n41576, 
        n41575, n41574, n41573, n41572, n41571, n41570, n41569, 
        n41568, n41567, n41566, n41565, n41564, n41563, n41562, 
        n41561, n41560, n41559, n41558, n41557, n41556, n41555, 
        n41554, n41553, n41552, n41551, n41550, n41549, n41548, 
        n41547, n41546, n41545, n41544, n41543, n41542, n41541, 
        n41540, n41539, n41538, n41537, n41536, n41535, n41534, 
        n41533, n41532, n41531, n41530, n41529, n52366, n41528, 
        n41527, n41526, n41525, n41524, n41523, n41522, n41521, 
        n41520, n41519, n41518, n41517, n41516, n41515, n41514, 
        n41513, n41512, n41511, n41510, n41509, n41508, n41507, 
        n41506, n30122, n41505, n41504, n41503, n48691, n8_adj_5432, 
        n7_adj_5433, n46584, n48685, n48675, n47285, n48665, n48659, 
        n40717, n41194, n41193, n36786, n48653, n40716, n48647, 
        n30124, n41192, n41191, n48643, n40415, n41190, n51068, 
        n48641, n40715, n52342, n36584, n40714, n28252, n28489, 
        n48627, n41189, n41188, n40384, n41187, n41186, n41185, 
        n41184, n36942, n48625, n20694, n40414, n40713, n40383, 
        n36580, n41459, n41458, n35782, n40712, n41457, n48619, 
        n41183, n41456, n48385, n28287, n48615, n41455, n41454, 
        n40711, n41182, n40413, n41453, n40710, n40412, n48607, 
        n41452, n41451, n41181, n40411, n41450, n40410, n36578, 
        n41449, n48601, n52319, n41448, n41447, n41446, n40409, 
        n41180, n41179, n41445, n41444, n41443, n41442, n48595, 
        n41178, n48589, n41441, n41440, n41439, n41438, n41177, 
        n40408, n41437, n36574, n48368, n50080, n40709, n41176, 
        n41175, n41174, n48579, n41173, n40708, n41172, n46575, 
        n46649, n41171, n48577, n41170, n48575, n41169, n41168, 
        n48573, n40391, n41167, n48571, n48567, n28484, n40407, 
        n48565, n41166, n41165, n48561, n52297, n48559, n41164, 
        n30123, n40406, n48549, n48360, n41163, n40390, n48547, 
        n48545, n48543, n48541, n40707, n41162, n48535, n46335, 
        n25701, n41161, n46638, n48529, n40382, n45602, n45666, 
        n48525, n39, n40, n47398, n52150, n41160, n48519, n48517, 
        n41159, n41158, n40706, n40705, n41157, n52704, n48505, 
        n41156, n41155, n41154, n48499, n52276, n48493, n48487, 
        n48481, n48479, n5_adj_5434, n46556;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n41584), .I0(n2927), 
            .I1(VCC_net), .CO(n41585));
    SB_LUT4 i16996_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n29618), 
            .I3(GND_net), .O(n30685));   // verilog/coms.v(127[12] 300[6])
    defparam i16996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16997_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n29618), 
            .I3(GND_net), .O(n30686));   // verilog/coms.v(127[12] 300[6])
    defparam i16997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16998_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n29618), 
            .I3(GND_net), .O(n30687));   // verilog/coms.v(127[12] 300[6])
    defparam i16998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n41583), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n41583), .I0(n2928), 
            .I1(VCC_net), .CO(n41584));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n41622), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16999_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30688));   // verilog/coms.v(127[12] 300[6])
    defparam i16999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17000_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30689));   // verilog/coms.v(127[12] 300[6])
    defparam i17000_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE dti_177 (.Q(dti), .C(CLK_c), .E(n29564), .D(dti_N_416));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n41582), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n41582), .I0(n2929), 
            .I1(GND_net), .CO(n41583));
    SB_LUT4 i17001_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30690));   // verilog/coms.v(127[12] 300[6])
    defparam i17001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17002_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30691));   // verilog/coms.v(127[12] 300[6])
    defparam i17002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17003_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30692));   // verilog/coms.v(127[12] 300[6])
    defparam i17003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17004_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30693));   // verilog/coms.v(127[12] 300[6])
    defparam i17004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17005_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30694));   // verilog/coms.v(127[12] 300[6])
    defparam i17005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17006_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30695));   // verilog/coms.v(127[12] 300[6])
    defparam i17006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17007_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30696));   // verilog/coms.v(127[12] 300[6])
    defparam i17007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17008_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30697));   // verilog/coms.v(127[12] 300[6])
    defparam i17008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17009_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30698));   // verilog/coms.v(127[12] 300[6])
    defparam i17009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17010_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30699));   // verilog/coms.v(127[12] 300[6])
    defparam i17010_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17011_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30700));   // verilog/coms.v(127[12] 300[6])
    defparam i17011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17012_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30701));   // verilog/coms.v(127[12] 300[6])
    defparam i17012_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 mux_236_i3_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 mux_236_i4_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4103[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n41581), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_24 (.CI(n40434), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n40435));
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n41581), .I0(n2930), 
            .I1(GND_net), .CO(n41582));
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i17013_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30702));   // verilog/coms.v(127[12] 300[6])
    defparam i17013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17014_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30703));   // verilog/coms.v(127[12] 300[6])
    defparam i17014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17015_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30704));   // verilog/coms.v(127[12] 300[6])
    defparam i17015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17016_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30705));   // verilog/coms.v(127[12] 300[6])
    defparam i17016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17017_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30706));   // verilog/coms.v(127[12] 300[6])
    defparam i17017_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n41622), .I0(n3016), 
            .I1(VCC_net), .CO(n41623));
    SB_LUT4 i17018_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30707));   // verilog/coms.v(127[12] 300[6])
    defparam i17018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n41580), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n41621), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n41580), .I0(n2931), 
            .I1(VCC_net), .CO(n41581));
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.GND_net(GND_net), .timer({timer}), 
            .CLK_c(CLK_c), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .neopxl_color({neopxl_color}), .VCC_net(VCC_net), .n2956(n2956), 
            .n30251(n30251), .n30250(n30250), .n30249(n30249), .n30248(n30248), 
            .n30247(n30247), .n30246(n30246), .n30245(n30245), .n30244(n30244), 
            .n30243(n30243), .n30242(n30242), .n30241(n30241), .n30240(n30240), 
            .n30239(n30239), .n30238(n30238), .n30237(n30237), .n30236(n30236), 
            .n30235(n30235), .n30234(n30234), .n30233(n30233), .n30232(n30232), 
            .n30231(n30231), .n30230(n30230), .n30229(n30229), .n30228(n30228), 
            .n30227(n30227), .n30226(n30226), .n30225(n30225), .n30224(n30224), 
            .n30223(n30223), .n30222(n30222), .n30221(n30221), .NEOPXL_c(NEOPXL_c), 
            .LED_c(LED_c), .n30122(n30122)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n41579), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n41621), .I0(n3017), 
            .I1(VCC_net), .CO(n41622));
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n41579), .I0(n2932), 
            .I1(GND_net), .CO(n41580));
    SB_CARRY add_224_8 (.CI(n40418), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n40419));
    SB_LUT4 i17019_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30708));   // verilog/coms.v(127[12] 300[6])
    defparam i17019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n41578), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17020_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30709));   // verilog/coms.v(127[12] 300[6])
    defparam i17020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i5_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i17021_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30710));   // verilog/coms.v(127[12] 300[6])
    defparam i17021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17022_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30711));   // verilog/coms.v(127[12] 300[6])
    defparam i17022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n41620), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n40417), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n41620), .I0(n3018), 
            .I1(VCC_net), .CO(n41621));
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17023_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30712));   // verilog/coms.v(127[12] 300[6])
    defparam i17023_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n41578), .I0(n2933), 
            .I1(VCC_net), .CO(n41579));
    SB_LUT4 i17024_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30713));   // verilog/coms.v(127[12] 300[6])
    defparam i17024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17025_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30714));   // verilog/coms.v(127[12] 300[6])
    defparam i17025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17026_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30715));   // verilog/coms.v(127[12] 300[6])
    defparam i17026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17027_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30716));   // verilog/coms.v(127[12] 300[6])
    defparam i17027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17028_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30717));   // verilog/coms.v(127[12] 300[6])
    defparam i17028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i6_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i7_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i8_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n41578));
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n52565), .I1(n2808), 
            .I2(VCC_net), .I3(n41577), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i17029_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30718));   // verilog/coms.v(127[12] 300[6])
    defparam i17029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n41576), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n41619), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17030_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30719));   // verilog/coms.v(127[12] 300[6])
    defparam i17030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16497_4_lut (.I0(n29684), .I1(r_Bit_Index_adj_5508[0]), .I2(n45512), 
            .I3(r_SM_Main_adj_5506[1]), .O(n30186));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16497_4_lut.LUT_INIT = 16'h4644;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n41576), .I0(n2809), 
            .I1(VCC_net), .CO(n41577));
    SB_LUT4 i17032_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30721));   // verilog/coms.v(127[12] 300[6])
    defparam i17032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n41575), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n40433), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17033_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30722));   // verilog/coms.v(127[12] 300[6])
    defparam i17033_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n41575), .I0(n2810), 
            .I1(VCC_net), .CO(n41576));
    SB_LUT4 i17034_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30723));   // verilog/coms.v(127[12] 300[6])
    defparam i17034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17035_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30724));   // verilog/coms.v(127[12] 300[6])
    defparam i17035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17036_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30725));   // verilog/coms.v(127[12] 300[6])
    defparam i17036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17037_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30726));   // verilog/coms.v(127[12] 300[6])
    defparam i17037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17038_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30727));   // verilog/coms.v(127[12] 300[6])
    defparam i17038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17039_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30728));   // verilog/coms.v(127[12] 300[6])
    defparam i17039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17040_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30729));   // verilog/coms.v(127[12] 300[6])
    defparam i17040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17041_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30730));   // verilog/coms.v(127[12] 300[6])
    defparam i17041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n41574), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i9_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i17042_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30731));   // verilog/coms.v(127[12] 300[6])
    defparam i17042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17043_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30732));   // verilog/coms.v(127[12] 300[6])
    defparam i17043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17044_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30733));   // verilog/coms.v(127[12] 300[6])
    defparam i17044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17045_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30734));   // verilog/coms.v(127[12] 300[6])
    defparam i17045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17046_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30735));   // verilog/coms.v(127[12] 300[6])
    defparam i17046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5280));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17047_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30736));   // verilog/coms.v(127[12] 300[6])
    defparam i17047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17048_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30737));   // verilog/coms.v(127[12] 300[6])
    defparam i17048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i17049_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30738));   // verilog/coms.v(127[12] 300[6])
    defparam i17049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17050_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30739));   // verilog/coms.v(127[12] 300[6])
    defparam i17050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17051_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30740));   // verilog/coms.v(127[12] 300[6])
    defparam i17051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17052_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30741));   // verilog/coms.v(127[12] 300[6])
    defparam i17052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17053_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30742));   // verilog/coms.v(127[12] 300[6])
    defparam i17053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17054_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n48368), .I3(GND_net), 
            .O(n30743));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i17054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17055_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n48368), .I3(GND_net), 
            .O(n30744));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i17055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n36514), .I1(n45666), .I2(state_adj_5493[0]), 
            .I3(read), .O(n45170));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut.LUT_INIT = 16'h8280;
    SB_LUT4 i30747_3_lut (.I0(n4_adj_5360), .I1(n7609), .I2(n46297), .I3(GND_net), 
            .O(n46310));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5279));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30825_4_lut (.I0(n7_adj_5283), .I1(state_adj_5493[0]), .I2(n6_adj_5292), 
            .I3(state_adj_5517[0]), .O(n46391));
    defparam i30825_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_3_lut (.I0(state_adj_5493[1]), .I1(read), .I2(n45666), 
            .I3(GND_net), .O(n12_adj_5383));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1672 (.I0(n36514), .I1(n12_adj_5383), .I2(state_adj_5493[0]), 
            .I3(n45666), .O(n45186));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1672.LUT_INIT = 16'h88a8;
    SB_LUT4 unary_minus_10_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5278));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16519_3_lut (.I0(current[5]), .I1(data_adj_5497[5]), .I2(n47264), 
            .I3(GND_net), .O(n30208));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i10_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16520_3_lut (.I0(current[4]), .I1(data_adj_5497[4]), .I2(n47264), 
            .I3(GND_net), .O(n30209));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16521_3_lut (.I0(current[3]), .I1(data_adj_5497[3]), .I2(n47264), 
            .I3(GND_net), .O(n30210));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i11_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i17058_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n48360), .I3(GND_net), 
            .O(n30747));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17059_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n48360), .I3(GND_net), 
            .O(n30748));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17060_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n48360), .I3(GND_net), 
            .O(n30749));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17061_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n48360), .I3(GND_net), 
            .O(n30750));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16522_3_lut (.I0(current[2]), .I1(data_adj_5497[2]), .I2(n47264), 
            .I3(GND_net), .O(n30211));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17062_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n48360), .I3(GND_net), 
            .O(n30751));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17063_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n48360), .I3(GND_net), 
            .O(n30752));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i12_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16523_3_lut (.I0(current[1]), .I1(data_adj_5497[1]), .I2(n47264), 
            .I3(GND_net), .O(n30212));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17064_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n48360), .I3(GND_net), 
            .O(n30753));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i17064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7264), .I2(n29730), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n44714));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_238_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n7264), .I1(n21929), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n46291));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'heaee;
    SB_LUT4 i2_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(n35695), .I2(\ID_READOUT_FSM.state [1]), 
            .I3(n46291), .O(n29730));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 add_224_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n40418), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i13_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16527_3_lut (.I0(n29730), .I1(\ID_READOUT_FSM.state [0]), .I2(n7264), 
            .I3(GND_net), .O(n30216));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16527_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 mux_236_i14_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n45412));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'hd054;
    SB_LUT4 mux_236_i15_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16452_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[7]), .I2(n35840), 
            .I3(n28440), .O(n30141));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16452_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16532_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n2956), .I3(GND_net), .O(n30221));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16533_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n2956), .I3(GND_net), .O(n30222));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16534_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n2956), .I3(GND_net), .O(n30223));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16535_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n2956), .I3(GND_net), .O(n30224));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16536_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n2956), .I3(GND_net), .O(n30225));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16537_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n2956), .I3(GND_net), .O(n30226));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16538_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n2956), .I3(GND_net), .O(n30227));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16539_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n2956), .I3(GND_net), .O(n30228));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16540_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n2956), .I3(GND_net), .O(n30229));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i16_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16541_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n2956), .I3(GND_net), .O(n30230));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16542_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n2956), .I3(GND_net), .O(n30231));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i17_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16543_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n2956), .I3(GND_net), .O(n30232));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16544_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n2956), .I3(GND_net), .O(n30233));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16453_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[8]), .I2(n9_adj_5344), 
            .I3(n28432), .O(n30142));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16453_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16545_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n2956), .I3(GND_net), .O(n30234));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16546_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n2956), .I3(GND_net), .O(n30235));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i18_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16547_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n2956), .I3(GND_net), .O(n30236));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16548_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n2956), .I3(GND_net), .O(n30237));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16549_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n2956), .I3(GND_net), .O(n30238));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16549_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n41574), .I0(n2811), 
            .I1(VCC_net), .CO(n41575));
    SB_LUT4 i16550_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n2956), .I3(GND_net), .O(n30239));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16454_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[9]), .I2(n5_adj_5315), 
            .I3(n28432), .O(n30143));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16454_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16455_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[10]), .I2(n5_adj_5316), 
            .I3(n28432), .O(n30144));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16455_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16456_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[11]), .I2(n35840), 
            .I3(n28432), .O(n30145));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16456_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16457_4_lut (.I0(state_7__N_4103[3]), .I1(data[3]), .I2(n4_adj_5350), 
            .I3(n28416), .O(n30146));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16457_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16551_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n2956), .I3(GND_net), .O(n30240));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16458_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[12]), .I2(n9_adj_5344), 
            .I3(n28429), .O(n30147));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n41573), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n41573), .I0(n2812), 
            .I1(VCC_net), .CO(n41574));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n41572), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n41572), .I0(n2813), 
            .I1(VCC_net), .CO(n41573));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n41571), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n41619), .I0(n3019), 
            .I1(VCC_net), .CO(n41620));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n41618), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n41618), .I0(n3020), 
            .I1(VCC_net), .CO(n41619));
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n41617), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i19_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16459_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[15]), .I2(n35840), 
            .I3(n28429), .O(n30148));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16459_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n41571), .I0(n2814), 
            .I1(VCC_net), .CO(n41572));
    SB_LUT4 mux_238_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n41570), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16461_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5347), 
            .I3(n28484), .O(n30150));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16461_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16462_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5271), 
            .I3(n28489), .O(n30151));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16462_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n41570), .I0(n2815), 
            .I1(VCC_net), .CO(n41571));
    SB_LUT4 i16463_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5271), 
            .I3(n28484), .O(n30152));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16463_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16464_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n28489), 
            .O(n30153));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16464_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36837_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52472));
    defparam i36837_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n41569), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16465_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n28484), 
            .O(n30154));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16465_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n41569), .I0(n2816), 
            .I1(VCC_net), .CO(n41570));
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n41568), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n41568), .I0(n2817), 
            .I1(VCC_net), .CO(n41569));
    SB_LUT4 i22086_2_lut (.I0(n25788), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n35762));
    defparam i22086_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16466_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n35741), 
            .I3(n28489), .O(n30155));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16466_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n41567), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n41617), .I0(n3021), 
            .I1(VCC_net), .CO(n41618));
    SB_LUT4 mux_238_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n41567), .I0(n2818), 
            .I1(VCC_net), .CO(n41568));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n41566), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n41566), .I0(n2819), 
            .I1(VCC_net), .CO(n41567));
    SB_LUT4 encoder0_position_31__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i20_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n7066), 
            .D(n1077), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n7066), 
            .D(n1078), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16467_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n35741), 
            .I3(n28484), .O(n30156));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16467_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16468_4_lut (.I0(state_7__N_4103[3]), .I1(data[0]), .I2(n10_adj_5431), 
            .I3(n28421), .O(n30157));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16468_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_10_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5277));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16469_4_lut (.I0(state_7__N_4103[3]), .I1(data[2]), .I2(n4_adj_5350), 
            .I3(n28421), .O(n30158));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16469_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16470_4_lut (.I0(state_7__N_4103[3]), .I1(data[1]), .I2(n10_adj_5431), 
            .I3(n28416), .O(n30159));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16470_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n41565), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16471_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30160));   // verilog/coms.v(127[12] 300[6])
    defparam i16471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16472_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n29618), 
            .I3(GND_net), .O(n30161));   // verilog/coms.v(127[12] 300[6])
    defparam i16472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16473_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n29618), 
            .I3(GND_net), .O(n30162));   // verilog/coms.v(127[12] 300[6])
    defparam i16473_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n41565), .I0(n2820), 
            .I1(VCC_net), .CO(n41566));
    SB_LUT4 i16474_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n47127), .I3(GND_net), .O(n30163));   // verilog/coms.v(127[12] 300[6])
    defparam i16474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n41564), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n41564), .I0(n2821), 
            .I1(VCC_net), .CO(n41565));
    SB_LUT4 mux_236_i21_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i22_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16476_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30165));   // verilog/coms.v(127[12] 300[6])
    defparam i16476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16477_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30166));   // verilog/coms.v(127[12] 300[6])
    defparam i16477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30766_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46329));
    defparam i30766_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i34373_4_lut (.I0(n42259), .I1(n42261), .I2(n771), .I3(n3303), 
            .O(n49949));
    defparam i34373_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n25438), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(n46338), .I1(n39), .I2(n49949), .I3(n45649), 
            .O(n40));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'hcc4c;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n54), .I1(n40), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n46329), .O(n44944));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'hccdc;
    SB_LUT4 mux_238_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i23_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i24_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16552_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n2956), .I3(GND_net), .O(n30241));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16479_3_lut (.I0(current[0]), .I1(data_adj_5497[0]), .I2(n47264), 
            .I3(GND_net), .O(n30168));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(enable_slow_N_4190), .I1(data_ready), 
            .I2(state_adj_5493[1]), .I3(state_adj_5493[0]), .O(n45294));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'hccd0;
    SB_LUT4 i16481_4_lut (.I0(rw), .I1(state_adj_5493[0]), .I2(state_adj_5493[1]), 
            .I3(n5609), .O(n30170));   // verilog/eeprom.v(26[8] 58[4])
    defparam i16481_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 unary_minus_10_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5276));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16553_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n2956), .I3(GND_net), .O(n30242));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16554_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n2956), .I3(GND_net), .O(n30243));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16555_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n2956), .I3(GND_net), .O(n30244));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16482_3_lut (.I0(CS_c), .I1(state_adj_5499[0]), .I2(state_adj_5499[1]), 
            .I3(GND_net), .O(n30171));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16482_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i37086_4_lut (.I0(n15_adj_5325), .I1(clk_out), .I2(state_adj_5499[0]), 
            .I3(state_adj_5499[1]), .O(n9_adj_5387));   // verilog/tli4970.v(33[10] 66[6])
    defparam i37086_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i23133_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n36820));
    defparam i23133_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16484_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5506[1]), .I2(n20694), 
            .I3(n4_adj_5349), .O(n30173));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16484_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i16485_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4087[0]), 
            .I3(enable_slow_N_4190), .O(n30174));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16485_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i36515_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52150));
    defparam i36515_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093_adj_5366), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36530_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52165));
    defparam i36530_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(n46623), .I1(n2118), .I2(n2122), .I3(n48805), 
            .O(n47917));
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n41563), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n41563), .I0(n2822), 
            .I1(VCC_net), .CO(n41564));
    SB_LUT4 i30736_3_lut (.I0(encoder0_position[26]), .I1(n46298), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36549_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52184));
    defparam i36549_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n41562), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n41562), .I0(n2823), 
            .I1(VCC_net), .CO(n41563));
    SB_LUT4 i1_3_lut_adj_1679 (.I0(n5_adj_5326), .I1(n3_adj_5361), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n48899));
    defparam i1_3_lut_adj_1679.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n41561), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n41561), .I0(n2824), 
            .I1(VCC_net), .CO(n41562));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n41560), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n41560), .I0(n2825), 
            .I1(VCC_net), .CO(n41561));
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n41559), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n41559), .I0(n2826), 
            .I1(VCC_net), .CO(n41560));
    SB_LUT4 i30748_3_lut (.I0(encoder0_position[29]), .I1(n46310), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_23 (.CI(n40433), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n40434));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n41558), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n41616), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n41558), .I0(n2827), 
            .I1(VCC_net), .CO(n41559));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n41557), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5358), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36565_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52200));
    defparam i36565_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n7066), 
            .D(n1079), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n41557), .I0(n2828), 
            .I1(VCC_net), .CO(n41558));
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n41556), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n41556), .I0(n2829), 
            .I1(GND_net), .CO(n41557));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n41555), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n41555), .I0(n2830), 
            .I1(GND_net), .CO(n41556));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n41554), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n41554), .I0(n2831), 
            .I1(VCC_net), .CO(n41555));
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n41553), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5359), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n405));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36587_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52222));
    defparam i36587_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5360), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n41553), .I0(n2832), 
            .I1(GND_net), .CO(n41554));
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n41552), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17), 
            .I3(n40474), .O(pwm_setpoint_23__N_191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n41552), .I0(n2833), 
            .I1(VCC_net), .CO(n41553));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n41552));
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n52531), .I1(n2709), 
            .I2(VCC_net), .I3(n41551), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5361), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n2117), .I1(n2119), .I2(n2120), .I3(n48601), 
            .O(n48607));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n41550), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n41550), .I0(n2710), 
            .I1(VCC_net), .CO(n41551));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n41549), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n41549), .I0(n2711), 
            .I1(VCC_net), .CO(n41550));
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n7066), 
            .D(n1080), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16556_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n2956), .I3(GND_net), .O(n30245));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16557_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n2956), .I3(GND_net), .O(n30246));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16557_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n7066), 
            .D(n1081), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n41548), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n41548), .I0(n2712), 
            .I1(VCC_net), .CO(n41549));
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n41547), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n41547), .I0(n2713), 
            .I1(VCC_net), .CO(n41548));
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n41546), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n41546), .I0(n2714), 
            .I1(VCC_net), .CO(n41547));
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n41616), .I0(n3022), 
            .I1(VCC_net), .CO(n41617));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n41615), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n41545), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5330), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n41545), .I0(n2715), 
            .I1(VCC_net), .CO(n41546));
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n41544), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n41544), .I0(n2716), 
            .I1(VCC_net), .CO(n41545));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n41543), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n41543), .I0(n2717), 
            .I1(VCC_net), .CO(n41544));
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n41615), .I0(n3023), 
            .I1(VCC_net), .CO(n41616));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n41542), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n41542), .I0(n2718), 
            .I1(VCC_net), .CO(n41543));
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n41541), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n41541), .I0(n2719), 
            .I1(VCC_net), .CO(n41542));
    SB_LUT4 i4829_2_lut (.I0(n2_adj_5362), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4829_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36606_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52241));
    defparam i36606_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16558_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n2956), .I3(GND_net), .O(n30247));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16559_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n2956), .I3(GND_net), .O(n30248));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16560_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n2956), .I3(GND_net), .O(n30249));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16561_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n2956), .I3(GND_net), .O(n30250));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n41614), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n41614), .I0(n3024), 
            .I1(VCC_net), .CO(n41615));
    SB_LUT4 encoder0_position_31__I_0_i777_rep_44_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i777_rep_44_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16562_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n2956), .I3(GND_net), .O(n30251));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n41540), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n41540), .I0(n2720), 
            .I1(VCC_net), .CO(n41541));
    SB_CARRY add_224_7 (.CI(n40417), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n40418));
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n41613), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n41539), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n41539), .I0(n2721), 
            .I1(VCC_net), .CO(n41540));
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n41613), .I0(n3025), 
            .I1(VCC_net), .CO(n41614));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n41538), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n41538), .I0(n2722), 
            .I1(VCC_net), .CO(n41539));
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n41537), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_10 (.CI(n40474), .I0(GND_net), .I1(n17), 
            .CO(n40475));
    SB_LUT4 add_224_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n40416), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n41537), .I0(n2723), 
            .I1(VCC_net), .CO(n41538));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n41536), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n40432), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n41536), .I0(n2724), 
            .I1(VCC_net), .CO(n41537));
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n41535), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n41535), .I0(n2725), 
            .I1(VCC_net), .CO(n41536));
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n41534), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n41534), .I0(n2726), 
            .I1(VCC_net), .CO(n41535));
    SB_LUT4 encoder0_position_31__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025_adj_5377));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n41533), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n41533), .I0(n2727), 
            .I1(VCC_net), .CO(n41534));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n41532), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n41532), .I0(n2728), 
            .I1(VCC_net), .CO(n41533));
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n41531), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint__i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_191[0]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_i1380_3_lut (.I0(n2025_adj_5377), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n41612), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n41531), .I0(n2729), 
            .I1(GND_net), .CO(n41532));
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n41612), .I0(n3026), 
            .I1(VCC_net), .CO(n41613));
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n41611), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n41530), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n41530), .I0(n2730), 
            .I1(GND_net), .CO(n41531));
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n41529), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n41529), .I0(n2731), 
            .I1(VCC_net), .CO(n41530));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n41528), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n41528), .I0(n2732), 
            .I1(GND_net), .CO(n41529));
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n41527), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_22 (.CI(n40432), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n40433));
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n41527), .I0(n2733), 
            .I1(VCC_net), .CO(n41528));
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n41527));
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n41611), .I0(n3027), 
            .I1(VCC_net), .CO(n41612));
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n7066), 
            .D(n1105), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n52502), .I1(n2610), 
            .I2(VCC_net), .I3(n41526), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n41525), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n41525), .I0(n2611), 
            .I1(VCC_net), .CO(n41526));
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n7066), 
            .D(n1082), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n41524), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n41524), .I0(n2612), 
            .I1(VCC_net), .CO(n41525));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n41523), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n41523), .I0(n2613), 
            .I1(VCC_net), .CO(n41524));
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n41522), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n7066), 
            .D(n1106), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n41522), .I0(n2614), 
            .I1(VCC_net), .CO(n41523));
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n41521), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n41521), .I0(n2615), 
            .I1(VCC_net), .CO(n41522));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n7066), 
            .D(n1108), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 unary_minus_10_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n40473), .O(pwm_setpoint_23__N_191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n41520), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n41520), .I0(n2616), 
            .I1(VCC_net), .CO(n41521));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n41519), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n41519), .I0(n2617), 
            .I1(VCC_net), .CO(n41520));
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n41518), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n41610), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n41518), .I0(n2618), 
            .I1(VCC_net), .CO(n41519));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n41517), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n5_adj_5381), .I1(n122), .I2(n3807), 
            .I3(n63_adj_5380), .O(n6_adj_5429));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'heaaa;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n41517), .I0(n2619), 
            .I1(VCC_net), .CO(n41518));
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n7066), 
            .D(n1083), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n41516), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n41516), .I0(n2620), 
            .I1(VCC_net), .CO(n41517));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n41515), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n41610), .I0(n3028), 
            .I1(VCC_net), .CO(n41611));
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n41515), .I0(n2621), 
            .I1(VCC_net), .CO(n41516));
    SB_LUT4 i3_4_lut (.I0(n53135), .I1(n6_adj_5429), .I2(n46), .I3(n4452), 
            .O(n8_adj_5430));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hcfce;
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n41514), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n41514), .I0(n2622), 
            .I1(VCC_net), .CO(n41515));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n41513), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n41513), .I0(n2623), 
            .I1(VCC_net), .CO(n41514));
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n41512), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n41512), .I0(n2624), 
            .I1(VCC_net), .CO(n41513));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n41511), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n41609), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n41511), .I0(n2625), 
            .I1(VCC_net), .CO(n41512));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n41510), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n41510), .I0(n2626), 
            .I1(VCC_net), .CO(n41511));
    SB_LUT4 i36641_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52276));
    defparam i36641_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8_adj_5430), .I2(n63), .I3(n5_adj_5434), 
            .O(n52967));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n41509), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_9 (.CI(n40473), .I0(GND_net), .I1(n18), 
            .CO(n40474));
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n41509), .I0(n2627), 
            .I1(VCC_net), .CO(n41510));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n41508), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n41508), .I0(n2628), 
            .I1(VCC_net), .CO(n41509));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n41507), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n41507), .I0(n2629), 
            .I1(GND_net), .CO(n41508));
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n41609), .I0(n3029), 
            .I1(GND_net), .CO(n41610));
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n41506), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n41506), .I0(n2630), 
            .I1(GND_net), .CO(n41507));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n41505), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n41505), .I0(n2631), 
            .I1(VCC_net), .CO(n41506));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n41504), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n41504), .I0(n2632), 
            .I1(GND_net), .CO(n41505));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n41503), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n41503), .I0(n2633), 
            .I1(VCC_net), .CO(n41504));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n41608), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n41608), .I0(n3030), 
            .I1(GND_net), .CO(n41609));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n41607), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n41607), .I0(n3031), 
            .I1(VCC_net), .CO(n41608));
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n41606), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n41503));
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n41606), .I0(n3032), 
            .I1(GND_net), .CO(n41607));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n41605), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n41605), .I0(n3033), 
            .I1(VCC_net), .CO(n41606));
    SB_LUT4 i36961_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52596));
    defparam i36961_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5275), 
            .I3(n40472), .O(pwm_setpoint_23__N_191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36662_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52297));
    defparam i36662_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n7066), 
            .D(n1084), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 add_224_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n40431), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36684_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52319));
    defparam i36684_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5290));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5291));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n7066), 
            .D(n1085), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n41605));
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n52596), .I1(n2907), 
            .I2(VCC_net), .I3(n41604), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n40392), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n41603), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_6 (.CI(n40416), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n40417));
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n41603), .I0(n2908), 
            .I1(VCC_net), .CO(n41604));
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n41602), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n41602), .I0(n2909), 
            .I1(VCC_net), .CO(n41603));
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n7066), 
            .D(n1107), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY add_224_21 (.CI(n40431), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n40432));
    SB_LUT4 add_224_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n40430), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n40384), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_20 (.CI(n40430), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n40431));
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n41601), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n41601), .I0(n2910), 
            .I1(VCC_net), .CO(n41602));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n41600), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_13 (.CI(n40392), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n40393));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n7066), 
            .D(n1086), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i36735_4_lut (.I0(n2116), .I1(n2115), .I2(n48607), .I3(n47917), 
            .O(n2148));
    defparam i36735_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n41600), .I0(n2911), 
            .I1(VCC_net), .CO(n41601));
    SB_CARRY unary_minus_10_add_3_8 (.CI(n40472), .I0(GND_net), .I1(n19_adj_5275), 
            .CO(n40473));
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n40429), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36707_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52342));
    defparam i36707_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37030_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52665));
    defparam i37030_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n41599), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5276), 
            .I3(n40471), .O(pwm_setpoint_23__N_191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_19 (.CI(n40429), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n40430));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n41599), .I0(n2912), 
            .I1(VCC_net), .CO(n41600));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5293));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36731_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52366));
    defparam i36731_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n41598), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n7066), 
            .D(n1087), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n7066), 
            .D(n1088), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5294));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_7 (.CI(n40471), .I0(GND_net), .I1(n20_adj_5276), 
            .CO(n40472));
    SB_LUT4 add_224_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n40415), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n41598), .I0(n2913), 
            .I1(VCC_net), .CO(n41599));
    SB_LUT4 unary_minus_10_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5277), 
            .I3(n40470), .O(pwm_setpoint_23__N_191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n41597), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5295));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36756_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52391));
    defparam i36756_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5296));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n41597), .I0(n2914), 
            .I1(VCC_net), .CO(n41598));
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n7066), 
            .D(n1089), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n7066), 
            .D(n1090), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n40428), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n41596), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2187_add_4_9_lut (.I0(n51113), .I1(n35762), .I2(dti_counter[7]), 
            .I3(n41738), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n52472), .I1(n2511), 
            .I2(VCC_net), .I3(n41459), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n41458), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n41458), .I0(n2512), 
            .I1(VCC_net), .CO(n41459));
    SB_LUT4 unary_minus_10_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5275));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_6 (.CI(n40470), .I0(GND_net), .I1(n21_adj_5277), 
            .CO(n40471));
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n41457), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n41457), .I0(n2513), 
            .I1(VCC_net), .CO(n41458));
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n41456), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n41456), .I0(n2514), 
            .I1(VCC_net), .CO(n41457));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n41455), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n41455), .I0(n2515), 
            .I1(VCC_net), .CO(n41456));
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n41596), .I0(n2915), 
            .I1(VCC_net), .CO(n41597));
    SB_LUT4 add_145_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n40391), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n41454), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16564_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30253));   // verilog/coms.v(127[12] 300[6])
    defparam i16564_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n41454), .I0(n2516), 
            .I1(VCC_net), .CO(n41455));
    SB_CARRY add_224_18 (.CI(n40428), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n40429));
    SB_LUT4 i16565_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30254));   // verilog/coms.v(127[12] 300[6])
    defparam i16565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16566_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30255));   // verilog/coms.v(127[12] 300[6])
    defparam i16566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n41453), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n41453), .I0(n2517), 
            .I1(VCC_net), .CO(n41454));
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n41452), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_5 (.CI(n40415), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n40416));
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n41452), .I0(n2518), 
            .I1(VCC_net), .CO(n41453));
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n41451), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16567_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30256));   // verilog/coms.v(127[12] 300[6])
    defparam i16567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n41595), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n41451), .I0(n2519), 
            .I1(VCC_net), .CO(n41452));
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n41450), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2187_add_4_8_lut (.I0(n51112), .I1(n35762), .I2(dti_counter[6]), 
            .I3(n41737), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n41450), .I0(n2520), 
            .I1(VCC_net), .CO(n41451));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n41449), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n40427), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_12 (.CI(n40391), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n40392));
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n41449), .I0(n2521), 
            .I1(VCC_net), .CO(n41450));
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n41448), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n41595), .I0(n2916), 
            .I1(VCC_net), .CO(n41596));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n41594), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n41448), .I0(n2522), 
            .I1(VCC_net), .CO(n41449));
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n41594), .I0(n2917), 
            .I1(VCC_net), .CO(n41595));
    SB_CARRY dti_counter_2187_add_4_8 (.CI(n41737), .I0(n35762), .I1(dti_counter[6]), 
            .CO(n41738));
    SB_LUT4 add_224_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n40414), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n41447), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n41593), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n41593), .I0(n2918), 
            .I1(VCC_net), .CO(n41594));
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n41447), .I0(n2523), 
            .I1(VCC_net), .CO(n41448));
    SB_LUT4 unary_minus_10_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n41446), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n41446), .I0(n2524), 
            .I1(VCC_net), .CO(n41447));
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n41445), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(244[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36867_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52502));
    defparam i36867_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
            .E(VCC_net), .D(n30216));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 mux_238_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n41592), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2187_add_4_7_lut (.I0(n51111), .I1(n35762), .I2(dti_counter[5]), 
            .I3(n41736), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n41445), .I0(n2525), 
            .I1(VCC_net), .CO(n41446));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n41444), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n41444), .I0(n2526), 
            .I1(VCC_net), .CO(n41445));
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n41592), .I0(n2919), 
            .I1(VCC_net), .CO(n41593));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n41591), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n41443), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n41443), .I0(n2527), 
            .I1(VCC_net), .CO(n41444));
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n41442), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n41442), .I0(n2528), 
            .I1(VCC_net), .CO(n41443));
    SB_CARRY dti_counter_2187_add_4_7 (.CI(n41736), .I0(n35762), .I1(dti_counter[5]), 
            .CO(n41737));
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n41441), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n41441), .I0(n2529), 
            .I1(GND_net), .CO(n41442));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n41440), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n41440), .I0(n2530), 
            .I1(GND_net), .CO(n41441));
    SB_LUT4 unary_minus_10_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5278), 
            .I3(n40469), .O(pwm_setpoint_23__N_191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n41439), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n41439), .I0(n2531), 
            .I1(VCC_net), .CO(n41440));
    SB_LUT4 i16568_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30257));   // verilog/coms.v(127[12] 300[6])
    defparam i16568_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n41591), .I0(n2920), 
            .I1(VCC_net), .CO(n41592));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n41590), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n41438), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_4 (.CI(n40414), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n40415));
    SB_CARRY unary_minus_10_add_3_5 (.CI(n40469), .I0(GND_net), .I1(n22_adj_5278), 
            .CO(n40470));
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n41438), .I0(n2532), 
            .I1(GND_net), .CO(n41439));
    SB_CARRY add_145_5 (.CI(n40384), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n40385));
    SB_LUT4 dti_counter_2187_add_4_6_lut (.I0(n51110), .I1(n35762), .I2(dti_counter[4]), 
            .I3(n41735), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n41437), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n41437), .I0(n2533), 
            .I1(VCC_net), .CO(n41438));
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n41590), .I0(n2921), 
            .I1(VCC_net), .CO(n41591));
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2187_add_4_6 (.CI(n41735), .I0(n35762), .I1(dti_counter[4]), 
            .CO(n41736));
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n41437));
    SB_LUT4 dti_counter_2187_add_4_5_lut (.I0(n51109), .I1(n35762), .I2(dti_counter[3]), 
            .I3(n41734), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n41589), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_17 (.CI(n40427), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n40428));
    SB_LUT4 add_224_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n40426), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2187_add_4_5 (.CI(n41734), .I0(n35762), .I1(dti_counter[3]), 
            .CO(n41735));
    SB_LUT4 unary_minus_10_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n41589), .I0(n2922), 
            .I1(VCC_net), .CO(n41590));
    SB_LUT4 unary_minus_10_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5279), 
            .I3(n40468), .O(pwm_setpoint_23__N_191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4512_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(107[7:14])
    defparam i4512_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_4 (.CI(n40468), .I0(GND_net), .I1(n23_adj_5279), 
            .CO(n40469));
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n41588), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1682 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n48385));
    defparam i3_4_lut_adj_1682.LUT_INIT = 16'h0004;
    SB_LUT4 unary_minus_10_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5280), 
            .I3(n40467), .O(pwm_setpoint_23__N_191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_3 (.CI(n40467), .I0(GND_net), .I1(n24_adj_5280), 
            .CO(n40468));
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n41588), .I0(n2923), 
            .I1(VCC_net), .CO(n41589));
    SB_CARRY add_224_16 (.CI(n40426), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n40427));
    SB_LUT4 dti_counter_2187_add_4_4_lut (.I0(n51108), .I1(n35762), .I2(dti_counter[2]), 
            .I3(n41733), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n41587), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25_adj_5281), 
            .I3(VCC_net), .O(pwm_setpoint_23__N_191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16508_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5347), 
            .I3(n28489), .O(n30197));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16508_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16509_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[0]), .I2(n11_adj_5346), 
            .I3(state_7__N_4293), .O(n30198));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16509_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_10_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5274));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n48360));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i16511_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n48360), .I3(GND_net), 
            .O(n30200));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16512_3_lut (.I0(current[12]), .I1(data_adj_5497[12]), .I2(n47264), 
            .I3(GND_net), .O(n30201));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16512_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n41587), .I0(n2924), 
            .I1(VCC_net), .CO(n41588));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n41586), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16581_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30270));   // verilog/coms.v(127[12] 300[6])
    defparam i16581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16513_3_lut (.I0(current[11]), .I1(data_adj_5497[11]), .I2(n47264), 
            .I3(GND_net), .O(n30202));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16514_3_lut (.I0(current[10]), .I1(data_adj_5497[10]), .I2(n47264), 
            .I3(GND_net), .O(n30203));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16514_3_lut.LUT_INIT = 16'hacac;
    SB_DFFSR pwm_setpoint__i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_191[23]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_191[22]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY unary_minus_10_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5281), 
            .CO(n40467));
    SB_LUT4 unary_minus_10_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_224_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n40425), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n40413), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_15 (.CI(n40425), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n40426));
    SB_CARRY add_224_3 (.CI(n40413), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n40414));
    SB_LUT4 unary_minus_10_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR pwm_setpoint__i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_191[21]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_191[20]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_191[19]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY dti_counter_2187_add_4_4 (.CI(n41733), .I0(n35762), .I1(dti_counter[2]), 
            .CO(n41734));
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n41586), .I0(n2925), 
            .I1(VCC_net), .CO(n41587));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n41585), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2187_add_4_3_lut (.I0(n51107), .I1(n35762), .I2(dti_counter[1]), 
            .I3(n41732), .O(n54_adj_5382)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2187_add_4_3 (.CI(n41732), .I0(n35762), .I1(dti_counter[1]), 
            .CO(n41733));
    SB_LUT4 unary_minus_10_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n41585), .I0(n2926), 
            .I1(VCC_net), .CO(n41586));
    SB_DFFSR pwm_setpoint__i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_191[18]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 dti_counter_2187_add_4_2_lut (.I0(n51093), .I1(n1958), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2187_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_DFFSR pwm_setpoint__i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_191[17]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY dti_counter_2187_add_4_2 (.CI(VCC_net), .I0(n1958), .I1(dti_counter[0]), 
            .CO(n41732));
    SB_LUT4 add_224_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n40424), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint__i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_191[16]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_191[15]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_191[14]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n41584), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint__i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_191[13]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_191[12]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_191[11]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_191[10]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_191[9]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_191[8]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_191[7]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_191[6]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_191[5]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_191[4]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_191[3]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_191[2]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_191[1]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_CARRY add_224_14 (.CI(n40424), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n40425));
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16582_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30271));   // verilog/coms.v(127[12] 300[6])
    defparam i16582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n40419), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n7066), 
            .D(n1091), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n40820), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_224_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n40423), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2), .I3(n40727), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_279), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5313), .I3(n40726), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n40726), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5313), .CO(n40727));
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5312), .I3(n40725), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_13 (.CI(n40423), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n40424));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5327), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n40819), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i981_rep_52_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i981_rep_52_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n40422), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_279), 
            .CO(n40413));
    SB_LUT4 unary_minus_10_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR GHC_184 (.Q(GHC), .C(CLK_c), .E(n29588), .D(GHC_N_403), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632_adj_5376));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632_adj_5376), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23263_4_lut (.I0(n829), .I1(n828), .I2(n36820), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i23263_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 add_145_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n40390), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n40412), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n40819), .I0(n928), 
            .I1(VCC_net), .CO(n40820));
    SB_LUT4 encoder0_position_31__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_11 (.CI(n40421), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n40422));
    SB_LUT4 encoder0_position_31__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n40725), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5312), .CO(n40726));
    SB_LUT4 unary_minus_10_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n52445), .I1(n2412), 
            .I2(VCC_net), .I3(n41331), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n41330), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n41330), .I0(n2413), 
            .I1(VCC_net), .CO(n41331));
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n41329), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n41329), .I0(n2414), 
            .I1(VCC_net), .CO(n41330));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n41328), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n41328), .I0(n2415), 
            .I1(VCC_net), .CO(n41329));
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n41327), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n41327), .I0(n2416), 
            .I1(VCC_net), .CO(n41328));
    SB_LUT4 unary_minus_10_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5311), .I3(n40724), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n40818), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n41326), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n41326), .I0(n2417), 
            .I1(VCC_net), .CO(n41327));
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n41325), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n40724), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5311), .CO(n40725));
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n41325), .I0(n2418), 
            .I1(VCC_net), .CO(n41326));
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n41324), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n40411), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n41324), .I0(n2419), 
            .I1(VCC_net), .CO(n41325));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5310), .I3(n40723), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHB_182 (.Q(GHB), .C(CLK_c), .E(n29588), .D(GHB_N_389), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n41323), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n40818), .I0(n929), 
            .I1(GND_net), .CO(n40819));
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n41323), .I0(n2420), 
            .I1(VCC_net), .CO(n41324));
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n40817), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHA_180 (.Q(GHA), .C(CLK_c), .E(n29588), .D(GHA_N_367), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i16583_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30272));   // verilog/coms.v(127[12] 300[6])
    defparam i16583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n41322), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16584_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30273));   // verilog/coms.v(127[12] 300[6])
    defparam i16584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16585_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30274));   // verilog/coms.v(127[12] 300[6])
    defparam i16585_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n41322), .I0(n2421), 
            .I1(VCC_net), .CO(n41323));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n41321), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n40817), .I0(n930), 
            .I1(GND_net), .CO(n40818));
    SB_LUT4 i16586_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30275));   // verilog/coms.v(127[12] 300[6])
    defparam i16586_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n41321), .I0(n2422), 
            .I1(VCC_net), .CO(n41322));
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n41320), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16587_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30276));   // verilog/coms.v(127[12] 300[6])
    defparam i16587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5297));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16588_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30277));   // verilog/coms.v(127[12] 300[6])
    defparam i16588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36782_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52417));
    defparam i36782_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n40723), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5310), .CO(n40724));
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n40816), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16589_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30278));   // verilog/coms.v(127[12] 300[6])
    defparam i16589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n41320), .I0(n2423), 
            .I1(VCC_net), .CO(n41321));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n41319), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5309), .I3(n40722), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16590_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30279));   // verilog/coms.v(127[12] 300[6])
    defparam i16590_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n40722), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5309), .CO(n40723));
    SB_LUT4 i16591_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30280));   // verilog/coms.v(127[12] 300[6])
    defparam i16591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16592_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30281));   // verilog/coms.v(127[12] 300[6])
    defparam i16592_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n41319), .I0(n2424), 
            .I1(VCC_net), .CO(n41320));
    SB_LUT4 i37034_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52669));
    defparam i37034_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n41318), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16593_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30282));   // verilog/coms.v(127[12] 300[6])
    defparam i16593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37069_1_lut (.I0(n36942), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52704));
    defparam i37069_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n41318), .I0(n2425), 
            .I1(VCC_net), .CO(n41319));
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n40816), .I0(n931), 
            .I1(VCC_net), .CO(n40817));
    SB_LUT4 encoder0_position_31__I_0_i2191_3_lut (.I0(n3220), .I1(n3287), 
            .I2(n3237), .I3(GND_net), .O(n31_adj_5426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n40815), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5308), .I3(n40721), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(n3224), .I1(n31_adj_5426), .I2(n3291), 
            .I3(n3237), .O(n48543));
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n3225), .I1(n19_adj_5425), .I2(n3292), 
            .I3(n3237), .O(n48545));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n3222), .I1(n13_adj_5422), .I2(n3289), 
            .I3(n3237), .O(n48549));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n3221), .I1(n15_adj_5423), .I2(n3288), 
            .I3(n3237), .O(n48547));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'heefc;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 mux_238_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22807_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n36486));
    defparam i22807_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n41317), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n41317), .I0(n2426), 
            .I1(VCC_net), .CO(n41318));
    SB_LUT4 i23005_4_lut (.I0(n36486), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n36688));
    defparam i23005_4_lut.LUT_INIT = 16'h88a0;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n40815), .I0(n932), 
            .I1(GND_net), .CO(n40816));
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n40814), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n40721), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5308), .CO(n40722));
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33_adj_5427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n3223), .I1(n17_adj_5424), .I2(n3290), 
            .I3(n3237), .O(n48541));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2189_3_lut (.I0(n3218), .I1(n3285), 
            .I2(n3237), .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1688 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5289));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i4_4_lut_adj_1688.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095_adj_5368), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_rep_43_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n50107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i837_rep_43_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_rep_53_3_lut (.I0(n50107), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i904_rep_53_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_5357), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n4_adj_5360), .I1(n5_adj_5359), .I2(n731), 
            .I3(n6_adj_5358), .O(n5_adj_5326));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_1690 (.I0(n3_adj_5361), .I1(n2_adj_5362), .I2(n5_adj_5326), 
            .I3(GND_net), .O(n46297));
    defparam i1_3_lut_adj_1690.LUT_INIT = 16'h8080;
    SB_LUT4 i30749_3_lut (.I0(n3_adj_5361), .I1(n7608), .I2(n46297), .I3(GND_net), 
            .O(n46312));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30750_3_lut (.I0(encoder0_position[30]), .I1(n46312), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i702_rep_45_3_lut (.I0(n1027), .I1(n1094_adj_5367), 
            .I2(n1059), .I3(GND_net), .O(n50109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i702_rep_45_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5307), .I3(n40720), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16580_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30269));   // verilog/coms.v(127[12] 300[6])
    defparam i16580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n48547), .I1(n48549), .I2(n48545), 
            .I3(n48543), .O(n48559));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n40814), .I0(n933), 
            .I1(VCC_net), .CO(n40815));
    SB_CARRY add_224_12 (.CI(n40422), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n40423));
    SB_LUT4 add_224_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n40421), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n41316), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2654_25_lut (.I0(n52137), .I1(n2_adj_5388), .I2(n1059), 
            .I3(n41715), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_5289), .I2(control_mode[2]), 
            .I3(GND_net), .O(n28407));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n40720), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5307), .CO(n40721));
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n51068), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5379));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n41316), .I0(n2427), 
            .I1(VCC_net), .CO(n41317));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n41315), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n2926), .I1(n2923), .I2(n2927), .I3(n2922), 
            .O(n48717));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n48559), .I1(n35), .I2(n48541), .I3(n33_adj_5427), 
            .O(n48561));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2186_3_lut (.I0(n3215), .I1(n3282), 
            .I2(n3237), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5306), .I3(n40719), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23121_4_lut (.I0(n36688), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n36808));
    defparam i23121_4_lut.LUT_INIT = 16'heefa;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n41315), .I0(n2428), 
            .I1(VCC_net), .CO(n41316));
    SB_LUT4 i1_2_lut_adj_1694 (.I0(n28252), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5341));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_adj_1694.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n41314), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n40383), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n3216), .I1(n37), .I2(n3283), .I3(n3237), 
            .O(n48969));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n36808), .I1(n41), .I2(n48561), .I3(n5_adj_5379), 
            .O(n48565));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfefc;
    SB_LUT4 add_2654_24_lut (.I0(n52150), .I1(n2_adj_5388), .I2(n1158), 
            .I3(n41714), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n40719), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5306), .CO(n40720));
    SB_CARRY add_2654_24 (.CI(n41714), .I0(n2_adj_5388), .I1(n1158), .CO(n41715));
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n41314), .I0(n2429), 
            .I1(GND_net), .CO(n41315));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n41313), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1697 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n28407), .I3(GND_net), .O(n15_adj_5287));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i2_3_lut_adj_1697.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_238_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_224_9 (.CI(n40419), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n40420));
    SB_LUT4 add_2654_23_lut (.I0(n52165), .I1(n2_adj_5388), .I2(n1257), 
            .I3(n41713), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_23 (.CI(n41713), .I0(n2_adj_5388), .I1(n1257), .CO(n41714));
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n41313), .I0(n2430), 
            .I1(GND_net), .CO(n41314));
    SB_LUT4 encoder0_position_31__I_0_i2183_3_lut (.I0(n3212), .I1(n3279), 
            .I2(n3237), .I3(GND_net), .O(n47));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n3214), .I1(n48565), .I2(n3281), .I3(n3237), 
            .O(n48567));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'heefc;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5421), .D(commutation_state_7__N_216[0]), .S(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY add_145_32 (.CI(n40411), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n40412));
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n2925), .I1(n2928), .I2(n2920), .I3(n2924), 
            .O(n48719));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n41312), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2654_22_lut (.I0(n52184), .I1(n2_adj_5388), .I2(n1356), 
            .I3(n41712), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n41312), .I0(n2431), 
            .I1(VCC_net), .CO(n41313));
    SB_LUT4 encoder0_position_31__I_0_i2182_3_lut (.I0(n3211), .I1(n3278), 
            .I2(n3237), .I3(GND_net), .O(n49_adj_5428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n3213), .I1(n48969), .I2(n3280), .I3(n3237), 
            .O(n48971));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'heefc;
    SB_LUT4 i36160_3_lut (.I0(n2925), .I1(n2992), .I2(n2940), .I3(GND_net), 
            .O(n3024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36160_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_22 (.CI(n41712), .I0(n2_adj_5388), .I1(n1356), .CO(n41713));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n41311), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5342), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2654_21_lut (.I0(n52200), .I1(n2_adj_5388), .I2(n1455), 
            .I3(n41711), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i709_rep_56_3_lut (.I0(n935), .I1(n1101_adj_5374), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i709_rep_56_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n40814));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5305), .I3(n40718), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_21 (.CI(n41711), .I0(n2_adj_5388), .I1(n1455), .CO(n41712));
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n41311), .I0(n2432), 
            .I1(GND_net), .CO(n41312));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n41310), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n41310), .I0(n2433), 
            .I1(VCC_net), .CO(n41311));
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n40718), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5305), .CO(n40719));
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n48719), .I1(n48717), .I2(n2919), .I3(n2921), 
            .O(n48723));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i23131_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n36818));
    defparam i23131_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n2916), .I1(n2917), .I2(n48723), .I3(n2918), 
            .O(n48729));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n48729), .I1(n2929), .I2(n36818), .I3(n2930), 
            .O(n48731));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n48731), 
            .O(n48737));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n48737), 
            .O(n48743));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hfffe;
    SB_LUT4 i36966_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n48743), 
            .O(n2940));
    defparam i36966_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16579_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30268));   // verilog/coms.v(127[12] 300[6])
    defparam i16579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23), .I2(encoder0_position[31]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_20_lut (.I0(n52222), .I1(n2_adj_5388), .I2(n1554), 
            .I3(n41710), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n41310));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5304), .I3(n40717), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_20 (.CI(n41710), .I0(n2_adj_5388), .I1(n1554), .CO(n41711));
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n40717), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5304), .CO(n40718));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5303), .I3(n40716), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1044_rep_39_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1044_rep_39_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30745_3_lut (.I0(n5_adj_5359), .I1(n7610), .I2(n46297), .I3(GND_net), 
            .O(n46308));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n48971), .I1(n49_adj_5428), .I2(n48567), 
            .I3(n47), .O(n48571));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n3210), .I1(n48571), .I2(n3277), .I3(n3237), 
            .O(n48573));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n40716), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5303), .CO(n40717));
    SB_LUT4 add_2654_19_lut (.I0(n52241), .I1(n2_adj_5388), .I2(n1653), 
            .I3(n41709), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_145_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n40410), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n3209), .I1(n48573), .I2(n3276), .I3(n3237), 
            .O(n48575));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5302), .I3(n40715), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2654_19 (.CI(n41709), .I0(n2_adj_5388), .I1(n1653), .CO(n41710));
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n2225), .I1(n2228), .I2(n2226), .I3(n2224), 
            .O(n48911));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n3208), .I1(n48575), .I2(n3275), .I3(n3237), 
            .O(n48577));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n3207), .I1(n48577), .I2(n3274), .I3(n3237), 
            .O(n48579));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i37072_4_lut (.I0(n61), .I1(n49998), .I2(n59), .I3(n48579), 
            .O(n36942));
    defparam i37072_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY add_145_11 (.CI(n40390), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n40391));
    SB_LUT4 add_145_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n40389), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n40715), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5302), .CO(n40716));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5301), .I3(n40714), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n40714), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5301), .CO(n40715));
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_18_lut (.I0(n52276), .I1(n2_adj_5388), .I2(n1752), 
            .I3(n41708), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_18 (.CI(n41708), .I0(n2_adj_5388), .I1(n1752), .CO(n41709));
    SB_LUT4 i36156_3_lut (.I0(n1727), .I1(n1794), .I2(n1752), .I3(GND_net), 
            .O(n1826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_17_lut (.I0(n52297), .I1(n2_adj_5388), .I2(n1851), 
            .I3(n41707), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i769_rep_55_3_lut (.I0(n50109), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i769_rep_55_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_17 (.CI(n41707), .I0(n2_adj_5388), .I1(n1851), .CO(n41708));
    SB_CARRY add_145_4 (.CI(n40383), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n40384));
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_31 (.CI(n40410), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n40411));
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5300), .I3(n40713), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n40713), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5300), .CO(n40714));
    SB_LUT4 add_2654_16_lut (.I0(n52319), .I1(n2_adj_5388), .I2(n1950), 
            .I3(n41706), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5343), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n934));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i641_rep_46_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i641_rep_46_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100_adj_5373), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_16 (.CI(n41706), .I0(n2_adj_5388), .I1(n1950), .CO(n41707));
    SB_LUT4 add_2654_15_lut (.I0(n52342), .I1(n2_adj_5388), .I2(n2049), 
            .I3(n41705), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_15 (.CI(n41705), .I0(n2_adj_5388), .I1(n2049), .CO(n41706));
    SB_LUT4 add_2654_14_lut (.I0(n52366), .I1(n2_adj_5388), .I2(n2148), 
            .I3(n41704), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_14 (.CI(n41704), .I0(n2_adj_5388), .I1(n2148), .CO(n41705));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22), .I2(encoder0_position[31]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2654_13_lut (.I0(n52391), .I1(n2_adj_5388), .I2(n2247), 
            .I3(n41703), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_13 (.CI(n41703), .I0(n2_adj_5388), .I1(n2247), .CO(n41704));
    SB_LUT4 add_2654_12_lut (.I0(n52417), .I1(n2_adj_5388), .I2(n2346), 
            .I3(n41702), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_12 (.CI(n41702), .I0(n2_adj_5388), .I1(n2346), .CO(n41703));
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36154_3_lut (.I0(n1627), .I1(n1694), .I2(n1653), .I3(GND_net), 
            .O(n1726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i36154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5299), .I3(n40712), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_10 (.CI(n40389), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n40390));
    SB_LUT4 i30746_3_lut (.I0(encoder0_position[28]), .I1(n46308), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_145_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n40382), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5348), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n834));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23055_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n36740));
    defparam i23055_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i573_rep_47_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i573_rep_47_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099_adj_5372), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1712 (.I0(n3225), .I1(n3218), .I2(n3219), .I3(GND_net), 
            .O(n49111));
    defparam i1_3_lut_adj_1712.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_11_lut (.I0(n52445), .I1(n2_adj_5388), .I2(n2445), 
            .I3(n41701), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i23123_4_lut (.I0(n957), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n36810));
    defparam i23123_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n3216), .I1(n49111), .I2(n3220), .I3(n3221), 
            .O(n49115));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1714 (.I0(n3229), .I1(n3230), .I2(GND_net), .I3(GND_net), 
            .O(n49163));
    defparam i1_2_lut_adj_1714.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n3223), .I1(n3227), .I2(n3228), .I3(n3226), 
            .O(n49133));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n3217), .I1(n49133), .I2(n3222), .I3(n3224), 
            .O(n49137));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n3213), .I1(n3214), .I2(n3215), .I3(n49137), 
            .O(n49143));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n3209), .I1(n3210), .I2(n3211), .I3(n49143), 
            .O(n49149));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n3212), .I1(n49163), .I2(n49115), .I3(n36810), 
            .O(n49119));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n3207), .I1(n3206), .I2(n3208), .I3(n49149), 
            .O(n48240));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_CARRY add_2654_11 (.CI(n41701), .I0(n2_adj_5388), .I1(n2445), .CO(n41702));
    SB_LUT4 i37067_4_lut (.I0(n3205), .I1(n3204), .I2(n48240), .I3(n49119), 
            .O(n3237));
    defparam i37067_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2041_3_lut (.I0(n3006), .I1(n3073), 
            .I2(n3039), .I3(GND_net), .O(n3105));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_10_lut (.I0(n52472), .I1(n2_adj_5388), .I2(n2544), 
            .I3(n41700), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2042_rep_50_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2042_rep_50_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16433_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n2956), .I3(GND_net), .O(n30122));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16434_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n48368), .I3(GND_net), 
            .O(n30123));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16434_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_10 (.CI(n41700), .I0(n2_adj_5388), .I1(n2544), .CO(n41701));
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16435_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30124));   // verilog/coms.v(127[12] 300[6])
    defparam i16435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n40420), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n40712), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5299), .CO(n40713));
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i975_rep_61_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i975_rep_61_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23113_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n36800));
    defparam i23113_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1721 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n48685));
    defparam i1_2_lut_adj_1721.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n927), .I1(n48685), .I2(n928), .I3(n36800), 
            .O(n960));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfefa;
    SB_LUT4 add_2654_9_lut (.I0(n52502), .I1(n2_adj_5388), .I2(n2643), 
            .I3(n41699), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_9 (.CI(n41699), .I0(n2_adj_5388), .I1(n2643), .CO(n41700));
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_8_lut (.I0(n52531), .I1(n2_adj_5388), .I2(n2742), 
            .I3(n41698), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n40409), .O(n1080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1857_rep_16_3_lut (.I0(n2793), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n50080));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1857_rep_16_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35866_3_lut (.I0(n2924), .I1(n2991), .I2(n2940), .I3(GND_net), 
            .O(n3023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i35866_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30735_3_lut (.I0(n7_adj_5357), .I1(n7612), .I2(n46297), .I3(GND_net), 
            .O(n46298));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098_adj_5371), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16442_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[1]), .I2(n10_adj_5345), 
            .I3(n28437), .O(n30131));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16442_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16443_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[2]), .I2(n5_adj_5316), 
            .I3(n28444), .O(n30132));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16443_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5298), .I3(n40711), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i22967_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n36650));
    defparam i22967_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16444_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[3]), .I2(n35840), 
            .I3(n28444), .O(n30133));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16444_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16445_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[4]), .I2(n9_adj_5344), 
            .I3(n28440), .O(n30134));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16445_4_lut.LUT_INIT = 16'hccca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i16446_4_lut (.I0(state_7__N_4103[3]), .I1(data[7]), .I2(n35782), 
            .I3(n28416), .O(n30135));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16446_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n3124), .I1(n3122), .I2(n3121), .I3(n3128), 
            .O(n48479));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i16447_4_lut (.I0(state_7__N_4103[3]), .I1(data[6]), .I2(n35782), 
            .I3(n28421), .O(n30136));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16447_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n3118), .I1(n3120), .I2(n3119), .I3(n3127), 
            .O(n48481));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n3125), .I1(n3116), .I2(n3126), .I3(n3123), 
            .O(n47854));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 i23011_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n36694));
    defparam i23011_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n47854), .I1(n3117), .I2(n48481), .I3(n48479), 
            .O(n48487));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n3129), .I1(n36694), .I2(n3130), .I3(n3131), 
            .O(n46667));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n3114), .I1(n46667), .I2(n48487), .I3(n3115), 
            .O(n48493));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n48493), 
            .O(n48499));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n48499), 
            .O(n48505));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 i37033_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n48505), 
            .O(n3138));
    defparam i37033_4_lut.LUT_INIT = 16'h0001;
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_8 (.CI(n41698), .I0(n2_adj_5388), .I1(n2742), .CO(n41699));
    SB_LUT4 add_2654_7_lut (.I0(n52565), .I1(n2_adj_5388), .I2(n2841), 
            .I3(n41697), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_7 (.CI(n41697), .I0(n2_adj_5388), .I1(n2841), .CO(n41698));
    SB_LUT4 add_2654_6_lut (.I0(n52596), .I1(n2_adj_5388), .I2(n2940), 
            .I3(n41696), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_6 (.CI(n41696), .I0(n2_adj_5388), .I1(n2940), .CO(n41697));
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_5_lut (.I0(n52631), .I1(n2_adj_5388), .I2(n3039), 
            .I3(n41695), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_5 (.CI(n41695), .I0(n2_adj_5388), .I1(n3039), .CO(n41696));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n40711), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5298), .CO(n40712));
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2654_4_lut (.I0(n52665), .I1(n2_adj_5388), .I2(n3138), 
            .I3(n41694), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_4 (.CI(n41694), .I0(n2_adj_5388), .I1(n3138), .CO(n41695));
    SB_LUT4 add_2654_3_lut (.I0(n52669), .I1(n2_adj_5388), .I2(n3237), 
            .I3(n41693), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2654_3 (.CI(n41693), .I0(n2_adj_5388), .I1(n3237), .CO(n41694));
    SB_LUT4 add_2654_2_lut (.I0(n52704), .I1(n2_adj_5388), .I2(n36942), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2654_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2654_2 (.CI(VCC_net), .I0(n2_adj_5388), .I1(n36942), 
            .CO(n41693));
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(n52669), .I1(n3204), 
            .I2(VCC_net), .I3(n41692), .O(n49998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n41691), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n41691), .I0(n3205), 
            .I1(VCC_net), .CO(n41692));
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n41690), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n41690), .I0(n3206), 
            .I1(VCC_net), .CO(n41691));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n41689), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n41689), .I0(n3207), 
            .I1(VCC_net), .CO(n41690));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n52417), .I1(n2313), 
            .I2(VCC_net), .I3(n41259), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n41688), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n41688), .I0(n3208), 
            .I1(VCC_net), .CO(n41689));
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n41687), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n41687), .I0(n3209), 
            .I1(VCC_net), .CO(n41688));
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n41686), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n41686), .I0(n3210), 
            .I1(VCC_net), .CO(n41687));
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n41685), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n41258), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n41685), .I0(n3211), 
            .I1(VCC_net), .CO(n41686));
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n41258), .I0(n2314), 
            .I1(VCC_net), .CO(n41259));
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n41257), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n41257), .I0(n2315), 
            .I1(VCC_net), .CO(n41258));
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n41256), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n41256), .I0(n2316), 
            .I1(VCC_net), .CO(n41257));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n41255), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n41255), .I0(n2317), 
            .I1(VCC_net), .CO(n41256));
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n41684), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n41254), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n41684), .I0(n3212), 
            .I1(VCC_net), .CO(n41685));
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n41254), .I0(n2318), 
            .I1(VCC_net), .CO(n41255));
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5297), .I3(n40710), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n41683), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n41253), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n41253), .I0(n2319), 
            .I1(VCC_net), .CO(n41254));
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n41252), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n41252), .I0(n2320), 
            .I1(VCC_net), .CO(n41253));
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30737_3_lut (.I0(n6_adj_5358), .I1(n7611), .I2(n46297), .I3(GND_net), 
            .O(n46300));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30737_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n41683), .I0(n3213), 
            .I1(VCC_net), .CO(n41684));
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n41251), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30738_3_lut (.I0(encoder0_position[27]), .I1(n46300), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i30738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n41682), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n41682), .I0(n3214), 
            .I1(VCC_net), .CO(n41683));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n41681), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n2222), .I1(n48911), .I2(n2223), .I3(n2227), 
            .O(n48915));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n41681), .I0(n3215), 
            .I1(VCC_net), .CO(n41682));
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n41680), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n41251), .I0(n2321), 
            .I1(VCC_net), .CO(n41252));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n41250), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n40710), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5297), .CO(n40711));
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n41250), .I0(n2322), 
            .I1(VCC_net), .CO(n41251));
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n41680), .I0(n3216), 
            .I1(VCC_net), .CO(n41681));
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n41679), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n41679), .I0(n3217), 
            .I1(VCC_net), .CO(n41680));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n41249), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n41249), .I0(n2323), 
            .I1(VCC_net), .CO(n41250));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n41248), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n41248), .I0(n2324), 
            .I1(VCC_net), .CO(n41249));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n41247), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n41678), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n41247), .I0(n2325), 
            .I1(VCC_net), .CO(n41248));
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n41246), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n41246), .I0(n2326), 
            .I1(VCC_net), .CO(n41247));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n41245), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n41245), .I0(n2327), 
            .I1(VCC_net), .CO(n41246));
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n1029), .I1(n36650), .I2(n1030), .I3(n1031), 
            .O(n46564));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n41244), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n41244), .I0(n2328), 
            .I1(VCC_net), .CO(n41245));
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n41678), .I0(n3218), 
            .I1(VCC_net), .CO(n41679));
    SB_LUT4 add_145_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n40388), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n41243), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n41243), .I0(n2329), 
            .I1(GND_net), .CO(n41244));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n41242), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n41242), .I0(n2330), 
            .I1(GND_net), .CO(n41243));
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n41677), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n41677), .I0(n3219), 
            .I1(VCC_net), .CO(n41678));
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n41676), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n41676), .I0(n3220), 
            .I1(VCC_net), .CO(n41677));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n41675), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n41241), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n41241), .I0(n2331), 
            .I1(VCC_net), .CO(n41242));
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n41240), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n41675), .I0(n3221), 
            .I1(VCC_net), .CO(n41676));
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n41240), .I0(n2332), 
            .I1(GND_net), .CO(n41241));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n41674), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n41239), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n41239), .I0(n2333), 
            .I1(VCC_net), .CO(n41240));
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n30200));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF read_189 (.Q(read), .C(CLK_c), .D(n48385));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2187__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36996_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52631));
    defparam i36996_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n3022), .I1(n3027), .I2(n3021), .I3(n3023), 
            .O(n49071));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1734 (.I0(n3020), .I1(n3019), .I2(n3024), .I3(GND_net), 
            .O(n49069));
    defparam i1_3_lut_adj_1734.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n3016), .I1(n3017), .I2(n3018), .I3(n3026), 
            .O(n49093));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 i23016_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n36700));
    defparam i23016_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n49069), .I1(n49071), .I2(n3025), .I3(n3028), 
            .O(n49075));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n3029), .I1(n36700), .I2(n3030), .I3(n3031), 
            .O(n46707));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n3013), .I1(n3015), .I2(n46707), .I3(n49075), 
            .O(n49081));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097_adj_5370), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n3008), .I1(n3010), .I2(n3014), .I3(n49093), 
            .O(n49099));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n3009), .I1(n3011), .I2(n3012), .I3(n49081), 
            .O(n49087));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36999_4_lut (.I0(n3006), .I1(n49087), .I2(n49099), .I3(n3007), 
            .O(n3039));
    defparam i36999_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36930_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52565));
    defparam i36930_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n2229), .I1(n36740), .I2(n2230), .I3(n2231), 
            .O(n46649));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'ha080;
    SB_LUT4 i36505_4_lut (.I0(n1026), .I1(n46564), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i36505_4_lut.LUT_INIT = 16'h0001;
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n7066), 
            .D(n1092), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23099_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n36786));
    defparam i23099_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1742 (.I0(n50109), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n48615));
    defparam i1_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1743 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n48779));
    defparam i1_2_lut_adj_1743.LUT_INIT = 16'h8888;
    SB_LUT4 i36519_4_lut (.I0(n48779), .I1(n1125), .I2(n48615), .I3(n36786), 
            .O(n1158));
    defparam i36519_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096_adj_5369), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22903_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n36584));
    defparam i22903_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1744 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n48793));
    defparam i1_3_lut_adj_1744.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n1229), .I1(n36584), .I2(n1230), .I3(n1231), 
            .O(n46559));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n41239));
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n41674), .I0(n3222), 
            .I1(VCC_net), .CO(n41675));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n41673), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n41673), .I0(n3223), 
            .I1(VCC_net), .CO(n41674));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n41672), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n41672), .I0(n3224), 
            .I1(VCC_net), .CO(n41673));
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n41671), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n41671), .I0(n3225), 
            .I1(VCC_net), .CO(n41672));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n41670), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5296), .I3(n40709), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n41670), .I0(n3226), 
            .I1(VCC_net), .CO(n41671));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n41669), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n40709), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5296), .CO(n40710));
    SB_CARRY add_145_30 (.CI(n40409), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n40410));
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n41669), .I0(n3227), 
            .I1(VCC_net), .CO(n41670));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n41668), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36896_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52531));
    defparam i36896_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n41668), .I0(n3228), 
            .I1(VCC_net), .CO(n41669));
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n52391), .I1(n2214), 
            .I2(VCC_net), .I3(n41228), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n41227), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5295), .I3(n40708), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n41227), .I0(n2215), 
            .I1(VCC_net), .CO(n41228));
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n41226), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n41226), .I0(n2216), 
            .I1(VCC_net), .CO(n41227));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n40708), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5295), .CO(n40709));
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n41225), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_9 (.CI(n40388), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n40389));
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n41225), .I0(n2217), 
            .I1(VCC_net), .CO(n41226));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n41224), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n41224), .I0(n2218), 
            .I1(VCC_net), .CO(n41225));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_3 (.CI(n40382), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n40383));
    SB_LUT4 unary_minus_10_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n41223), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n41223), .I0(n2219), 
            .I1(VCC_net), .CO(n41224));
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n41667), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n41222), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n41222), .I0(n2220), 
            .I1(VCC_net), .CO(n41223));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n41221), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n41667), .I0(n3229), 
            .I1(GND_net), .CO(n41668));
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n41221), .I0(n2221), 
            .I1(VCC_net), .CO(n41222));
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n41666), .O(n51068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n41666), .I0(n3230), 
            .I1(GND_net), .CO(n41667));
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n41220), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n41220), .I0(n2222), 
            .I1(VCC_net), .CO(n41221));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5294), .I3(n40707), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n40707), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5294), .CO(n40708));
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n41219), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n41219), .I0(n2223), 
            .I1(VCC_net), .CO(n41220));
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n41665), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n41218), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n41218), .I0(n2224), 
            .I1(VCC_net), .CO(n41219));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n41217), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n41665), .I0(n3231), 
            .I1(VCC_net), .CO(n41666));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n41664), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n41664), .I0(n3232), 
            .I1(GND_net), .CO(n41665));
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n41217), .I0(n2225), 
            .I1(VCC_net), .CO(n41218));
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n41663), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n41216), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n41216), .I0(n2226), 
            .I1(VCC_net), .CO(n41217));
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n41215), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n41663), .I0(n3233), 
            .I1(VCC_net), .CO(n41664));
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n41215), .I0(n2227), 
            .I1(VCC_net), .CO(n41216));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n41214), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n41214), .I0(n2228), 
            .I1(VCC_net), .CO(n41215));
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n41213), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n40408), .O(n1081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n41213), .I0(n2229), 
            .I1(GND_net), .CO(n41214));
    SB_CARRY add_145_29 (.CI(n40408), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n40409));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n41212), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n41212), .I0(n2230), 
            .I1(GND_net), .CO(n41213));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n41211), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n41662), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n41211), .I0(n2231), 
            .I1(VCC_net), .CO(n41212));
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n41210), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n41210), .I0(n2232), 
            .I1(GND_net), .CO(n41211));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n41209), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n41209), .I0(n2233), 
            .I1(VCC_net), .CO(n41210));
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n41209));
    SB_LUT4 add_145_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n40387), .O(n1102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n52366), .I1(n2115), 
            .I2(VCC_net), .I3(n41208), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n41207), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n41207), .I0(n2116), 
            .I1(VCC_net), .CO(n41208));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n41206), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n40407), .O(n1082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5293), .I3(n40706), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_28 (.CI(n40407), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n40408));
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n41206), .I0(n2117), 
            .I1(VCC_net), .CO(n41207));
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n41205), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n41662), .I0(n957), 
            .I1(GND_net), .CO(n41663));
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n41205), .I0(n2118), 
            .I1(VCC_net), .CO(n41206));
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n41204), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n41204), .I0(n2119), 
            .I1(VCC_net), .CO(n41205));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n41203), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n41203), .I0(n2120), 
            .I1(VCC_net), .CO(n41204));
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n41202), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n41202), .I0(n2121), 
            .I1(VCC_net), .CO(n41203));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n41201), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n41201), .I0(n2122), 
            .I1(VCC_net), .CO(n41202));
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n2220), .I1(n46649), .I2(n2221), .I3(n48915), 
            .O(n48921));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n41200), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n41662));
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n41200), .I0(n2123), 
            .I1(VCC_net), .CO(n41201));
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n48921), 
            .O(n48927));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i36760_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n48927), 
            .O(n2247));
    defparam i36760_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n41199), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n41199), .I0(n2124), 
            .I1(VCC_net), .CO(n41200));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n41198), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n41198), .I0(n2125), 
            .I1(VCC_net), .CO(n41199));
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n41197), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n41197), .I0(n2126), 
            .I1(VCC_net), .CO(n41198));
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n2326), .I1(n2324), .I2(n2327), .I3(n2325), 
            .O(n48517));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n41196), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n41196), .I0(n2127), 
            .I1(VCC_net), .CO(n41197));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n41195), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1749 (.I0(n2322), .I1(n2328), .I2(n2323), .I3(GND_net), 
            .O(n48519));
    defparam i1_3_lut_adj_1749.LUT_INIT = 16'hfefe;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n7066), 
            .D(n1093), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n41195), .I0(n2128), 
            .I1(VCC_net), .CO(n41196));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n41194), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n41194), .I0(n2129), 
            .I1(GND_net), .CO(n41195));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n41193), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n41193), .I0(n2130), 
            .I1(GND_net), .CO(n41194));
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n41192), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n41192), .I0(n2131), 
            .I1(VCC_net), .CO(n41193));
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n41191), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n41191), .I0(n2132), 
            .I1(GND_net), .CO(n41192));
    SB_LUT4 add_145_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n40406), .O(n1083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n41190), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n41190), .I0(n2133), 
            .I1(VCC_net), .CO(n41191));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n41190));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n52665), .I1(n3105), 
            .I2(VCC_net), .I3(n41661), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_145_27 (.CI(n40406), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n40407));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n52342), .I1(n2016), 
            .I2(VCC_net), .I3(n41189), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n41188), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16569_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30258));   // verilog/coms.v(127[12] 300[6])
    defparam i16569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_8 (.CI(n40387), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n40388));
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n41188), .I0(n2017), 
            .I1(VCC_net), .CO(n41189));
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n41187), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n41187), .I0(n2018), 
            .I1(VCC_net), .CO(n41188));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n41186), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n41186), .I0(n2019), 
            .I1(VCC_net), .CO(n41187));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n41185), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n41185), .I0(n2020), 
            .I1(VCC_net), .CO(n41186));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n41184), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n41184), .I0(n2021), 
            .I1(VCC_net), .CO(n41185));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n41183), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n41183), .I0(n2022), 
            .I1(VCC_net), .CO(n41184));
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n41182), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n40405), .O(n1084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n41182), .I0(n2023), 
            .I1(VCC_net), .CO(n41183));
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n41181), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16570_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30259));   // verilog/coms.v(127[12] 300[6])
    defparam i16570_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_26 (.CI(n40405), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n40406));
    SB_LUT4 add_145_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n40404), .O(n1085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n41181), .I0(n2024), 
            .I1(VCC_net), .CO(n41182));
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n41660), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16571_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n29618), .I3(GND_net), .O(n30260));   // verilog/coms.v(127[12] 300[6])
    defparam i16571_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n41660), .I0(n3106), 
            .I1(VCC_net), .CO(n41661));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n41659), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025_adj_5377), 
            .I2(VCC_net), .I3(n41180), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n41180), .I0(n2025_adj_5377), 
            .I1(VCC_net), .CO(n41181));
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n41179), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n40706), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5293), .CO(n40707));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5291), .I3(n40705), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n41659), .I0(n3107), 
            .I1(VCC_net), .CO(n41660));
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n41179), .I0(n2026), 
            .I1(VCC_net), .CO(n41180));
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n41178), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n40705), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5291), .CO(n40706));
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n41178), .I0(n2027), 
            .I1(VCC_net), .CO(n41179));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5290), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_10 (.CI(n40420), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n40421));
    SB_CARRY add_145_25 (.CI(n40404), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n40405));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19), .I2(encoder0_position[31]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n41177), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n41177), .I0(n2028), 
            .I1(VCC_net), .CO(n41178));
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23145_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n36832));
    defparam i23145_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n41176), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n41658), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n41176), .I0(n2029), 
            .I1(GND_net), .CO(n41177));
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n41175), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n41175), .I0(n2030), 
            .I1(GND_net), .CO(n41176));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n41174), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n41658), .I0(n3108), 
            .I1(VCC_net), .CO(n41659));
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n41174), .I0(n2031), 
            .I1(VCC_net), .CO(n41175));
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n41173), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n41173), .I0(n2032), 
            .I1(GND_net), .CO(n41174));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n41172), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n41657), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n41172), .I0(n2033), 
            .I1(VCC_net), .CO(n41173));
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5290), .CO(n40705));
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n41172));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n52319), .I1(n1917), 
            .I2(VCC_net), .I3(n41171), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n41170), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n41170), .I0(n1918), 
            .I1(VCC_net), .CO(n41171));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n41169), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n41169), .I0(n1919), 
            .I1(VCC_net), .CO(n41170));
    SB_LUT4 encoder0_position_31__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36534_4_lut (.I0(n1225), .I1(n1224), .I2(n46559), .I3(n48793), 
            .O(n1257));
    defparam i36534_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_5319), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n941));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n41168), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n40403), .O(n1086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n41168), .I0(n1920), 
            .I1(VCC_net), .CO(n41169));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n41167), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n41167), .I0(n1921), 
            .I1(VCC_net), .CO(n41168));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n41166), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n2320), .I1(n2321), .I2(n48519), .I3(n48517), 
            .O(n48525));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n41166), .I0(n1922), 
            .I1(VCC_net), .CO(n41167));
    SB_LUT4 i1_2_lut_adj_1751 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n48903));
    defparam i1_2_lut_adj_1751.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n41165), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n41165), .I0(n1923), 
            .I1(VCC_net), .CO(n41166));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n41164), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n41164), .I0(n1924), 
            .I1(VCC_net), .CO(n41165));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n41163), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n41163), .I0(n1925), 
            .I1(VCC_net), .CO(n41164));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n41162), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n41162), .I0(n1926), 
            .I1(VCC_net), .CO(n41163));
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n48903), .I1(n2319), .I2(n48525), .I3(n36832), 
            .O(n48529));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'hfefc;
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n41161), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n41161), .I0(n1927), 
            .I1(VCC_net), .CO(n41162));
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n41160), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n41160), .I0(n1928), 
            .I1(VCC_net), .CO(n41161));
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n41159), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n41159), .I0(n1929), 
            .I1(GND_net), .CO(n41160));
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n41158), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n41158), .I0(n1930), 
            .I1(GND_net), .CO(n41159));
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n41157), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n41157), .I0(n1931), 
            .I1(VCC_net), .CO(n41158));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n41156), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n41156), .I0(n1932), 
            .I1(GND_net), .CO(n41157));
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n41657), .I0(n3109), 
            .I1(VCC_net), .CO(n41658));
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n41155), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n41155), .I0(n1933), 
            .I1(VCC_net), .CO(n41156));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n41155));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n52297), .I1(n1818), 
            .I2(VCC_net), .I3(n41154), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n41153), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n41656), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n41153), .I0(n1819), 
            .I1(VCC_net), .CO(n41154));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n41152), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n41152), .I0(n1820), 
            .I1(VCC_net), .CO(n41153));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n41151), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n41151), .I0(n1821), 
            .I1(VCC_net), .CO(n41152));
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195_adj_5375), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n41150), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n41150), .I0(n1822), 
            .I1(VCC_net), .CO(n41151));
    SB_CARRY add_145_24 (.CI(n40403), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n40404));
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n41149), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n41149), .I0(n1823), 
            .I1(VCC_net), .CO(n41150));
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n41656), .I0(n3110), 
            .I1(VCC_net), .CO(n41657));
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n41148), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLA_181 (.Q(INLA_c_0), .C(CLK_c), .E(n29588), .D(GLA_N_384), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n41148), .I0(n1824), 
            .I1(VCC_net), .CO(n41149));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n41147), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n41147), .I0(n1825), 
            .I1(VCC_net), .CO(n41148));
    SB_LUT4 encoder0_position_31__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n41146), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5320), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n41146), .I0(n1826), 
            .I1(VCC_net), .CO(n41147));
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n41145), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n40402), .O(n1087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n41145), .I0(n1827), 
            .I1(VCC_net), .CO(n41146));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n41144), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n41144), .I0(n1828), 
            .I1(VCC_net), .CO(n41145));
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n41143), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n41143), .I0(n1829), 
            .I1(GND_net), .CO(n41144));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n41142), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n41142), .I0(n1830), 
            .I1(GND_net), .CO(n41143));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n41655), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n41141), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n41141), .I0(n1831), 
            .I1(VCC_net), .CO(n41142));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n41140), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n41140), .I0(n1832), 
            .I1(GND_net), .CO(n41141));
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n41139), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n41139), .I0(n1833), 
            .I1(VCC_net), .CO(n41140));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n41139));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n52276), .I1(n1719), 
            .I2(VCC_net), .I3(n41138), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n41137), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n41655), .I0(n3111), 
            .I1(VCC_net), .CO(n41656));
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n41137), .I0(n1720), 
            .I1(VCC_net), .CO(n41138));
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n41136), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n41136), .I0(n1721), 
            .I1(VCC_net), .CO(n41137));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n41135), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n41135), .I0(n1722), 
            .I1(VCC_net), .CO(n41136));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n41134), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n41654), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n41134), .I0(n1723), 
            .I1(VCC_net), .CO(n41135));
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n41133), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n40386), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n41133), .I0(n1724), 
            .I1(VCC_net), .CO(n41134));
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n41132), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16572_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n29618), .I3(GND_net), .O(n30261));   // verilog/coms.v(127[12] 300[6])
    defparam i16572_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n41132), .I0(n1725), 
            .I1(VCC_net), .CO(n41133));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n41131), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n41131), .I0(n1726), 
            .I1(VCC_net), .CO(n41132));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n41130), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_23 (.CI(n40402), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n40403));
    SB_LUT4 i4472_4_lut (.I0(n28290), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5378));
    defparam i4472_4_lut.LUT_INIT = 16'hc8c0;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n41130), .I0(n1727), 
            .I1(VCC_net), .CO(n41131));
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n41129), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n41129), .I0(n1728), 
            .I1(VCC_net), .CO(n41130));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n41128), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1753 (.I0(n24_adj_5378), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n47285));
    defparam i2_4_lut_adj_1753.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1754 (.I0(n47285), .I1(delay_counter[18]), .I2(n28292), 
            .I3(GND_net), .O(n47822));
    defparam i2_3_lut_adj_1754.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n41654), .I0(n3112), 
            .I1(VCC_net), .CO(n41655));
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n41128), .I0(n1729), 
            .I1(GND_net), .CO(n41129));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n41653), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n41653), .I0(n3113), 
            .I1(VCC_net), .CO(n41654));
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n41652), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n41652), .I0(n3114), 
            .I1(VCC_net), .CO(n41653));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n41127), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n41127), .I0(n1730), 
            .I1(GND_net), .CO(n41128));
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n41126), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16448_4_lut (.I0(state_7__N_4103[3]), .I1(data[5]), .I2(n4_adj_5272), 
            .I3(n28416), .O(n30137));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16448_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n41126), .I0(n1731), 
            .I1(VCC_net), .CO(n41127));
    SB_LUT4 i2_4_lut_adj_1755 (.I0(delay_counter[23]), .I1(n47822), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5314));
    defparam i2_4_lut_adj_1755.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1756 (.I0(n7_adj_5314), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n28287), .O(n62));
    defparam i4_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n41125), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1757 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n28292));
    defparam i2_3_lut_adj_1757.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5420));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_5420), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n28287));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1758 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_5285));
    defparam i5_3_lut_adj_1758.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n41125), .I0(n1732), 
            .I1(GND_net), .CO(n41126));
    SB_LUT4 i16449_4_lut (.I0(state_7__N_4103[3]), .I1(data[4]), .I2(n4_adj_5272), 
            .I3(n28421), .O(n30138));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16449_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6_4_lut_adj_1759 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5284));
    defparam i6_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n41124), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n41124), .I0(n1733), 
            .I1(VCC_net), .CO(n41125));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n41124));
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n52241), .I1(n1620), 
            .I2(VCC_net), .I3(n41123), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n41651), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16450_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[5]), .I2(n6_adj_5317), 
            .I3(n28437), .O(n30139));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16450_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5284), .I1(delay_counter[2]), .I2(n14_adj_5285), 
            .I3(delay_counter[6]), .O(n28290));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n41122), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n41122), .I0(n1621), 
            .I1(VCC_net), .CO(n41123));
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n41651), .I0(n3115), 
            .I1(VCC_net), .CO(n41652));
    SB_LUT4 i8374_3_lut (.I0(n62), .I1(\ID_READOUT_FSM.state [0]), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n21929));
    defparam i8374_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 add_2591_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n40555), 
            .O(n7607)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1760 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5286));
    defparam i1_2_lut_adj_1760.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n41650), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1761 (.I0(delay_counter[9]), .I1(n4_adj_5286), 
            .I2(delay_counter[10]), .I3(n28290), .O(n47398));
    defparam i2_4_lut_adj_1761.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1762 (.I0(n47398), .I1(n28292), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n47283));
    defparam i2_4_lut_adj_1762.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5432));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n41650), .I0(n3116), 
            .I1(VCC_net), .CO(n41651));
    SB_LUT4 i2_4_lut_adj_1763 (.I0(delay_counter[22]), .I1(n47283), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5433));
    defparam i2_4_lut_adj_1763.LUT_INIT = 16'ha8a0;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n41649), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n41121), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n41121), .I0(n1622), 
            .I1(VCC_net), .CO(n41122));
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n41649), .I0(n3117), 
            .I1(VCC_net), .CO(n41650));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n41648), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n41120), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22230_4_lut (.I0(n7_adj_5433), .I1(delay_counter[31]), .I2(n28287), 
            .I3(n8_adj_5432), .O(n1195));   // verilog/TinyFPGA_B.v(378[14:38])
    defparam i22230_4_lut.LUT_INIT = 16'h3230;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n41120), .I0(n1623), 
            .I1(VCC_net), .CO(n41121));
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n41119), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n41119), .I0(n1624), 
            .I1(VCC_net), .CO(n41120));
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n41118), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n41648), .I0(n3118), 
            .I1(VCC_net), .CO(n41649));
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5386));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_145_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n41118), .I0(n1625), 
            .I1(VCC_net), .CO(n41119));
    SB_LUT4 i22899_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n36580));
    defparam i22899_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n50107), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n48675));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1765 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5385));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i6_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n1329), .I1(n36580), .I2(n1330), .I3(n1331), 
            .O(n46556));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'ha080;
    SB_LUT4 i36554_4_lut (.I0(n46556), .I1(n1323), .I2(n1324), .I3(n48675), 
            .O(n1356));
    defparam i36554_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22897_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n36578));
    defparam i22897_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1767 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n48815));
    defparam i1_2_lut_adj_1767.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n1429), .I1(n36578), .I2(n1430), .I3(n1431), 
            .O(n46575));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n41117), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n41117), .I0(n1626), 
            .I1(VCC_net), .CO(n41118));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n41116), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_5385), .I2(n10_adj_5386), 
            .I3(ID[6]), .O(n28264));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2591_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n40554), 
            .O(n7608)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n41116), .I0(n1627), 
            .I1(VCC_net), .CO(n41117));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n41115), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n41115), .I0(n1628), 
            .I1(VCC_net), .CO(n41116));
    SB_CARRY add_2591_6 (.CI(n40554), .I0(n622), .I1(GND_net), .CO(n40555));
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n41114), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n41114), .I0(n1629), 
            .I1(GND_net), .CO(n41115));
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n41113), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n41113), .I0(n1630), 
            .I1(GND_net), .CO(n41114));
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n41112), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n41112), .I0(n1631), 
            .I1(VCC_net), .CO(n41113));
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632_adj_5376), 
            .I2(GND_net), .I3(n41111), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n41111), .I0(n1632_adj_5376), 
            .I1(GND_net), .CO(n41112));
    SB_LUT4 add_2591_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n40553), 
            .O(n7609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16276_4_lut (.I0(n7066), .I1(n1195), .I2(n21929), .I3(n28265), 
            .O(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16276_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n41110), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n41110), .I0(n1633), 
            .I1(VCC_net), .CO(n41111));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n41110));
    SB_CARRY add_2591_5 (.CI(n40553), .I0(n623), .I1(VCC_net), .CO(n40554));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n52222), .I1(n1521), 
            .I2(VCC_net), .I3(n41109), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n41108), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2591_4_lut (.I0(GND_net), .I1(n405), .I2(GND_net), .I3(n40552), 
            .O(n7610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n41108), .I0(n1522), 
            .I1(VCC_net), .CO(n41109));
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n41107), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n41107), .I0(n1523), 
            .I1(VCC_net), .CO(n41108));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n50105), 
            .I2(VCC_net), .I3(n41106), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n41106), .I0(n50105), 
            .I1(VCC_net), .CO(n41107));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n41105), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n41105), .I0(n1525), 
            .I1(VCC_net), .CO(n41106));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n41104), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n41104), .I0(n1526), 
            .I1(VCC_net), .CO(n41105));
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n41647), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16515_3_lut (.I0(current[9]), .I1(data_adj_5497[9]), .I2(n47264), 
            .I3(GND_net), .O(n30204));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n41103), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n41103), .I0(n1527), 
            .I1(VCC_net), .CO(n41104));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n41102), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n41102), .I0(n1528), 
            .I1(VCC_net), .CO(n41103));
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n41647), .I0(n3119), 
            .I1(VCC_net), .CO(n41648));
    SB_CARRY add_145_7 (.CI(n40386), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n40387));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n41101), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n41101), .I0(n1529), 
            .I1(GND_net), .CO(n41102));
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n41100), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n41100), .I0(n1530), 
            .I1(GND_net), .CO(n41101));
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n41099), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n41646), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n48815), 
            .O(n48821));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n41099), .I0(n1531), 
            .I1(VCC_net), .CO(n41100));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n41098), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n41098), .I0(n1532), 
            .I1(GND_net), .CO(n41099));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n41097), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n41097), .I0(n1533), 
            .I1(VCC_net), .CO(n41098));
    SB_CARRY add_2591_4 (.CI(n40552), .I0(n405), .I1(GND_net), .CO(n40553));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n41646), .I0(n3120), 
            .I1(VCC_net), .CO(n41647));
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n41097));
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n52200), .I1(n1422), 
            .I2(VCC_net), .I3(n41096), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n41095), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16516_3_lut (.I0(current[8]), .I1(data_adj_5497[8]), .I2(n47264), 
            .I3(GND_net), .O(n30205));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2591_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n40551), 
            .O(n7611)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2591_3 (.CI(n40551), .I0(n625), .I1(VCC_net), .CO(n40552));
    SB_LUT4 add_2591_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7612)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2591_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2591_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n40551));
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n41095), .I0(n1423), 
            .I1(VCC_net), .CO(n41096));
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n48529), 
            .O(n48535));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 add_145_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n40401), .O(n1088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n41094), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n41094), .I0(n1424), 
            .I1(VCC_net), .CO(n41095));
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n41093), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36571_4_lut (.I0(n1423), .I1(n1422), .I2(n48821), .I3(n46575), 
            .O(n1455));
    defparam i36571_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n41093), .I0(n1425), 
            .I1(VCC_net), .CO(n41094));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n41092), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n41092), .I0(n1426), 
            .I1(VCC_net), .CO(n41093));
    SB_CARRY add_145_22 (.CI(n40401), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n40402));
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n41645), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n41091), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n41091), .I0(n1427), 
            .I1(VCC_net), .CO(n41092));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n41090), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n41645), .I0(n3121), 
            .I1(VCC_net), .CO(n41646));
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n41090), .I0(n1428), 
            .I1(VCC_net), .CO(n41091));
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n41089), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n41089), .I0(n1429), 
            .I1(GND_net), .CO(n41090));
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n41088), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n41088), .I0(n1430), 
            .I1(GND_net), .CO(n41089));
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n41087), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n41644), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n41087), .I0(n1431), 
            .I1(VCC_net), .CO(n41088));
    SB_LUT4 i6909_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_403));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i6909_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n41086), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n41086), .I0(n1432), 
            .I1(GND_net), .CO(n41087));
    SB_LUT4 i6911_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_412));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i6911_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n41085), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n41644), .I0(n3122), 
            .I1(VCC_net), .CO(n41645));
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n41085), .I0(n1433), 
            .I1(VCC_net), .CO(n41086));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n41085));
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n41643), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n41643), .I0(n3123), 
            .I1(VCC_net), .CO(n41644));
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1771 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n48619));
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'heeee;
    SB_LUT4 i23084_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n36770));
    defparam i23084_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n50105), .I1(n1525), .I2(n1526), .I3(n48619), 
            .O(n48625));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n1529), .I1(n48625), .I2(n36770), .I3(n1530), 
            .O(n48627));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n41642), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n40775), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n41642), .I0(n3124), 
            .I1(VCC_net), .CO(n41643));
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n40774), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n40774), .I0(n829), 
            .I1(GND_net), .CO(n40775));
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n41641), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n41641), .I0(n3125), 
            .I1(VCC_net), .CO(n41642));
    SB_LUT4 add_145_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n40400), .O(n1089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n41640), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n40773), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n40773), .I0(n830), 
            .I1(GND_net), .CO(n40774));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n40772), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n40772), .I0(n831), 
            .I1(VCC_net), .CO(n40773));
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n52184), .I1(n1323), 
            .I2(VCC_net), .I3(n41074), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n40771), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n40771), .I0(n832), 
            .I1(GND_net), .CO(n40772));
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n41073), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n41073), .I0(n1324), 
            .I1(VCC_net), .CO(n41074));
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n50107), 
            .I2(VCC_net), .I3(n41072), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n41072), .I0(n50107), 
            .I1(VCC_net), .CO(n41073));
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n41640), .I0(n3126), 
            .I1(VCC_net), .CO(n41641));
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n41071), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n41639), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n41071), .I0(n1326), 
            .I1(VCC_net), .CO(n41072));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n40770), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n40770), .I0(n833), 
            .I1(VCC_net), .CO(n40771));
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n41070), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n41639), .I0(n3127), 
            .I1(VCC_net), .CO(n41640));
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n41070), .I0(n1327), 
            .I1(VCC_net), .CO(n41071));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n41069), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_21 (.CI(n40400), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n40401));
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n41069), .I0(n1328), 
            .I1(VCC_net), .CO(n41070));
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n41068), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n41068), .I0(n1329), 
            .I1(GND_net), .CO(n41069));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n41067), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n41067), .I0(n1330), 
            .I1(GND_net), .CO(n41068));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n41066), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n41066), .I0(n1331), 
            .I1(VCC_net), .CO(n41067));
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n41065), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n41065), .I0(n1332), 
            .I1(GND_net), .CO(n41066));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n41064), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n40770));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n41638), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n41064), .I0(n1333), 
            .I1(VCC_net), .CO(n41065));
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n41064));
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n41638), .I0(n3128), 
            .I1(VCC_net), .CO(n41639));
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n52165), .I1(n1224), 
            .I2(VCC_net), .I3(n41063), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n41062), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n41062), .I0(n1225), 
            .I1(VCC_net), .CO(n41063));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n41061), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n41061), .I0(n1226), 
            .I1(VCC_net), .CO(n41062));
    SB_LUT4 i16573_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n29618), .I3(GND_net), .O(n30262));   // verilog/coms.v(127[12] 300[6])
    defparam i16573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n41060), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n7066), 
            .D(n1094), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n7066), 
            .D(n1095), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16574_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n29618), .I3(GND_net), .O(n30263));   // verilog/coms.v(127[12] 300[6])
    defparam i16574_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n41060), .I0(n1227), 
            .I1(VCC_net), .CO(n41061));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n41059), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n41059), .I0(n1228), 
            .I1(VCC_net), .CO(n41060));
    SB_LUT4 add_145_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n40385), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n41058), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n41058), .I0(n1229), 
            .I1(GND_net), .CO(n41059));
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n41057), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n41057), .I0(n1230), 
            .I1(GND_net), .CO(n41058));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n41637), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n41056), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n41056), .I0(n1231), 
            .I1(VCC_net), .CO(n41057));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n41055), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n41055), .I0(n1232), 
            .I1(GND_net), .CO(n41056));
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n41637), .I0(n3129), 
            .I1(GND_net), .CO(n41638));
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n41054), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n41054), .I0(n1233), 
            .I1(VCC_net), .CO(n41055));
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n41054));
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n52150), .I1(n1125), 
            .I2(VCC_net), .I3(n41053), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n41636), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n41636), .I0(n3130), 
            .I1(GND_net), .CO(n41637));
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n50109), 
            .I2(VCC_net), .I3(n41052), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n41052), .I0(n50109), 
            .I1(VCC_net), .CO(n41053));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n41051), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n41051), .I0(n1127), 
            .I1(VCC_net), .CO(n41052));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n41050), .O(n1195_adj_5375)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n41050), .I0(n1128), 
            .I1(VCC_net), .CO(n41051));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5298));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n41049), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n41049), .I0(n1129), 
            .I1(GND_net), .CO(n41050));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n41048), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n41048), .I0(n1130), 
            .I1(GND_net), .CO(n41049));
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n7066), 
            .D(n1096), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n41047), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n41047), .I0(n1131), 
            .I1(VCC_net), .CO(n41048));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n41046), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n41046), .I0(n1132), 
            .I1(GND_net), .CO(n41047));
    SB_LUT4 i35617_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n51093));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35617_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35692_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n51107));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35692_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35623_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n51108));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35623_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35622_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n51109));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35622_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n41045), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n41045), .I0(n1133), 
            .I1(VCC_net), .CO(n41046));
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n41045));
    SB_LUT4 i35621_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n51110));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35621_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35620_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n51111));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35620_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35619_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n51112));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35619_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i35618_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n51113));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i35618_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5288), 
            .I2(commutation_state_prev[0]), .I3(dti_N_416), .O(n29564));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_DFFESR GLB_183 (.Q(INLB_c_0), .C(CLK_c), .E(n29588), .D(GLB_N_398), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFFESR GLC_185 (.Q(INLC_c_0), .C(CLK_c), .E(n29588), .D(GLC_N_412), 
            .R(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i22087_1_lut_2_lut (.I0(n25788), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n1958));
    defparam i22087_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n41635), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n45412));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n44714));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n30753));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n30752));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n30751));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n30750));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n30749));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n30748));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n30747));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1774 (.I0(n3807), .I1(tx_transmit_N_3513), 
            .I2(n2025), .I3(n28383), .O(n45649));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1774.LUT_INIT = 16'haafe;
    SB_LUT4 i36786_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n48535), 
            .O(n2346));
    defparam i36786_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30771_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n46335));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i30771_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16575_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n29618), .I3(GND_net), .O(n30264));   // verilog/coms.v(127[12] 300[6])
    defparam i16575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6901_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_367));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6901_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i6903_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_384));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6903_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i6905_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_389));
    defparam i6905_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n41011), .O(n1093_adj_5366)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16576_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n29618), .I3(GND_net), .O(n30265));   // verilog/coms.v(127[12] 300[6])
    defparam i16576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16577_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n29618), .I3(GND_net), .O(n30266));   // verilog/coms.v(127[12] 300[6])
    defparam i16577_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n41635), .I0(n3131), 
            .I1(VCC_net), .CO(n41636));
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n41010), .O(n1094_adj_5367)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16578_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n29618), .I3(GND_net), .O(n30267));   // verilog/coms.v(127[12] 300[6])
    defparam i16578_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n41010), .I0(n1027), 
            .I1(VCC_net), .CO(n41011));
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n41009), .O(n1095_adj_5368)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n41009), .I0(n1028), 
            .I1(VCC_net), .CO(n41010));
    SB_LUT4 i6907_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_398));
    defparam i6907_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n41008), .O(n1096_adj_5369)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5288));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'h7bde;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n41008), .I0(n1029), 
            .I1(GND_net), .CO(n41009));
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n41007), .O(n1097_adj_5370)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n41007), .I0(n1030), 
            .I1(GND_net), .CO(n41008));
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n41006), .O(n1098_adj_5371)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5412));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n41006), .I0(n1031), 
            .I1(VCC_net), .CO(n41007));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n41005), .O(n1099_adj_5372)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_215), 
            .I3(n40489), .O(pwm_setpoint_23__N_191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n40399), .O(n1090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2187__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54_adj_5382));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n41005), .I0(n1032), 
            .I1(GND_net), .CO(n41006));
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n41004), .O(n1100_adj_5373)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_20 (.CI(n40399), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n40400));
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n41004), .I0(n1033), 
            .I1(VCC_net), .CO(n41005));
    SB_LUT4 unary_minus_10_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3), 
            .I3(n40488), .O(pwm_setpoint_23__N_191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101_adj_5374)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5411));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36810_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52445));
    defparam i36810_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n41634), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_adj_1776 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5365));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i2_2_lut_adj_1776.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n41004));
    SB_LUT4 i6_4_lut_adj_1777 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5363));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i6_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 add_145_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n40398), .O(n1091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n40382));
    SB_LUT4 i7_4_lut_adj_1778 (.I0(dti_counter[0]), .I1(n14_adj_5363), .I2(n10_adj_5365), 
            .I3(dti_counter[3]), .O(n25788));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i7_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_CARRY add_145_6 (.CI(n40385), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n40386));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5410));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5299));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_24 (.CI(n40488), .I0(GND_net), .I1(n3), 
            .CO(n40489));
    SB_LUT4 i36492_2_lut (.I0(n25788), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_416));
    defparam i36492_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5329), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4_adj_5273), 
            .I3(n40487), .O(pwm_setpoint_23__N_191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n41634), .I0(n3132), 
            .I1(GND_net), .CO(n41635));
    SB_CARRY add_145_19 (.CI(n40398), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n40399));
    SB_LUT4 encoder0_position_31__I_0_i845_rep_54_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i845_rep_54_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n41633), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1180_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5409));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n2423), .I1(n2427), .I2(n2422), .I3(n2425), 
            .O(n48945));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n2426), .I1(n48945), .I2(n2428), .I3(n2424), 
            .O(n48947));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i23143_4_lut (.I0(n949), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n36830));
    defparam i23143_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n2419), .I1(n2420), .I2(n48947), .I3(n2421), 
            .O(n48953));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i36592_4_lut (.I0(n1522), .I1(n1521), .I2(n48627), .I3(n1523), 
            .O(n1554));
    defparam i36592_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1782 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n49155));
    defparam i1_2_lut_adj_1782.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n2418), .I1(n49155), .I2(n48953), .I3(n36830), 
            .O(n48957));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n48957), 
            .O(n48963));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 i36813_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n48963), 
            .O(n2445));
    defparam i36813_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_rep_41_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n50105));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i972_rep_41_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n2522), .I1(n2525), .I2(n2528), .I3(n2527), 
            .O(n48753));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n2524), .I1(n2520), .I2(n2526), .I3(n2523), 
            .O(n47555));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 i23038_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n36722));
    defparam i23038_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n47555), .I1(n2519), .I2(n48753), .I3(n2521), 
            .O(n48759));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n2529), .I1(n36722), .I2(n2530), .I3(n2531), 
            .O(n46638));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n2517), .I1(n46638), .I2(n2518), .I3(n48759), 
            .O(n48765));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n48765), 
            .O(n48771));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i36841_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n48771), 
            .O(n2544));
    defparam i36841_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23028_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n36712));
    defparam i23028_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1791 (.I0(n2626), .I1(n2625), .I2(GND_net), .I3(GND_net), 
            .O(n48977));
    defparam i1_2_lut_adj_1791.LUT_INIT = 16'heeee;
    SB_LUT4 i22893_3_lut (.I0(n941), .I1(n1632_adj_5376), .I2(n1633), 
            .I3(GND_net), .O(n36574));
    defparam i22893_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n2624), .I1(n2628), .I2(n2622), .I3(n2627), 
            .O(n48981));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n2621), .I1(n48981), .I2(n48977), .I3(n2623), 
            .O(n48985));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n48831));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n2629), .I1(n36712), .I2(n2630), .I3(n2631), 
            .O(n46679));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n1629), .I1(n36574), .I2(n1630), .I3(n1631), 
            .O(n46584));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n2618), .I1(n2619), .I2(n2620), .I3(n48985), 
            .O(n48991));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n2616), .I1(n2617), .I2(n48991), .I3(n46679), 
            .O(n48997));
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n48997), 
            .O(n49003));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n46335));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5388), .I3(n41938), .O(n2_adj_5362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5389), .I3(n41937), .O(n3_adj_5361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n41937), 
            .I0(GND_net), .I1(n3_adj_5389), .CO(n41938));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5390), .I3(n41936), .O(n4_adj_5360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n41936), 
            .I0(GND_net), .I1(n4_adj_5390), .CO(n41937));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5391), .I3(n41935), .O(n5_adj_5359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n41935), 
            .I0(GND_net), .I1(n5_adj_5391), .CO(n41936));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5392), .I3(n41934), .O(n6_adj_5358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n41934), 
            .I0(GND_net), .I1(n6_adj_5392), .CO(n41935));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5393), .I3(n41933), .O(n7_adj_5357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n41933), 
            .I0(GND_net), .I1(n7_adj_5393), .CO(n41934));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5394), .I3(n41932), .O(n8_adj_5348)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n41932), 
            .I0(GND_net), .I1(n8_adj_5394), .CO(n41933));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5395), .I3(n41931), .O(n9_adj_5343)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n41931), 
            .I0(GND_net), .I1(n9_adj_5395), .CO(n41932));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5396), .I3(n41930), .O(n10_adj_5342)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n41930), 
            .I0(GND_net), .I1(n10_adj_5396), .CO(n41931));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5397), .I3(n41929), .O(n11_adj_5330)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n41929), 
            .I0(GND_net), .I1(n11_adj_5397), .CO(n41930));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5398), .I3(n41928), .O(n12_adj_5329)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n41928), 
            .I0(GND_net), .I1(n12_adj_5398), .CO(n41929));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5399), .I3(n41927), .O(n13_adj_5328)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n41927), 
            .I0(GND_net), .I1(n13_adj_5399), .CO(n41928));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5400), .I3(n41926), .O(n14_adj_5327)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n41926), 
            .I0(GND_net), .I1(n14_adj_5400), .CO(n41927));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5401), .I3(n41925), .O(n15_adj_5320)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n41925), 
            .I0(GND_net), .I1(n15_adj_5401), .CO(n41926));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5402), .I3(n41924), .O(n16_adj_5319)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n41924), 
            .I0(GND_net), .I1(n16_adj_5402), .CO(n41925));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5403), .I3(n41923), .O(n17_adj_5318)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n41923), 
            .I0(GND_net), .I1(n17_adj_5403), .CO(n41924));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5404), .I3(n41922), .O(n18_adj_5282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n41922), 
            .I0(GND_net), .I1(n18_adj_5404), .CO(n41923));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5405), .I3(n41921), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n41921), 
            .I0(GND_net), .I1(n19_adj_5405), .CO(n41922));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5406), .I3(n41920), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n41920), 
            .I0(GND_net), .I1(n20_adj_5406), .CO(n41921));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5407), .I3(n41919), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n41919), 
            .I0(GND_net), .I1(n21_adj_5407), .CO(n41920));
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5408), .I3(n41918), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n41918), 
            .I0(GND_net), .I1(n22_adj_5408), .CO(n41919));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5409), .I3(n41917), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36870_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n49003), 
            .O(n2643));
    defparam i36870_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n41917), 
            .I0(GND_net), .I1(n23_adj_5409), .CO(n41918));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5410), .I3(n41916), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n41916), 
            .I0(GND_net), .I1(n24_adj_5410), .CO(n41917));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5411), .I3(n41915), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n41915), 
            .I0(GND_net), .I1(n25_adj_5411), .CO(n41916));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5412), .I3(n41914), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5300));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n41914), 
            .I0(GND_net), .I1(n26_adj_5412), .CO(n41915));
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n7066), 
            .D(n1097), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5413), .I3(n41913), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n41913), 
            .I0(GND_net), .I1(n27_adj_5413), .CO(n41914));
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n7066), 
            .D(n1098), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5414), .I3(n41912), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5408));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n41912), 
            .I0(GND_net), .I1(n28_adj_5414), .CO(n41913));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5415), .I3(n41911), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n41911), 
            .I0(GND_net), .I1(n29_adj_5415), .CO(n41912));
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n7066), 
            .D(n1099), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5416), .I3(n41910), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n41910), 
            .I0(GND_net), .I1(n30_adj_5416), .CO(n41911));
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n7066), 
            .D(n1100), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5417), .I3(n41909), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n41909), 
            .I0(GND_net), .I1(n31_adj_5417), .CO(n41910));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5418), .I3(n41908), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n41908), 
            .I0(GND_net), .I1(n32_adj_5418), .CO(n41909));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5419), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5419), .CO(n41908));
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n7066), 
            .D(n1101), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF dti_counter_2187__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5301));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n1623), .I1(n46584), .I2(n1624), .I3(n48831), 
            .O(n48837));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 i36625_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n48837), 
            .O(n1653));
    defparam i36625_4_lut.LUT_INIT = 16'h0001;
    SB_DFF dti_counter_2187__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2187__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2187__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2187__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2187__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20), .I2(encoder0_position[31]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dir_175 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n7066), 
            .D(n1102), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n41633), .I0(n3133), 
            .I1(VCC_net), .CO(n41634));
    SB_LUT4 add_145_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n40397), .O(n1092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_23 (.CI(n40487), .I0(GND_net), .I1(n4_adj_5273), 
            .CO(n40488));
    SB_LUT4 unary_minus_10_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5), 
            .I3(n40486), .O(pwm_setpoint_23__N_191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_22 (.CI(n40486), .I0(GND_net), .I1(n5), 
            .CO(n40487));
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n41633));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5407));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6), 
            .I3(n40485), .O(pwm_setpoint_23__N_191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1858_rep_14_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1858_rep_14_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5302));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25), .I2(encoder0_position[31]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5406));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_18 (.CI(n40397), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n40398));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24), .I2(encoder0_position[31]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_21 (.CI(n40485), .I0(GND_net), .I1(n6), 
            .CO(n40486));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5303));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n40396), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5405));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7), 
            .I3(n40484), .O(pwm_setpoint_23__N_191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_17 (.CI(n40396), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n40397));
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(GND_net), .I1(n3006), 
            .I2(VCC_net), .I3(n41632), .O(n3073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n41631), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5304));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5305));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n40395), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_5318), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n942));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_16 (.CI(n40395), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n40396));
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n41631), .I0(n3007), 
            .I1(VCC_net), .CO(n41632));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n41630), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5421));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1801 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_216[0]));   // verilog/TinyFPGA_B.v(148[4] 150[7])
    defparam i1_3_lut_adj_1801.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n41630), .I0(n3008), 
            .I1(VCC_net), .CO(n41631));
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1039_rep_51_3_lut (.I0(n50105), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1039_rep_51_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1802 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5289), .I3(control_mode[2]), .O(n28252));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam i1_2_lut_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5404));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23026_3_lut (.I0(n952), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n36710));
    defparam i23026_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_5282), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n943));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n41629), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5306));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36502_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52137));
    defparam i36502_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1803 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n48691));
    defparam i1_3_lut_adj_1803.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_20 (.CI(n40484), .I0(GND_net), .I1(n7), 
            .CO(n40485));
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8), 
            .I3(n40483), .O(pwm_setpoint_23__N_191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5388));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5307));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1804 (.I0(n2725), .I1(n2720), .I2(n2727), .I3(GND_net), 
            .O(n48641));
    defparam i1_3_lut_adj_1804.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n41629), .I0(n3009), 
            .I1(VCC_net), .CO(n41630));
    SB_LUT4 add_145_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n40394), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21), .I2(encoder0_position[31]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23076_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n36762));
    defparam i23076_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n41628), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5403));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21932_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i21932_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n1723), .I1(n1724), .I2(n48691), .I3(n1725), 
            .O(n48697));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n2723), .I1(n2721), .I2(n2726), .I3(n2728), 
            .O(n48643));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i21931_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i21931_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_10_add_3_19 (.CI(n40483), .I0(GND_net), .I1(n8), 
            .CO(n40484));
    SB_LUT4 i22319_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i22319_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5308));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16517_3_lut (.I0(current[7]), .I1(data_adj_5497[7]), .I2(n47264), 
            .I3(GND_net), .O(n30206));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n40482), .O(pwm_setpoint_23__N_191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5309));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n41628), .I0(n3010), 
            .I1(VCC_net), .CO(n41629));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5402));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n41627), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_18 (.CI(n40482), .I0(GND_net), .I1(n9), 
            .CO(n40483));
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1807 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n48865));
    defparam i1_2_lut_adj_1807.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5310));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n48643), .I1(n48641), .I2(n2722), .I3(n2724), 
            .O(n48647));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5311));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_5328), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5401));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i913_rep_42_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i913_rep_42_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n41627), .I0(n3011), 
            .I1(VCC_net), .CO(n41628));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n41626), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n2729), .I1(n36710), .I2(n2730), .I3(n2731), 
            .O(n46644));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'ha080;
    SB_CARRY add_145_15 (.CI(n40394), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n40395));
    motorControl control (.GND_net(GND_net), .\Ki[2] (Ki[2]), .\Ki[0] (Ki[0]), 
            .\Ki[1] (Ki[1]), .\Ki[3] (Ki[3]), .PWMLimit({PWMLimit}), .\Ki[6] (Ki[6]), 
            .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Kp[5] (Kp[5]), .\Kp[1] (Kp[1]), 
            .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .IntegralLimit({IntegralLimit}), 
            .VCC_net(VCC_net), .setpoint({setpoint}), .motor_state({motor_state}), 
            .duty({duty}), .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(271[16] 283[4])
    SB_LUT4 add_145_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n40393), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16769_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n47127), .I3(GND_net), .O(n30458));   // verilog/coms.v(127[12] 300[6])
    defparam i16769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5400));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16770_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n47127), .I3(GND_net), .O(n30459));   // verilog/coms.v(127[12] 300[6])
    defparam i16770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16771_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n47127), .I3(GND_net), .O(n30460));   // verilog/coms.v(127[12] 300[6])
    defparam i16771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n41626), .I0(n3012), 
            .I1(VCC_net), .CO(n41627));
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n48865), .I1(n1722), .I2(n48697), .I3(n36762), 
            .O(n48701));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfefc;
    SB_LUT4 unary_minus_10_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10), 
            .I3(n40481), .O(pwm_setpoint_23__N_191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5399));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n41625), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_17 (.CI(n40481), .I0(GND_net), .I1(n10), 
            .CO(n40482));
    SB_LUT4 unary_minus_10_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11), 
            .I3(n40480), .O(pwm_setpoint_23__N_191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n2717), .I1(n2718), .I2(n48647), .I3(n2719), 
            .O(n48653));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_CARRY add_145_14 (.CI(n40393), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n40394));
    SB_CARRY unary_minus_10_add_3_16 (.CI(n40480), .I0(GND_net), .I1(n11), 
            .CO(n40481));
    SB_LUT4 i16772_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n47127), .I3(GND_net), .O(n30461));   // verilog/coms.v(127[12] 300[6])
    defparam i16772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n40479), .O(pwm_setpoint_23__N_191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_15 (.CI(n40479), .I0(GND_net), .I1(n12), 
            .CO(n40480));
    SB_LUT4 unary_minus_10_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13), 
            .I3(n40478), .O(pwm_setpoint_23__N_191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_14 (.CI(n40478), .I0(GND_net), .I1(n13), 
            .CO(n40479));
    SB_LUT4 i16518_3_lut (.I0(current[6]), .I1(data_adj_5497[6]), .I2(n47264), 
            .I3(GND_net), .O(n30207));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16773_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n47127), .I3(GND_net), .O(n30462));   // verilog/coms.v(127[12] 300[6])
    defparam i16773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(n2715), .I1(n2716), .I2(n48653), .I3(n46644), 
            .O(n48659));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i36645_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n48701), 
            .O(n1752));
    defparam i36645_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5398));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n40477), .O(pwm_setpoint_23__N_191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16774_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n47127), .I3(GND_net), .O(n30463));   // verilog/coms.v(127[12] 300[6])
    defparam i16774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16775_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n47127), .I3(GND_net), .O(n30464));   // verilog/coms.v(127[12] 300[6])
    defparam i16775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16244_2_lut (.I0(n29588), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29939));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i16244_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n7066), 
            .D(n1103), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5397));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16776_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n47127), .I3(GND_net), .O(n30465));   // verilog/coms.v(127[12] 300[6])
    defparam i16776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36354_4_lut (.I0(commutation_state[1]), .I1(n25788), .I2(dti), 
            .I3(commutation_state[2]), .O(n29588));
    defparam i36354_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 mux_238_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16777_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n47127), .I3(GND_net), .O(n30466));   // verilog/coms.v(127[12] 300[6])
    defparam i16777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5396));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16778_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n47127), .I3(GND_net), .O(n30467));   // verilog/coms.v(127[12] 300[6])
    defparam i16778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16779_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n47127), .I3(GND_net), .O(n30468));   // verilog/coms.v(127[12] 300[6])
    defparam i16779_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_13 (.CI(n40477), .I0(GND_net), .I1(n14), 
            .CO(n40478));
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n41625), .I0(n3013), 
            .I1(VCC_net), .CO(n41626));
    SB_LUT4 mux_238_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_10_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5274), 
            .I3(n40476), .O(pwm_setpoint_23__N_191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5395));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n7066), 
            .D(n1104), .R(n29965));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n48659), 
            .O(n48665));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i16780_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n47127), .I3(GND_net), .O(n30469));   // verilog/coms.v(127[12] 300[6])
    defparam i16780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n1825), .I1(n1827), .I2(n1828), .I3(n1826), 
            .O(n48847));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hfffe;
    SB_LUT4 i16781_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n47127), .I3(GND_net), .O(n30470));   // verilog/coms.v(127[12] 300[6])
    defparam i16781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36901_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n48665), 
            .O(n2742));
    defparam i36901_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5394));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16782_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n47127), .I3(GND_net), .O(n30471));   // verilog/coms.v(127[12] 300[6])
    defparam i16782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n41624), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n41624), .I0(n3014), 
            .I1(VCC_net), .CO(n41625));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n41623), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_12 (.CI(n40476), .I0(GND_net), .I1(n15_adj_5274), 
            .CO(n40477));
    SB_LUT4 unary_minus_10_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16), 
            .I3(n40475), .O(pwm_setpoint_23__N_191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16783_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n47127), .I3(GND_net), .O(n30472));   // verilog/coms.v(127[12] 300[6])
    defparam i16783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n40435), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_11 (.CI(n40475), .I0(GND_net), .I1(n16), 
            .CO(n40476));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5393));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n41623), .I0(n3015), 
            .I1(VCC_net), .CO(n41624));
    SB_LUT4 add_224_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n40434), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16784_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n47127), .I3(GND_net), .O(n30473));   // verilog/coms.v(127[12] 300[6])
    defparam i16784_3_lut.LUT_INIT = 16'hacac;
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23073_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n36758));
    defparam i23073_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16785_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n47127), .I3(GND_net), .O(n30474));   // verilog/coms.v(127[12] 300[6])
    defparam i16785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1815 (.I0(n1823), .I1(n1824), .I2(n48847), .I3(GND_net), 
            .O(n48851));
    defparam i1_3_lut_adj_1815.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5392));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16786_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n47127), .I3(GND_net), .O(n30475));   // verilog/coms.v(127[12] 300[6])
    defparam i16786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16787_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n47127), .I3(GND_net), .O(n30476));   // verilog/coms.v(127[12] 300[6])
    defparam i16787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5391));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16788_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n47127), .I3(GND_net), .O(n30477));   // verilog/coms.v(127[12] 300[6])
    defparam i16788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16789_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n47127), .I3(GND_net), .O(n30478));   // verilog/coms.v(127[12] 300[6])
    defparam i16789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5390));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16790_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n47127), .I3(GND_net), .O(n30479));   // verilog/coms.v(127[12] 300[6])
    defparam i16790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16791_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n47127), .I3(GND_net), .O(n30480));   // verilog/coms.v(127[12] 300[6])
    defparam i16791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5389));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16792_3_lut (.I0(\data_out_frame[27] [1]), .I1(n47698), .I2(n29783), 
            .I3(GND_net), .O(n30481));   // verilog/coms.v(127[12] 300[6])
    defparam i16792_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i16793_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n25701), .I3(GND_net), .O(n30482));   // verilog/coms.v(127[12] 300[6])
    defparam i16793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n1829), .I1(n36758), .I2(n1830), .I3(n1831), 
            .O(n46621));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'ha080;
    SB_LUT4 i16794_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n25701), .I3(GND_net), .O(n30483));   // verilog/coms.v(127[12] 300[6])
    defparam i16794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16795_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n25701), .I3(GND_net), .O(n30484));   // verilog/coms.v(127[12] 300[6])
    defparam i16795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16796_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n25701), .I3(GND_net), .O(n30485));   // verilog/coms.v(127[12] 300[6])
    defparam i16796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16797_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n25701), .I3(GND_net), .O(n30486));   // verilog/coms.v(127[12] 300[6])
    defparam i16797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16798_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n25701), .I3(GND_net), .O(n30487));   // verilog/coms.v(127[12] 300[6])
    defparam i16798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n1821), .I1(n1822), .I2(n46621), .I3(n48851), 
            .O(n48857));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 i16799_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n25701), .I3(GND_net), .O(n30488));   // verilog/coms.v(127[12] 300[6])
    defparam i16799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16800_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n25701), .I3(GND_net), .O(n30489));   // verilog/coms.v(127[12] 300[6])
    defparam i16800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36666_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n48857), 
            .O(n1851));
    defparam i36666_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16801_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n25701), .I3(GND_net), .O(n30490));   // verilog/coms.v(127[12] 300[6])
    defparam i16801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16802_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n25701), .I3(GND_net), .O(n30491));   // verilog/coms.v(127[12] 300[6])
    defparam i16802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16803_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n25701), .I3(GND_net), .O(n30492));   // verilog/coms.v(127[12] 300[6])
    defparam i16803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16804_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n25701), .I3(GND_net), .O(n30493));   // verilog/coms.v(127[12] 300[6])
    defparam i16804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16805_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n25701), .I3(GND_net), .O(n30494));   // verilog/coms.v(127[12] 300[6])
    defparam i16805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16806_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n25701), .I3(GND_net), .O(n30495));   // verilog/coms.v(127[12] 300[6])
    defparam i16806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16807_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n25701), .I3(GND_net), .O(n30496));   // verilog/coms.v(127[12] 300[6])
    defparam i16807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16808_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n25701), .I3(GND_net), .O(n30497));   // verilog/coms.v(127[12] 300[6])
    defparam i16808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16809_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n25701), .I3(GND_net), .O(n30498));   // verilog/coms.v(127[12] 300[6])
    defparam i16809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1818 (.I0(n2824), .I1(n2820), .I2(n2821), .I3(GND_net), 
            .O(n49025));
    defparam i1_3_lut_adj_1818.LUT_INIT = 16'hfefe;
    SB_LUT4 i16810_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n25701), .I3(GND_net), .O(n30499));   // verilog/coms.v(127[12] 300[6])
    defparam i16810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16811_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n25701), .I3(GND_net), .O(n30500));   // verilog/coms.v(127[12] 300[6])
    defparam i16811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16813_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n25701), .I3(GND_net), .O(n30502));   // verilog/coms.v(127[12] 300[6])
    defparam i16813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16814_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n25701), .I3(GND_net), .O(n30503));   // verilog/coms.v(127[12] 300[6])
    defparam i16814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16815_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n25701), .I3(GND_net), .O(n30504));   // verilog/coms.v(127[12] 300[6])
    defparam i16815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n2826), .I1(n2825), .I2(n2823), .I3(n2828), 
            .O(n49027));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i16816_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n25701), .I3(GND_net), .O(n30505));   // verilog/coms.v(127[12] 300[6])
    defparam i16816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16818_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n25701), .I3(GND_net), .O(n30507));   // verilog/coms.v(127[12] 300[6])
    defparam i16818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16819_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n25701), .I3(GND_net), .O(n30508));   // verilog/coms.v(127[12] 300[6])
    defparam i16819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16820_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n25701), .I3(GND_net), .O(n30509));   // verilog/coms.v(127[12] 300[6])
    defparam i16820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16821_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n25701), .I3(GND_net), .O(n30510));   // verilog/coms.v(127[12] 300[6])
    defparam i16821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16822_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n25701), .I3(GND_net), .O(n30511));   // verilog/coms.v(127[12] 300[6])
    defparam i16822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16823_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n25701), .I3(GND_net), .O(n30512));   // verilog/coms.v(127[12] 300[6])
    defparam i16823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16824_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n25701), .I3(GND_net), .O(n30513));   // verilog/coms.v(127[12] 300[6])
    defparam i16824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16825_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n25701), .I3(GND_net), .O(n30514));   // verilog/coms.v(127[12] 300[6])
    defparam i16825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n49027), .I1(n49025), .I2(n2822), .I3(n2827), 
            .O(n49031));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'hfffe;
    SB_LUT4 i16826_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n25701), .I3(GND_net), .O(n30515));   // verilog/coms.v(127[12] 300[6])
    defparam i16826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16827_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[12]), 
            .I2(n25701), .I3(GND_net), .O(n30516));   // verilog/coms.v(127[12] 300[6])
    defparam i16827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16828_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n25701), .I3(GND_net), .O(n30517));   // verilog/coms.v(127[12] 300[6])
    defparam i16828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23071_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n36756));
    defparam i23071_3_lut.LUT_INIT = 16'hc8c8;
    \grp_debouncer(3,1000)  debounce (.reg_B({reg_B}), .CLK_c(CLK_c), .n48368(n48368), 
            .data_i({hall1, hall2, hall3}), .n30744(n30744), .data_o({h1, 
            h2, h3}), .n30743(n30743), .n30123(n30123), .GND_net(GND_net), 
            .VCC_net(VCC_net));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    SB_LUT4 i16829_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n25701), .I3(GND_net), .O(n30518));   // verilog/coms.v(127[12] 300[6])
    defparam i16829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16830_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n25701), .I3(GND_net), .O(n30519));   // verilog/coms.v(127[12] 300[6])
    defparam i16830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23135_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n36822));
    defparam i23135_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16831_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n25701), .I3(GND_net), .O(n30520));   // verilog/coms.v(127[12] 300[6])
    defparam i16831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16832_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n25701), .I3(GND_net), .O(n30521));   // verilog/coms.v(127[12] 300[6])
    defparam i16832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(n1929), .I1(n36756), .I2(n1930), .I3(n1931), 
            .O(n46606));
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n2817), .I1(n2818), .I2(n49031), .I3(n2819), 
            .O(n49037));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n1925), .I1(n1926), .I2(n1928), .I3(n1927), 
            .O(n48589));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i16833_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n25701), .I3(GND_net), .O(n30522));   // verilog/coms.v(127[12] 300[6])
    defparam i16833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16451_4_lut (.I0(CS_MISO_c), .I1(data_adj_5497[6]), .I2(n5_adj_5316), 
            .I3(n28440), .O(n30140));   // verilog/tli4970.v(33[10] 66[6])
    defparam i16451_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(n46606), .I1(n1921), .I2(n1923), .I3(n1924), 
            .O(n48789));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i16834_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n25701), .I3(GND_net), .O(n30523));   // verilog/coms.v(127[12] 300[6])
    defparam i16834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16836_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n25701), .I3(GND_net), .O(n30525));   // verilog/coms.v(127[12] 300[6])
    defparam i16836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n28264), .I3(n1195), .O(n7264));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i16837_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n25701), .I3(GND_net), .O(n30526));   // verilog/coms.v(127[12] 300[6])
    defparam i16837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n28264), .I3(GND_net), .O(n28265));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i22019_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n28264), .I3(n1195), .O(n35695));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i22019_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n49037), .I1(n2829), .I2(n36822), .I3(n2830), 
            .O(n49039));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1826 (.I0(n1918), .I1(n1920), .I2(n1922), .I3(n48589), 
            .O(n48595));
    defparam i1_4_lut_adj_1826.LUT_INIT = 16'hfffe;
    SB_LUT4 i16838_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n25701), .I3(GND_net), .O(n30527));   // verilog/coms.v(127[12] 300[6])
    defparam i16838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16839_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n25701), .I3(GND_net), .O(n30528));   // verilog/coms.v(127[12] 300[6])
    defparam i16839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n28264), .I3(GND_net), .O(n7066));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 mux_238_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n49039), 
            .O(n49045));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 i16840_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n25701), .I3(GND_net), .O(n30529));   // verilog/coms.v(127[12] 300[6])
    defparam i16840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16841_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n25701), .I3(GND_net), .O(n30530));   // verilog/coms.v(127[12] 300[6])
    defparam i16841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16842_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n25701), .I3(GND_net), .O(n30531));   // verilog/coms.v(127[12] 300[6])
    defparam i16842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16843_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n25701), .I3(GND_net), .O(n30532));   // verilog/coms.v(127[12] 300[6])
    defparam i16843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16844_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n25701), .I3(GND_net), .O(n30533));   // verilog/coms.v(127[12] 300[6])
    defparam i16844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16845_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n25701), .I3(GND_net), .O(n30534));   // verilog/coms.v(127[12] 300[6])
    defparam i16845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16846_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n25701), .I3(GND_net), .O(n30535));   // verilog/coms.v(127[12] 300[6])
    defparam i16846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5312));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5313));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_279));   // verilog/TinyFPGA_B.v(321[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i16847_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n25701), .I3(GND_net), .O(n30536));   // verilog/coms.v(127[12] 300[6])
    defparam i16847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16848_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n25701), .I3(GND_net), .O(n30537));   // verilog/coms.v(127[12] 300[6])
    defparam i16848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36688_4_lut (.I0(n48595), .I1(n1917), .I2(n48789), .I3(n1919), 
            .O(n1950));
    defparam i36688_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n49045), 
            .O(n49051));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i23067_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n36752));
    defparam i23067_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16849_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n25701), .I3(GND_net), .O(n30538));   // verilog/coms.v(127[12] 300[6])
    defparam i16849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16850_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n25701), .I3(GND_net), .O(n30539));   // verilog/coms.v(127[12] 300[6])
    defparam i16850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16851_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n25701), .I3(GND_net), .O(n30540));   // verilog/coms.v(127[12] 300[6])
    defparam i16851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16852_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n25701), .I3(GND_net), .O(n30541));   // verilog/coms.v(127[12] 300[6])
    defparam i16852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36934_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n49051), 
            .O(n2841));
    defparam i36934_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16853_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n25701), .I3(GND_net), .O(n30542));   // verilog/coms.v(127[12] 300[6])
    defparam i16853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16854_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n25701), .I3(GND_net), .O(n30543));   // verilog/coms.v(127[12] 300[6])
    defparam i16854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1829 (.I0(n2027), .I1(n2026), .I2(GND_net), .I3(GND_net), 
            .O(n48875));
    defparam i1_2_lut_adj_1829.LUT_INIT = 16'heeee;
    SB_LUT4 i16855_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n25701), .I3(GND_net), .O(n30544));   // verilog/coms.v(127[12] 300[6])
    defparam i16855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16856_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n25701), 
            .I3(GND_net), .O(n30545));   // verilog/coms.v(127[12] 300[6])
    defparam i16856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16857_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n25701), 
            .I3(GND_net), .O(n30546));   // verilog/coms.v(127[12] 300[6])
    defparam i16857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16858_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n25701), 
            .I3(GND_net), .O(n30547));   // verilog/coms.v(127[12] 300[6])
    defparam i16858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16859_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n25701), 
            .I3(GND_net), .O(n30548));   // verilog/coms.v(127[12] 300[6])
    defparam i16859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16860_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n25701), 
            .I3(GND_net), .O(n30549));   // verilog/coms.v(127[12] 300[6])
    defparam i16860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16861_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n25701), 
            .I3(GND_net), .O(n30550));   // verilog/coms.v(127[12] 300[6])
    defparam i16861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut_4_lut (.I0(n2_adj_5362), 
            .I1(encoder0_position[31]), .I2(n48899), .I3(n7607), .O(n828));
    defparam encoder0_position_31__I_0_i500_4_lut_4_lut.LUT_INIT = 16'ha808;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2025_adj_5377), .I1(n48875), .I2(n2024), 
            .I3(n2028), .O(n48879));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    SB_LUT4 i16862_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n25701), 
            .I3(GND_net), .O(n30551));   // verilog/coms.v(127[12] 300[6])
    defparam i16862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16863_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n25701), 
            .I3(GND_net), .O(n30552));   // verilog/coms.v(127[12] 300[6])
    defparam i16863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16864_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n25701), 
            .I3(GND_net), .O(n30553));   // verilog/coms.v(127[12] 300[6])
    defparam i16864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16865_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n25701), 
            .I3(GND_net), .O(n30554));   // verilog/coms.v(127[12] 300[6])
    defparam i16865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16866_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n25701), 
            .I3(GND_net), .O(n30555));   // verilog/coms.v(127[12] 300[6])
    defparam i16866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16867_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n25701), 
            .I3(GND_net), .O(n30556));   // verilog/coms.v(127[12] 300[6])
    defparam i16867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n2029), .I1(n36752), .I2(n2030), .I3(n2031), 
            .O(n46642));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'ha080;
    SB_LUT4 i16868_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n25701), 
            .I3(GND_net), .O(n30557));   // verilog/coms.v(127[12] 300[6])
    defparam i16868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16869_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n25701), 
            .I3(GND_net), .O(n30558));   // verilog/coms.v(127[12] 300[6])
    defparam i16869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16870_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n25701), 
            .I3(GND_net), .O(n30559));   // verilog/coms.v(127[12] 300[6])
    defparam i16870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n48879), 
            .O(n48885));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i16871_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n25701), 
            .I3(GND_net), .O(n30560));   // verilog/coms.v(127[12] 300[6])
    defparam i16871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16872_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n25701), 
            .I3(GND_net), .O(n30561));   // verilog/coms.v(127[12] 300[6])
    defparam i16872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16873_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n25701), 
            .I3(GND_net), .O(n30562));   // verilog/coms.v(127[12] 300[6])
    defparam i16873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16874_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n25701), 
            .I3(GND_net), .O(n30563));   // verilog/coms.v(127[12] 300[6])
    defparam i16874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16875_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n25701), 
            .I3(GND_net), .O(n30564));   // verilog/coms.v(127[12] 300[6])
    defparam i16875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16876_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n25701), 
            .I3(GND_net), .O(n30565));   // verilog/coms.v(127[12] 300[6])
    defparam i16876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16877_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n25701), 
            .I3(GND_net), .O(n30566));   // verilog/coms.v(127[12] 300[6])
    defparam i16877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16878_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n25701), 
            .I3(GND_net), .O(n30567));   // verilog/coms.v(127[12] 300[6])
    defparam i16878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16879_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n25701), 
            .I3(GND_net), .O(n30568));   // verilog/coms.v(127[12] 300[6])
    defparam i16879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16880_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n25701), .I3(GND_net), .O(n30569));   // verilog/coms.v(127[12] 300[6])
    defparam i16880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16881_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n25701), .I3(GND_net), .O(n30570));   // verilog/coms.v(127[12] 300[6])
    defparam i16881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16882_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n25701), .I3(GND_net), .O(n30571));   // verilog/coms.v(127[12] 300[6])
    defparam i16882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16883_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n25701), .I3(GND_net), .O(n30572));   // verilog/coms.v(127[12] 300[6])
    defparam i16883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n2019), .I1(n2020), .I2(n48885), .I3(n46642), 
            .O(n48891));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i16884_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n25701), .I3(GND_net), .O(n30573));   // verilog/coms.v(127[12] 300[6])
    defparam i16884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16885_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n25701), .I3(GND_net), .O(n30574));   // verilog/coms.v(127[12] 300[6])
    defparam i16885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16886_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n25701), .I3(GND_net), .O(n30575));   // verilog/coms.v(127[12] 300[6])
    defparam i16886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16887_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n25701), .I3(GND_net), .O(n30576));   // verilog/coms.v(127[12] 300[6])
    defparam i16887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16888_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n25701), .I3(GND_net), .O(n30577));   // verilog/coms.v(127[12] 300[6])
    defparam i16888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16889_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n25701), .I3(GND_net), .O(n30578));   // verilog/coms.v(127[12] 300[6])
    defparam i16889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16890_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n25701), .I3(GND_net), .O(n30579));   // verilog/coms.v(127[12] 300[6])
    defparam i16890_3_lut.LUT_INIT = 16'hcaca;
    EEPROM eeprom (.\state[3] (state_adj_5517[3]), .n6(n6_adj_5292), .GND_net(GND_net), 
           .CLK_c(CLK_c), .n5608({n5609}), .\state[1] (state_adj_5493[1]), 
           .read(read), .\state[0] (state_adj_5493[0]), .enable_slow_N_4190(enable_slow_N_4190), 
           .\state[1]_adj_18 (state_adj_5517[1]), .\state[2] (state_adj_5517[2]), 
           .n7(n7_adj_5283), .n30170(n30170), .rw(rw), .n45294(n45294), 
           .data_ready(data_ready), .n45186(n45186), .n45170(n45170), 
           .n36514(n36514), .n46391(n46391), .n45666(n45666), .\state_7__N_4087[0] (state_7__N_4087[0]), 
           .sda_enable(sda_enable), .n4(n4_adj_5350), .scl_enable_N_4177(scl_enable_N_4177), 
           .scl_enable(scl_enable), .n6686(n6686), .n35782(n35782), .n8(n8_adj_5384), 
           .VCC_net(VCC_net), .\state[0]_adj_19 (state_adj_5517[0]), .n4_adj_20(n4_adj_5272), 
           .\saved_addr[0] (saved_addr[0]), .n6496(n6496), .n51120(n51120), 
           .n15(n15), .n10(n10_adj_5321), .n28421(n28421), .n28416(n28416), 
           .n10_adj_21(n10_adj_5431), .\state_7__N_4103[3] (state_7__N_4103[3]), 
           .n7227(n7227), .n30174(n30174), .n30159(n30159), .data({data}), 
           .n30158(n30158), .n30157(n30157), .n30146(n30146), .scl(scl), 
           .sda_out(sda_out), .n30138(n30138), .n30137(n30137), .n30136(n30136), 
           .n30135(n30135), .n10_adj_22(n10_adj_5364)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(387[10] 398[6])
    SB_LUT4 i16891_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n25701), .I3(GND_net), .O(n30580));   // verilog/coms.v(127[12] 300[6])
    defparam i16891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16892_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n25701), .I3(GND_net), .O(n30581));   // verilog/coms.v(127[12] 300[6])
    defparam i16892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16893_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n25701), .I3(GND_net), .O(n30582));   // verilog/coms.v(127[12] 300[6])
    defparam i16893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16894_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n25701), .I3(GND_net), .O(n30583));   // verilog/coms.v(127[12] 300[6])
    defparam i16894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16895_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n25701), .I3(GND_net), .O(n30584));   // verilog/coms.v(127[12] 300[6])
    defparam i16895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16896_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n25701), .I3(GND_net), .O(n30585));   // verilog/coms.v(127[12] 300[6])
    defparam i16896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16897_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n25701), .I3(GND_net), .O(n30586));   // verilog/coms.v(127[12] 300[6])
    defparam i16897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16898_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n25701), .I3(GND_net), .O(n30587));   // verilog/coms.v(127[12] 300[6])
    defparam i16898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16899_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n25701), .I3(GND_net), .O(n30588));   // verilog/coms.v(127[12] 300[6])
    defparam i16899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16900_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n25701), .I3(GND_net), .O(n30589));   // verilog/coms.v(127[12] 300[6])
    defparam i16900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16901_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n25701), .I3(GND_net), .O(n30590));   // verilog/coms.v(127[12] 300[6])
    defparam i16901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16902_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n25701), .I3(GND_net), .O(n30591));   // verilog/coms.v(127[12] 300[6])
    defparam i16902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16903_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n25701), .I3(GND_net), .O(n30592));   // verilog/coms.v(127[12] 300[6])
    defparam i16903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16904_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n25701), .I3(GND_net), .O(n30593));   // verilog/coms.v(127[12] 300[6])
    defparam i16904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16905_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n25701), .I3(GND_net), .O(n30594));   // verilog/coms.v(127[12] 300[6])
    defparam i16905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16906_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n25701), .I3(GND_net), .O(n30595));   // verilog/coms.v(127[12] 300[6])
    defparam i16906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16907_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n25701), .I3(GND_net), .O(n30596));   // verilog/coms.v(127[12] 300[6])
    defparam i16907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16908_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n25701), .I3(GND_net), .O(n30597));   // verilog/coms.v(127[12] 300[6])
    defparam i16908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16909_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n25701), .I3(GND_net), .O(n30598));   // verilog/coms.v(127[12] 300[6])
    defparam i16909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16910_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n25701), .I3(GND_net), .O(n30599));   // verilog/coms.v(127[12] 300[6])
    defparam i16910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n29660), 
            .I3(rx_data_ready), .O(n45162));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i16911_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n25701), .I3(GND_net), .O(n30600));   // verilog/coms.v(127[12] 300[6])
    defparam i16911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16912_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n25701), .I3(GND_net), .O(n30601));   // verilog/coms.v(127[12] 300[6])
    defparam i16912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16913_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n25701), .I3(GND_net), .O(n30602));   // verilog/coms.v(127[12] 300[6])
    defparam i16913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16914_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n25701), .I3(GND_net), .O(n30603));   // verilog/coms.v(127[12] 300[6])
    defparam i16914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16915_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n25701), .I3(GND_net), .O(n30604));   // verilog/coms.v(127[12] 300[6])
    defparam i16915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16916_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n25701), .I3(GND_net), .O(n30605));   // verilog/coms.v(127[12] 300[6])
    defparam i16916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16917_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n25701), .I3(GND_net), .O(n30606));   // verilog/coms.v(127[12] 300[6])
    defparam i16917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16918_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n25701), .I3(GND_net), .O(n30607));   // verilog/coms.v(127[12] 300[6])
    defparam i16918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16919_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n25701), .I3(GND_net), .O(n30608));   // verilog/coms.v(127[12] 300[6])
    defparam i16919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16920_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n25701), .I3(GND_net), .O(n30609));   // verilog/coms.v(127[12] 300[6])
    defparam i16920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16921_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n25701), .I3(GND_net), .O(n30610));   // verilog/coms.v(127[12] 300[6])
    defparam i16921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16922_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n25701), .I3(GND_net), .O(n30611));   // verilog/coms.v(127[12] 300[6])
    defparam i16922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16923_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n25701), .I3(GND_net), .O(n30612));   // verilog/coms.v(127[12] 300[6])
    defparam i16923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16924_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n25701), .I3(GND_net), .O(n30613));   // verilog/coms.v(127[12] 300[6])
    defparam i16924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16925_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n25701), .I3(GND_net), .O(n30614));   // verilog/coms.v(127[12] 300[6])
    defparam i16925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16926_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n25701), .I3(GND_net), .O(n30615));   // verilog/coms.v(127[12] 300[6])
    defparam i16926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16927_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n25701), .I3(GND_net), .O(n30616));   // verilog/coms.v(127[12] 300[6])
    defparam i16927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16928_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n25701), .I3(GND_net), .O(n30617));   // verilog/coms.v(127[12] 300[6])
    defparam i16928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16929_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n25701), .I3(GND_net), .O(n30618));   // verilog/coms.v(127[12] 300[6])
    defparam i16929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16930_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n25701), .I3(GND_net), .O(n30619));   // verilog/coms.v(127[12] 300[6])
    defparam i16930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16931_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n25701), .I3(GND_net), .O(n30620));   // verilog/coms.v(127[12] 300[6])
    defparam i16931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16932_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n25701), .I3(GND_net), .O(n30621));   // verilog/coms.v(127[12] 300[6])
    defparam i16932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16933_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n25701), .I3(GND_net), .O(n30622));   // verilog/coms.v(127[12] 300[6])
    defparam i16933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16934_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n25701), .I3(GND_net), .O(n30623));   // verilog/coms.v(127[12] 300[6])
    defparam i16934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5517[0]), .I1(n51120), .I2(n6686), 
            .I3(n10_adj_5321), .O(n8_adj_5384));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 i16935_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n25701), .I3(GND_net), .O(n30624));   // verilog/coms.v(127[12] 300[6])
    defparam i16935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16936_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n25701), .I3(GND_net), .O(n30625));   // verilog/coms.v(127[12] 300[6])
    defparam i16936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16937_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n25701), .I3(GND_net), .O(n30626));   // verilog/coms.v(127[12] 300[6])
    defparam i16937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16938_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n25701), .I3(GND_net), .O(n30627));   // verilog/coms.v(127[12] 300[6])
    defparam i16938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5273));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16939_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n25701), .I3(GND_net), .O(n30628));   // verilog/coms.v(127[12] 300[6])
    defparam i16939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16940_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n25701), .I3(GND_net), .O(n30629));   // verilog/coms.v(127[12] 300[6])
    defparam i16940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16941_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n25701), .I3(GND_net), .O(n30630));   // verilog/coms.v(127[12] 300[6])
    defparam i16941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16942_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n25701), .I3(GND_net), .O(n30631));   // verilog/coms.v(127[12] 300[6])
    defparam i16942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16943_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n25701), .I3(GND_net), .O(n30632));   // verilog/coms.v(127[12] 300[6])
    defparam i16943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16944_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n25701), .I3(GND_net), .O(n30633));   // verilog/coms.v(127[12] 300[6])
    defparam i16944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5506[1]), .I1(r_SM_Main_adj_5506[0]), 
            .I2(r_SM_Main_adj_5506[2]), .I3(r_SM_Main_2__N_3613[1]), .O(n53023));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_4_lut_adj_1834 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main_2__N_3542[2]), .O(n45602));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_4_lut_adj_1834.LUT_INIT = 16'h2000;
    TLI4970 tli (.\data[15] (data_adj_5497[15]), .\state[1] (state_adj_5499[1]), 
            .\state[0] (state_adj_5499[0]), .n47264(n47264), .GND_net(GND_net), 
            .n6(n6_adj_5317), .n15(n15_adj_5325), .n5(n5_adj_5315), .n5_adj_13(n5_adj_5316), 
            .n35840(n35840), .CLK_c(CLK_c), .n30212(n30212), .current({current}), 
            .n30211(n30211), .n30210(n30210), .n30209(n30209), .n30208(n30208), 
            .n30207(n30207), .n30206(n30206), .n30205(n30205), .n30204(n30204), 
            .n30203(n30203), .n30202(n30202), .n30201(n30201), .n30198(n30198), 
            .\data[0] (data_adj_5497[0]), .n10(n10_adj_5345), .n9(n9_adj_5344), 
            .n11(n11_adj_5346), .state_7__N_4293(state_7__N_4293), .n9_adj_14(n9_adj_5387), 
            .clk_out(clk_out), .n30171(n30171), .CS_c(CS_c), .n30168(n30168), 
            .n30148(n30148), .n30147(n30147), .\data[12] (data_adj_5497[12]), 
            .n30145(n30145), .\data[11] (data_adj_5497[11]), .n30144(n30144), 
            .\data[10] (data_adj_5497[10]), .n30143(n30143), .\data[9] (data_adj_5497[9]), 
            .n28429(n28429), .n28432(n28432), .n30142(n30142), .\data[8] (data_adj_5497[8]), 
            .n30141(n30141), .\data[7] (data_adj_5497[7]), .n28437(n28437), 
            .n30140(n30140), .\data[6] (data_adj_5497[6]), .n30139(n30139), 
            .\data[5] (data_adj_5497[5]), .n30134(n30134), .\data[4] (data_adj_5497[4]), 
            .n30133(n30133), .\data[3] (data_adj_5497[3]), .n30132(n30132), 
            .\data[2] (data_adj_5497[2]), .n30131(n30131), .\data[1] (data_adj_5497[1]), 
            .n28444(n28444), .VCC_net(VCC_net), .CS_CLK_c(CS_CLK_c), .n28440(n28440)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(400[11] 406[4])
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.b_prev(b_prev), .GND_net(GND_net), 
            .a_new({a_new[1], Open_0}), .direction_N_3907(direction_N_3907), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1668(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .n30218(n30218), .n1632(n1632), .encoder0_position({encoder0_position}), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(285[57] 292[6])
    SB_LUT4 i16945_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n25701), .I3(GND_net), .O(n30634));   // verilog/coms.v(127[12] 300[6])
    defparam i16945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36711_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n48891), 
            .O(n2049));
    defparam i36711_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16946_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n25701), .I3(GND_net), .O(n30635));   // verilog/coms.v(127[12] 300[6])
    defparam i16946_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i16947_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n25701), .I3(GND_net), .O(n30636));   // verilog/coms.v(127[12] 300[6])
    defparam i16947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16948_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n25701), .I3(GND_net), .O(n30637));   // verilog/coms.v(127[12] 300[6])
    defparam i16948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35865_3_lut_4_lut (.I0(n2841), .I1(n2742), .I2(n2726), .I3(n50080), 
            .O(n2924));
    defparam i35865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16530_3_lut_4_lut (.I0(n1673), .I1(b_prev_adj_5323), .I2(a_new_adj_5469[1]), 
            .I3(direction_N_3907_adj_5324), .O(n30219));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16530_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i16949_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n25701), .I3(GND_net), .O(n30638));   // verilog/coms.v(127[12] 300[6])
    defparam i16949_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(1,500000)  quad_counter1 (.b_prev(b_prev_adj_5323), 
            .GND_net(GND_net), .a_new({a_new_adj_5469[1], Open_1}), .direction_N_3907(direction_N_3907_adj_5324), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1668(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .n30219(n30219), .n1673(n1673), .encoder1_position({encoder1_position}), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(294[57] 301[6])
    SB_LUT4 i16529_3_lut_4_lut (.I0(n1632), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3907), .O(n30218));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16529_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i16950_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n25701), .I3(GND_net), .O(n30639));   // verilog/coms.v(127[12] 300[6])
    defparam i16950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16951_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n25701), .I3(GND_net), .O(n30640));   // verilog/coms.v(127[12] 300[6])
    defparam i16951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16952_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n25701), .I3(GND_net), .O(n30641));   // verilog/coms.v(127[12] 300[6])
    defparam i16952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16953_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n25701), .I3(GND_net), .O(n30642));   // verilog/coms.v(127[12] 300[6])
    defparam i16953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23065_3_lut (.I0(n946), .I1(n2132), .I2(n2133), .I3(GND_net), 
            .O(n36750));
    defparam i23065_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i16954_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n25701), .I3(GND_net), .O(n30643));   // verilog/coms.v(127[12] 300[6])
    defparam i16954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16955_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n25701), .I3(GND_net), .O(n30644));   // verilog/coms.v(127[12] 300[6])
    defparam i16955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16956_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n25701), .I3(GND_net), .O(n30645));   // verilog/coms.v(127[12] 300[6])
    defparam i16956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16957_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n25701), .I3(GND_net), .O(n30646));   // verilog/coms.v(127[12] 300[6])
    defparam i16957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16958_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n25701), .I3(GND_net), .O(n30647));   // verilog/coms.v(127[12] 300[6])
    defparam i16958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16959_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n25701), .I3(GND_net), .O(n30648));   // verilog/coms.v(127[12] 300[6])
    defparam i16959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16960_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n25701), 
            .I3(GND_net), .O(n30649));   // verilog/coms.v(127[12] 300[6])
    defparam i16960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16961_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n25701), 
            .I3(GND_net), .O(n30650));   // verilog/coms.v(127[12] 300[6])
    defparam i16961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16962_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n25701), 
            .I3(GND_net), .O(n30651));   // verilog/coms.v(127[12] 300[6])
    defparam i16962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16963_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n25701), 
            .I3(GND_net), .O(n30652));   // verilog/coms.v(127[12] 300[6])
    defparam i16963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16964_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n25701), 
            .I3(GND_net), .O(n30653));   // verilog/coms.v(127[12] 300[6])
    defparam i16964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16965_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n25701), 
            .I3(GND_net), .O(n30654));   // verilog/coms.v(127[12] 300[6])
    defparam i16965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16966_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n25701), 
            .I3(GND_net), .O(n30655));   // verilog/coms.v(127[12] 300[6])
    defparam i16966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16967_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n25701), 
            .I3(GND_net), .O(n30656));   // verilog/coms.v(127[12] 300[6])
    defparam i16967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16968_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n29618), 
            .I3(GND_net), .O(n30657));   // verilog/coms.v(127[12] 300[6])
    defparam i16968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16969_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n29618), 
            .I3(GND_net), .O(n30658));   // verilog/coms.v(127[12] 300[6])
    defparam i16969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16970_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n29618), 
            .I3(GND_net), .O(n30659));   // verilog/coms.v(127[12] 300[6])
    defparam i16970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16971_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n29618), 
            .I3(GND_net), .O(n30660));   // verilog/coms.v(127[12] 300[6])
    defparam i16971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16972_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n29618), 
            .I3(GND_net), .O(n30661));   // verilog/coms.v(127[12] 300[6])
    defparam i16972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16973_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n29618), 
            .I3(GND_net), .O(n30662));   // verilog/coms.v(127[12] 300[6])
    defparam i16973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16974_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n29618), 
            .I3(GND_net), .O(n30663));   // verilog/coms.v(127[12] 300[6])
    defparam i16974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5287), .I3(n15_adj_5341), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16975_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n29618), 
            .I3(GND_net), .O(n30664));   // verilog/coms.v(127[12] 300[6])
    defparam i16975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16976_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n29618), 
            .I3(GND_net), .O(n30665));   // verilog/coms.v(127[12] 300[6])
    defparam i16976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16977_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n29618), 
            .I3(GND_net), .O(n30666));   // verilog/coms.v(127[12] 300[6])
    defparam i16977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16978_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n29618), 
            .I3(GND_net), .O(n30667));   // verilog/coms.v(127[12] 300[6])
    defparam i16978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16979_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n29618), 
            .I3(GND_net), .O(n30668));   // verilog/coms.v(127[12] 300[6])
    defparam i16979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16980_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n29618), 
            .I3(GND_net), .O(n30669));   // verilog/coms.v(127[12] 300[6])
    defparam i16980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16981_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n29618), 
            .I3(GND_net), .O(n30670));   // verilog/coms.v(127[12] 300[6])
    defparam i16981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16982_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n29618), 
            .I3(GND_net), .O(n30671));   // verilog/coms.v(127[12] 300[6])
    defparam i16982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16500_4_lut (.I0(n29701), .I1(r_Bit_Index[0]), .I2(n45507), 
            .I3(r_SM_Main[1]), .O(n30189));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16500_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i1_4_lut_adj_1835 (.I0(n2125), .I1(n2127), .I2(n2128), .I3(n2126), 
            .O(n48805));
    defparam i1_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 i16984_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n29618), 
            .I3(GND_net), .O(n30673));   // verilog/coms.v(127[12] 300[6])
    defparam i16984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16985_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n29618), 
            .I3(GND_net), .O(n30674));   // verilog/coms.v(127[12] 300[6])
    defparam i16985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n2129), .I1(n36750), .I2(n2130), .I3(n2131), 
            .O(n46623));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'ha080;
    SB_LUT4 i16986_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n29618), 
            .I3(GND_net), .O(n30675));   // verilog/coms.v(127[12] 300[6])
    defparam i16986_3_lut.LUT_INIT = 16'hcaca;
    coms neopxl_color_23__I_0 (.n30269(n30269), .PWMLimit({PWMLimit}), .CLK_c(CLK_c), 
         .n30268(n30268), .n30267(n30267), .n30266(n30266), .n30265(n30265), 
         .n30264(n30264), .GND_net(GND_net), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\FRAME_MATCHER.state ({Open_2, 
         Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, Open_9, 
         Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, Open_16, 
         Open_17, Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
         Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, Open_30, 
         Open_31, Open_32, \FRAME_MATCHER.state [0]}), .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .n30263(n30263), 
         .n30262(n30262), .n30261(n30261), .rx_data_ready(rx_data_ready), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .n30260(n30260), .n30259(n30259), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n30258(n30258), 
         .\data_out_frame[20] ({\data_out_frame[20] [7:5], Open_33, \data_out_frame[20] [3:2], 
         Open_34, Open_35}), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), .\data_in[3] ({\data_in[3] }), 
         .\data_in[2] ({\data_in[2] }), .n771(n771), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .n4452(n4452), .n28383(n28383), .n63(n63), .n3807(n3807), .setpoint({setpoint}), 
         .n30257(n30257), .n63_adj_3(n63_adj_5380), .n3303(n3303), .n122(n122), 
         .n42261(n42261), .n5(n5_adj_5381), .n53135(n53135), .n30256(n30256), 
         .n30255(n30255), .n30254(n30254), .n30253(n30253), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .n52967(n52967), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .tx_transmit_N_3513(tx_transmit_N_3513), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[21][4] (\data_out_frame[21] [4]), 
         .\data_out_frame[20][1] (\data_out_frame[20] [1]), .\data_out_frame[21][1] (\data_out_frame[21] [1]), 
         .\data_out_frame[21][2] (\data_out_frame[21] [2]), .ID({ID}), .DE_c(DE_c), 
         .LED_c(LED_c), .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n47698(n47698), .\data_out_frame[21][0] (\data_out_frame[21] [0]), 
         .\data_out_frame[27][1] (\data_out_frame[27] [1]), .n29783(n29783), 
         .\data_out_frame[20][0] (\data_out_frame[20] [0]), .\data_out_frame[21][3] (\data_out_frame[21] [3]), 
         .n25438(n25438), .n42259(n42259), .rx_data({rx_data}), .tx_active(tx_active), 
         .n2025(n2025), .n54(n54), .n46(n46), .n46338(n46338), .\state[2] (state_adj_5517[2]), 
         .\state[3] (state_adj_5517[3]), .n10(n10_adj_5364), .n44944(n44944), 
         .n30166(n30166), .n30165(n30165), .control_mode({control_mode}), 
         .n30163(n30163), .neopxl_color({neopxl_color}), .n30162(n30162), 
         .\Ki[0] (Ki[0]), .n30161(n30161), .\Kp[0] (Kp[0]), .n30160(n30160), 
         .n30742(n30742), .IntegralLimit({IntegralLimit}), .n30741(n30741), 
         .n30740(n30740), .n30739(n30739), .n30738(n30738), .n30737(n30737), 
         .n30736(n30736), .n30735(n30735), .n30734(n30734), .n30733(n30733), 
         .n30732(n30732), .n30731(n30731), .\state[0] (state_adj_5517[0]), 
         .\state[1] (state_adj_5517[1]), .enable_slow_N_4190(enable_slow_N_4190), 
         .n7227(n7227), .n30730(n30730), .n30729(n30729), .n30728(n30728), 
         .n30727(n30727), .n30726(n30726), .n30725(n30725), .n30724(n30724), 
         .n30723(n30723), .n30722(n30722), .n30721(n30721), .n30719(n30719), 
         .n30718(n30718), .n30717(n30717), .n30716(n30716), .n30715(n30715), 
         .n30714(n30714), .n30713(n30713), .n30712(n30712), .n30711(n30711), 
         .n30710(n30710), .n30709(n30709), .n30708(n30708), .n30707(n30707), 
         .n30706(n30706), .n30705(n30705), .n30704(n30704), .n30703(n30703), 
         .n30702(n30702), .n30701(n30701), .n30700(n30700), .n30699(n30699), 
         .n30698(n30698), .n30697(n30697), .n30696(n30696), .n30695(n30695), 
         .n30694(n30694), .n30693(n30693), .n30692(n30692), .n30691(n30691), 
         .n30690(n30690), .n30689(n30689), .n30688(n30688), .n30687(n30687), 
         .\Kp[1] (Kp[1]), .n30686(n30686), .\Kp[2] (Kp[2]), .n30685(n30685), 
         .\Kp[3] (Kp[3]), .n30684(n30684), .\Kp[4] (Kp[4]), .n30683(n30683), 
         .\Kp[5] (Kp[5]), .n30682(n30682), .\Kp[6] (Kp[6]), .n30681(n30681), 
         .\Kp[7] (Kp[7]), .n30680(n30680), .\Kp[8] (Kp[8]), .n30679(n30679), 
         .\Kp[9] (Kp[9]), .n30678(n30678), .\Kp[10] (Kp[10]), .n30677(n30677), 
         .\Kp[11] (Kp[11]), .n30676(n30676), .\Kp[12] (Kp[12]), .n30675(n30675), 
         .\Kp[13] (Kp[13]), .n30674(n30674), .\Kp[14] (Kp[14]), .n30673(n30673), 
         .\Kp[15] (Kp[15]), .n30671(n30671), .\Ki[1] (Ki[1]), .n30670(n30670), 
         .\Ki[2] (Ki[2]), .n30669(n30669), .\Ki[3] (Ki[3]), .n30668(n30668), 
         .\Ki[4] (Ki[4]), .n30667(n30667), .\Ki[5] (Ki[5]), .n30666(n30666), 
         .\Ki[6] (Ki[6]), .n30665(n30665), .\Ki[7] (Ki[7]), .n30664(n30664), 
         .\Ki[8] (Ki[8]), .n30663(n30663), .\Ki[9] (Ki[9]), .n30662(n30662), 
         .\Ki[10] (Ki[10]), .n30661(n30661), .\Ki[11] (Ki[11]), .n30660(n30660), 
         .\Ki[12] (Ki[12]), .n30659(n30659), .\Ki[13] (Ki[13]), .n30658(n30658), 
         .\Ki[14] (Ki[14]), .n30657(n30657), .\Ki[15] (Ki[15]), .n30656(n30656), 
         .n30655(n30655), .n30654(n30654), .n30653(n30653), .n30652(n30652), 
         .n30651(n30651), .n30650(n30650), .n30649(n30649), .n30648(n30648), 
         .n30647(n30647), .n30646(n30646), .n30645(n30645), .n30644(n30644), 
         .n30643(n30643), .n30642(n30642), .n30641(n30641), .n30640(n30640), 
         .n30639(n30639), .n30638(n30638), .n30637(n30637), .n30636(n30636), 
         .n30635(n30635), .n30634(n30634), .n30633(n30633), .n30632(n30632), 
         .n30631(n30631), .n30630(n30630), .n30629(n30629), .n30628(n30628), 
         .n30627(n30627), .n30626(n30626), .n30625(n30625), .n30624(n30624), 
         .n30623(n30623), .n30622(n30622), .n30621(n30621), .n30620(n30620), 
         .n30619(n30619), .n30618(n30618), .n30617(n30617), .n30616(n30616), 
         .n30615(n30615), .n30614(n30614), .n30613(n30613), .n30612(n30612), 
         .n30611(n30611), .n30610(n30610), .n30609(n30609), .n30608(n30608), 
         .n30607(n30607), .n30606(n30606), .n30605(n30605), .n30604(n30604), 
         .n30603(n30603), .n30602(n30602), .n30601(n30601), .n30600(n30600), 
         .n30599(n30599), .n30598(n30598), .n30597(n30597), .n30596(n30596), 
         .n30595(n30595), .n30594(n30594), .n30593(n30593), .n30592(n30592), 
         .n30591(n30591), .n30590(n30590), .n30589(n30589), .n30588(n30588), 
         .n30587(n30587), .n30586(n30586), .n30585(n30585), .n30584(n30584), 
         .n30583(n30583), .n30582(n30582), .n30581(n30581), .n30580(n30580), 
         .n30579(n30579), .n30578(n30578), .n30577(n30577), .n30576(n30576), 
         .n30575(n30575), .n30574(n30574), .n30573(n30573), .n30572(n30572), 
         .n30571(n30571), .n30570(n30570), .n30569(n30569), .n30568(n30568), 
         .n30567(n30567), .n30566(n30566), .n30565(n30565), .n30564(n30564), 
         .n30563(n30563), .n30562(n30562), .n30561(n30561), .n30560(n30560), 
         .n30559(n30559), .n30558(n30558), .n30557(n30557), .n30556(n30556), 
         .n30555(n30555), .n30554(n30554), .n30553(n30553), .n30552(n30552), 
         .n30551(n30551), .n30550(n30550), .n30549(n30549), .n30548(n30548), 
         .n30547(n30547), .n30546(n30546), .n30545(n30545), .n30544(n30544), 
         .n30543(n30543), .n30542(n30542), .n30541(n30541), .n30540(n30540), 
         .n30539(n30539), .n30538(n30538), .n30537(n30537), .n30536(n30536), 
         .n30535(n30535), .n30534(n30534), .n30533(n30533), .n30532(n30532), 
         .n30531(n30531), .n30530(n30530), .n30529(n30529), .n30528(n30528), 
         .n30527(n30527), .n30526(n30526), .n30525(n30525), .n30523(n30523), 
         .n30522(n30522), .n30521(n30521), .n30520(n30520), .n30519(n30519), 
         .n30518(n30518), .n30517(n30517), .n30516(n30516), .n30515(n30515), 
         .n30514(n30514), .n30513(n30513), .n30512(n30512), .n30511(n30511), 
         .n30510(n30510), .n30509(n30509), .n30508(n30508), .n30507(n30507), 
         .n30505(n30505), .n30504(n30504), .n30503(n30503), .n30502(n30502), 
         .n30500(n30500), .n30499(n30499), .n30498(n30498), .n30497(n30497), 
         .n30496(n30496), .n30495(n30495), .n30494(n30494), .n30493(n30493), 
         .n30492(n30492), .n30491(n30491), .n30490(n30490), .n30489(n30489), 
         .n30488(n30488), .n30487(n30487), .n30486(n30486), .n30485(n30485), 
         .n30484(n30484), .n30483(n30483), .n30482(n30482), .n30481(n30481), 
         .n30480(n30480), .n30479(n30479), .n30478(n30478), .n30477(n30477), 
         .n30476(n30476), .n30475(n30475), .n30474(n30474), .n30473(n30473), 
         .n30472(n30472), .n30471(n30471), .n30470(n30470), .n30469(n30469), 
         .n30468(n30468), .n30467(n30467), .n30466(n30466), .n30465(n30465), 
         .n30464(n30464), .n30463(n30463), .n30462(n30462), .n30461(n30461), 
         .n30460(n30460), .n30459(n30459), .n30458(n30458), .n30124(n30124), 
         .n30282(n30282), .n30281(n30281), .n30280(n30280), .n30279(n30279), 
         .n30278(n30278), .n30277(n30277), .n30276(n30276), .n30275(n30275), 
         .n30274(n30274), .n30273(n30273), .n30272(n30272), .n29618(n29618), 
         .n30271(n30271), .n30270(n30270), .n15(n15), .scl_enable_N_4177(scl_enable_N_4177), 
         .n6496(n6496), .n5_adj_4(n5_adj_5434), .n45649(n45649), .\displacement[4] (displacement[4]), 
         .n25701(n25701), .n47127(n47127), .n46329(n46329), .r_SM_Main({r_SM_Main_adj_5506}), 
         .n20694(n20694), .\r_Bit_Index[0] (r_Bit_Index_adj_5508[0]), .tx_o(tx_o), 
         .n29684(n29684), .n45512(n45512), .\r_SM_Main_2__N_3613[1] (r_SM_Main_2__N_3613[1]), 
         .n53023(n53023), .n30173(n30173), .n4(n4_adj_5349), .n30186(n30186), 
         .VCC_net(VCC_net), .tx_enable(tx_enable), .n29701(n29701), .n4_adj_5(n4_adj_5271), 
         .n4_adj_6(n4), .\r_Bit_Index[0]_adj_7 (r_Bit_Index[0]), .n28484(n28484), 
         .n35741(n35741), .r_SM_Main_adj_12({r_SM_Main}), .r_Rx_Data(r_Rx_Data), 
         .\r_SM_Main_2__N_3542[2] (r_SM_Main_2__N_3542[2]), .RX_N_10(RX_N_10), 
         .n28489(n28489), .n4_adj_11(n4_adj_5347), .n30197(n30197), .n45507(n45507), 
         .n30156(n30156), .n30155(n30155), .n30154(n30154), .n30153(n30153), 
         .n30152(n30152), .n30151(n30151), .n30150(n30150), .n45602(n45602), 
         .n29660(n29660), .n30189(n30189), .n45162(n45162)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(238[8] 261[4])
    SB_LUT4 i1_3_lut_adj_1837 (.I0(n2121), .I1(n2123), .I2(n2124), .I3(GND_net), 
            .O(n48601));
    defparam i1_3_lut_adj_1837.LUT_INIT = 16'hfefe;
    SB_LUT4 i16987_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n29618), 
            .I3(GND_net), .O(n30676));   // verilog/coms.v(127[12] 300[6])
    defparam i16987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5281));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16988_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n29618), 
            .I3(GND_net), .O(n30677));   // verilog/coms.v(127[12] 300[6])
    defparam i16988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16989_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n29618), 
            .I3(GND_net), .O(n30678));   // verilog/coms.v(127[12] 300[6])
    defparam i16989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16990_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n29618), 
            .I3(GND_net), .O(n30679));   // verilog/coms.v(127[12] 300[6])
    defparam i16990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16991_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n29618), 
            .I3(GND_net), .O(n30680));   // verilog/coms.v(127[12] 300[6])
    defparam i16991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16992_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n29618), 
            .I3(GND_net), .O(n30681));   // verilog/coms.v(127[12] 300[6])
    defparam i16992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i1_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16993_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n29618), 
            .I3(GND_net), .O(n30682));   // verilog/coms.v(127[12] 300[6])
    defparam i16993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i2_3_lut_4_lut (.I0(n28252), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16994_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n29618), 
            .I3(GND_net), .O(n30683));   // verilog/coms.v(127[12] 300[6])
    defparam i16994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16995_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n29618), 
            .I3(GND_net), .O(n30684));   // verilog/coms.v(127[12] 300[6])
    defparam i16995_3_lut.LUT_INIT = 16'hcaca;
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .pwm_setpoint({pwm_setpoint}), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (GND_net, timer, CLK_c, \neo_pixel_transmitter.t0 , 
            neopxl_color, VCC_net, n2956, n30251, n30250, n30249, 
            n30248, n30247, n30246, n30245, n30244, n30243, n30242, 
            n30241, n30240, n30239, n30238, n30237, n30236, n30235, 
            n30234, n30233, n30232, n30231, n30230, n30229, n30228, 
            n30227, n30226, n30225, n30224, n30223, n30222, n30221, 
            NEOPXL_c, LED_c, n30122) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]timer;
    input CLK_c;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input [23:0]neopxl_color;
    input VCC_net;
    output n2956;
    input n30251;
    input n30250;
    input n30249;
    input n30248;
    input n30247;
    input n30246;
    input n30245;
    input n30244;
    input n30243;
    input n30242;
    input n30241;
    input n30240;
    input n30239;
    input n30238;
    input n30237;
    input n30236;
    input n30235;
    input n30234;
    input n30233;
    input n30232;
    input n30231;
    input n30230;
    input n30229;
    input n30228;
    input n30227;
    input n30226;
    input n30225;
    input n30224;
    input n30223;
    input n30222;
    input n30221;
    output NEOPXL_c;
    input LED_c;
    input n30122;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [31:0]n133;
    
    wire n41756, n41757, \neo_pixel_transmitter.done_N_736 , n52965, 
        \neo_pixel_transmitter.done , start_N_727, n14, start, n75, 
        n125;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n51481, n46444, n51482, n38635, n46512, n46516, \neo_pixel_transmitter.done_N_742 ;
    wire [31:0]n255;
    
    wire n29590;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n30005, n41755, n41754, n41753, n41752;
    wire [31:0]n1;
    
    wire n41751, n50211, n50212, n50218, n50217, n2621, n52730, 
        n2495;
    wire [31:0]n2555;
    
    wire n2522, n2594, n2503, n2602, n2504, n2603, n2497, n2596, 
        n2494, n2593, n41750, n2491, n2590, n2499, n2598, n2507, 
        n2606, n2502, n2601, n2496, n2595, n2501, n2600, n2500, 
        n2599, n2508, n2607, n2492, n2591, n2509, n2608, n2498, 
        n2597, n2609, n2493, n2592, n2505, n2604, n2490, n2589, 
        n2506, n2605, n2588, n36, n25_adj_5154, n34, n40, n38, 
        n39, n37, n1103, n4, n40584, n1037;
    wire [31:0]n1070;
    
    wire n1005, n40583, n2406;
    wire [31:0]n2456;
    
    wire n2423, n2397, n2398, n2408, n2401, n2404, n2405, n2409, 
        n2400, n2407, n2403, n2402, n2396, n2391, n2395, n2393, 
        n2394, n2392, n2399, n26_adj_5155, n33_adj_5156, n2489, 
        n22_adj_5157, n38_adj_5158, n36_adj_5159, n37_adj_5160, n35, 
        n41749, n1006, n40582, n41748, n132, n45645, n1007, n40581, 
        n41747, n41746, n2308;
    wire [31:0]n2357;
    
    wire n2324, n2307, n2306, n41745, n41744, n2304, n2305, n2303, 
        n2298, n2296, n2297, n2295, n2294, n2293, n2292, n1008, 
        n40580, n2301, n41743, n2300, n1009, n40579, n2302, n2299, 
        n41742, n2309, n27_adj_5161, n33_adj_5162, n32_adj_5163, n2390, 
        n31_adj_5164, n35_adj_5165, n37_adj_5166, n41741, n43736, 
        n52230, n2205;
    wire [31:0]n2258;
    
    wire n2225, n2208, n41740, n2197, n2201, n2207, n2206, n2209, 
        n2203, n2202, n2200, n2199, n2193, n2204, n2198, n2195, 
        n2196, n2194, n30_adj_5168, n41739, n36610, n2291, n34_adj_5169, 
        n32_adj_5170, n33_adj_5171, n31_adj_5172, n2100;
    wire [31:0]n2159;
    
    wire n2126, n2098, n2099, n2097, n2108, n2103, n2105, n2109, 
        n2106, n2102, n2101, n2107, n2104, n2096, n2095, n2094, 
        n2192, n28_adj_5173, n36608, n32_adj_5174, n30_adj_5175, n31_adj_5176, 
        n29_adj_5177, n2004;
    wire [31:0]n2060;
    
    wire n2027, n1997, n1996, n1998, n2002, n1999, n2005, n2008, 
        n2006, n2000, n2001, n2009, n2003, n2007, n1995, n2093, 
        n18_adj_5178, n36606, n30_adj_5179, n28_adj_5180, n29_adj_5181, 
        n27_adj_5182, n1898;
    wire [31:0]n1961;
    
    wire n1928, n1897, n1896, n1902, n1900, n1901, n1899, n1908, 
        n1903, n1909, n1907, n1906, n1905, n1904, n36604, n28_adj_5183, 
        n26_adj_5184, n27_adj_5185, n1994, n25_adj_5186, n36602, n26_adj_5187, 
        n24_adj_5188, n25_adj_5189, n1895, n23_adj_5190, n51038, n38580, 
        n12_adj_5191, n1829, n52729, n40466, n40465, n40464, n1202, 
        n41731, n1136;
    wire [31:0]n1169;
    
    wire n1104, n41730, n1105, n41729, n1106, n41728, n1107, n41727, 
        n1108, n41726, n40463, n40462, n1109, n41725, n1400, n1301, 
        n41724, n1334;
    wire [31:0]n1367;
    
    wire n1302, n41723, n1303, n41722, n1304, n41721;
    wire [3:0]state_3__N_528;
    
    wire n7_adj_5192, n38562, n1305, n41720, n40461, n1306, n41719, 
        n1307, n41718, n40460, n1308, n41717, n1309, n41716;
    wire [31:0]n971;
    
    wire n28470, n40630, n49915, n40629, n49913, n40628, n49911, 
        n42258, n1235;
    wire [31:0]n1268;
    
    wire n1203, n42257, n1204, n42256, n1205, n42255, n1206, n42254, 
        n1207, n42253, n1208, n42252, n1209, n42251, n1697, n1598, 
        n42250, n1631;
    wire [31:0]n1664;
    
    wire n1599, n42249, n1600, n42248, n1601, n42247, n1602, n42246, 
        n1603, n42245, n1604, n42244, n1605, n42243, n1606, n42242, 
        n1607, n42241, n1608, n42240, n1609, n42239, n1796, n42238, 
        n1730;
    wire [31:0]n1763;
    
    wire n1698, n42237, n1707, n1806, n1700, n1799, n1709, n1808, 
        n1708, n1807, n1699, n1798, n1797, n1704, n1803, n1702, 
        n1801, n42236, n42235, n1809, n1701, n42234, n42233, n1703, 
        n42232, n42231, n1705, n42230, n1706, n42229, n42228, 
        n1800, n42227, n42226, n42225, n42224, n42223, n1804, 
        n42222, n42221, n42220, n1802, n42219, n42218, n42217, 
        n1805, n24_adj_5194, n17_adj_5195, n42216, n40627, n49909, 
        n22_adj_5196, n40626, n49907, n26_adj_5197, n42215, n42214, 
        n42213, n42212, n42211, n42210, n42209, n42208, n42207, 
        n42206, n42205, n52930, n50183, n42204, n42203, n42202, 
        n42201, n42200, n42199, n42198, n42197, n42196, n52888, 
        n42195, n50261, n42194, n42193, n42192, n42191, n42190, 
        n42189, n42188, n42187, n42186, n42185, n42184, n42183, 
        n42182, n42181, n40625, n49905, n40459, n42180, n42179, 
        n42178, n42177, n42176, n42175, n42174, n42173, n42172, 
        n42171, n42170, n42169, n42168, n42167, n42166, n42165, 
        n42164, n42163, n42162, n42161, n42160, n42159, n42158, 
        n40624, n49903, n807, n838, n12165, n46352, n50068, n906, 
        n42157, n42156, n42155, n42154, n42153, n26840, n739, 
        n26854, n36796, n708, n46742, n13435, n608, n52882, n42152, 
        n42151, n40623, n49901, n42150, n29881, n42149, n42148, 
        n42147, n46442, n49527, n42146, n40458, n46437, n7_adj_5198, 
        n40622, n49899, n42145, n42144, n40457, n40704, n42143, 
        n50267, n42142, n42141, n42140, n40456, n42139, n42138, 
        n42137, n40621, n49897, n42136, n42135, n42134, n42133, 
        n42132, n40455, n40703, n40702, n40701, n42131, n40620, 
        n49895, n40700, n42130, n42129, n42128, n42127, n40619, 
        n49893, n40618, n49891, n42126, n42125, n42124, n40454, 
        n42123, n42122, n42121, n42120, n42119, n42118, n40617, 
        n49889, n42117, n40453, n42116, n40616, n49887, n42115, 
        n42114, n40452, n42113, n42112, n42111, n42110, n42109, 
        n40615, n49885, n42108, n42107, n42106, n42105, n42104, 
        n40614, n49883, n40613, n49881, n42103, n42102, n42101, 
        n42100, n42099, n42098, n42097, n40612, n49879, n42096, 
        n42095, n42094, n42093, n42092, n42091, n42090, n40451, 
        n42089, n42088, n18_adj_5199, n21_adj_5200, n20_adj_5201, 
        n42087, n24_adj_5202, n40611;
    wire [31:0]one_wire_N_679;
    
    wire n42086, n40610, n2687, n42085, n2688, n42084, n2689, 
        n42083, n2690, n42082, n2691, n42081, n2692, n42080, n2693, 
        n42079, n40450, n1505;
    wire [31:0]n1565;
    
    wire n1532, n1509, n1508, n1503, n2694, n42078, n40449, n2695, 
        n42077, n2696, n42076, n2697, n42075, n2698, n42074, n2699, 
        n42073, n2700, n42072, n40609, n2701, n42071, n2702, n42070, 
        n38636, n2703, n42069, n2704, n42068, n2705, n42067, n2706, 
        n42066, n2707, n42065, n2708, n42064, n2709, n40448, n2786, 
        n42063, n2720;
    wire [31:0]n2753;
    
    wire n42062, n1502, n1501, n1500, n40608, n42061, n42060, 
        n42059, n1506, n42058, n1507, n42057, n42056, n42055, 
        n42054, n1407;
    wire [31:0]n1466;
    
    wire n1433, n40447, n1499, n41084, n42053, n42052, n42051, 
        n1401, n41083, n42050, n42049, n42048, n42047, n1402, 
        n41082, n42046, n40607, n1403, n41081, n52810, n52813, 
        n42045, n1404, n41080, n42044, n42043, n42042, n42041, 
        n40446, n2885, n42040, n2819, n1405, n41079;
    wire [31:0]n2852;
    
    wire n2787, n42039, n2788, n42038, n2789, n42037, n1406, n41078, 
        n49873, n40606, n49871, n40445, n2790, n42036, n2791, 
        n42035, n1408, n2792, n42034, n2793, n42033, n2794, n42032, 
        n2795, n42031, n2796, n42030, n2797, n42029, n2798, n42028, 
        n41077, n41076, n2799, n42027, n1409, n41075, n40605, 
        n49869, n2800, n42026, n2801, n42025, n2802, n42024, n1504, 
        n2803, n42023, n40604, n2804, n42022, n16_adj_5203, n18_adj_5204, 
        n13_adj_5205, n2805, n42021, n2806, n42020, n40444, n2807, 
        n42019, n2808, n42018, n2809, n42017, n2984, n42016, n2918;
    wire [31:0]n2951;
    
    wire n2886, n42015, n36636, n18_adj_5206, n2887, n42014, n16_adj_5207, 
        n20_adj_5208, n2888, n42013, n16_adj_5209, n40603, n19_adj_5210, 
        n18_adj_5211, n2889, n42012, n22_adj_5213, n2890, n42011, 
        n38574, n98, n46, n44, n45, n43, n42, n41, n52, n47, 
        n43659, n42573, n42886, n2891, n42010, n40602, n2892, 
        n42009, n2893, n42008, n2894, n42007, n51058, n18_adj_5214, 
        n2895, n42006, n51053, n40601, n4_adj_5215, n40600, n2896, 
        n42005, n2897, n42004, n40443, n2898, n42003, n2899, n42002, 
        n2900, n42001, n2901, n42000, n2902, n41999, n2903, n41998, 
        n40442, n41044, n2904, n41997, n2905, n41996, n2906, n41995, 
        n2907, n41994, n41043, n41042, n41041, n41040, n41039, 
        n41038, n2908, n41993, n41037, n41036, n41035, n41034, 
        n48388, n55, n121, n46488, n8_adj_5216, n7_adj_5217, n40441, 
        n2909, n41992, n40440, n3083, n41991, n3017;
    wire [31:0]n3050;
    
    wire n2985, n41990, n2986, n41989, n2987, n41988, n2988, n41987, 
        n2989, n41986, n2990, n41985, n2991, n41984, n2992, n41983, 
        n2993, n41982, n2994, n41981, n2995, n41980, n2996, n41979, 
        n2997, n41978, n2998, n41977, n2999, n41976, n3000, n41975, 
        n3001, n41974, n3002, n41973, n3003, n41972, n3004, n41971, 
        n3005, n41970, n3006, n41969, n3007, n41968, n3008, n41967, 
        n3009, n41966, n50010, n41965, n3116;
    wire [31:0]n3149;
    
    wire n3084, n41964, n3085, n41963, n3086, n41962, n3087, n41961, 
        n3088, n41960, n3089, n41959, n3090, n41958, n3091, n41957, 
        n3092, n41956, n3093, n41955, n3094, n41954, n3095, n41953, 
        n3096, n41952, n3097, n41951, n3098, n41950, n3099, n41949, 
        n3100, n41948, n3101, n41947, n3102, n41946, n3103, n41945, 
        n3104, n41944, n3105, n41943, n3106, n41942, n3107, n41941, 
        n3108, n41940, n3109, n41939, n52768, n40439, n40438, 
        n52735, n52771, n40437, n40436, n41769, n41768, n41767, 
        n41766, n41765, n41764, n41763, n41762, n41761, n41760, 
        n41759, n41758, n128, n28_adj_5218, n38_adj_5219, n36_adj_5220, 
        n42_adj_5221, n40_adj_5222, n41_adj_5223, n39_adj_5224, n32_adj_5225, 
        n39_adj_5226, n26_adj_5227, n38_adj_5228, n44_adj_5229, n42_adj_5230, 
        n43_adj_5231, n41_adj_5232, n30_adj_5233, n39_adj_5234, n38_adj_5235, 
        n43_adj_5236, n42_adj_5237, n41_adj_5238, n45_adj_5239, n47_adj_5240, 
        n34_adj_5241, n44_adj_5242, n40_adj_5243, n45_adj_5244, n42_adj_5245, 
        n48, n41_adj_5246, n49, n36_adj_5247, n46_adj_5248, n42_adj_5249, 
        n33_adj_5250, n43_adj_5251, n50, n48_adj_5252, n49_adj_5253, 
        n47_adj_5254, n21_adj_5255, n25_adj_5256, n11_adj_5257, n49309, 
        n15_adj_5258, n29_adj_5259, n49313, n49315, n49317, n49311, 
        n49319, n33_adj_5260, n3209, n49327, n49329, n35_adj_5261, 
        n37_adj_5262, n49335, n49337, n49339, n49341, n49343, n49345, 
        n49347, n49349, n49351, n49353, n49355, n59, n61, n51034, 
        n10_adj_5263;
    wire [4:0]color_bit_N_722;
    
    wire n51115, n11_adj_5264, n13_adj_5265, n10_adj_5266, n16_adj_5267, 
        n11_adj_5268, n10_adj_5269, n12_adj_5270, n52732;
    
    SB_LUT4 timer_2188_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n41756), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_20 (.CI(n41756), .I0(GND_net), .I1(timer[18]), 
            .CO(n41757));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n52965), .D(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(n14), .D(start_N_727));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i36048_4_lut (.I0(n75), .I1(n125), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n51481));
    defparam i36048_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i35847_3_lut (.I0(state[1]), .I1(n51481), .I2(n46444), .I3(GND_net), 
            .O(n51482));
    defparam i35847_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i53_4_lut (.I0(n46444), .I1(n38635), .I2(state[1]), .I3(n125), 
            .O(n46512));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i56_4_lut (.I0(n46512), .I1(n51482), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n46516));
    defparam i56_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_742 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n29590), .D(n255[1]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n29590), .D(n255[2]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n29590), .D(n255[3]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n29590), .D(n255[4]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n29590), .D(n255[5]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n29590), .D(n255[6]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n29590), .D(n255[7]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n29590), .D(n255[8]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n29590), .D(n255[9]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n29590), 
            .D(n255[10]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n29590), 
            .D(n255[11]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n29590), 
            .D(n255[12]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n29590), 
            .D(n255[13]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n29590), 
            .D(n255[14]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n29590), 
            .D(n255[15]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n29590), 
            .D(n255[16]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n29590), 
            .D(n255[17]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n29590), 
            .D(n255[18]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n29590), 
            .D(n255[19]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n29590), 
            .D(n255[20]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n29590), 
            .D(n255[21]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n29590), 
            .D(n255[22]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n29590), 
            .D(n255[23]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n29590), 
            .D(n255[24]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n29590), 
            .D(n255[25]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n29590), 
            .D(n255[26]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n29590), 
            .D(n255[27]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n29590), 
            .D(n255[28]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n29590), 
            .D(n255[29]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n29590), 
            .D(n255[30]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n29590), 
            .D(n255[31]), .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2188_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n41755), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_19 (.CI(n41755), .I0(GND_net), .I1(timer[17]), 
            .CO(n41756));
    SB_LUT4 timer_2188_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n41754), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_18 (.CI(n41754), .I0(GND_net), .I1(timer[16]), 
            .CO(n41755));
    SB_LUT4 timer_2188_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n41753), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_17 (.CI(n41753), .I0(GND_net), .I1(timer[15]), 
            .CO(n41754));
    SB_LUT4 timer_2188_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n41752), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_16 (.CI(n41752), .I0(GND_net), .I1(timer[14]), 
            .CO(n41753));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2188_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n41751), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34577_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50211));
    defparam i34577_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_15 (.CI(n41751), .I0(GND_net), .I1(timer[13]), 
            .CO(n41752));
    SB_LUT4 i34578_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50212));
    defparam i34578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34584_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50218));
    defparam i34584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34583_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n50217));
    defparam i34583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i37095_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52730));
    defparam i37095_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1749_3_lut (.I0(n2495), .I1(n2555[25]), .I2(n2522), 
            .I3(GND_net), .O(n2594));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1757_3_lut (.I0(n2503), .I1(n2555[17]), .I2(n2522), 
            .I3(GND_net), .O(n2602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1758_3_lut (.I0(n2504), .I1(n2555[16]), .I2(n2522), 
            .I3(GND_net), .O(n2603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1751_3_lut (.I0(n2497), .I1(n2555[23]), .I2(n2522), 
            .I3(GND_net), .O(n2596));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1748_3_lut (.I0(n2494), .I1(n2555[26]), .I2(n2522), 
            .I3(GND_net), .O(n2593));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n41750), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1745_3_lut (.I0(n2491), .I1(n2555[29]), .I2(n2522), 
            .I3(GND_net), .O(n2590));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1753_3_lut (.I0(n2499), .I1(n2555[21]), .I2(n2522), 
            .I3(GND_net), .O(n2598));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1761_3_lut (.I0(n2507), .I1(n2555[13]), .I2(n2522), 
            .I3(GND_net), .O(n2606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1756_3_lut (.I0(n2502), .I1(n2555[18]), .I2(n2522), 
            .I3(GND_net), .O(n2601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1750_3_lut (.I0(n2496), .I1(n2555[24]), .I2(n2522), 
            .I3(GND_net), .O(n2595));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1755_3_lut (.I0(n2501), .I1(n2555[19]), .I2(n2522), 
            .I3(GND_net), .O(n2600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1754_3_lut (.I0(n2500), .I1(n2555[20]), .I2(n2522), 
            .I3(GND_net), .O(n2599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1762_3_lut (.I0(n2508), .I1(n2555[12]), .I2(n2522), 
            .I3(GND_net), .O(n2607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1746_3_lut (.I0(n2492), .I1(n2555[28]), .I2(n2522), 
            .I3(GND_net), .O(n2591));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1763_3_lut (.I0(n2509), .I1(n2555[11]), .I2(n2522), 
            .I3(GND_net), .O(n2608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1752_3_lut (.I0(n2498), .I1(n2555[22]), .I2(n2522), 
            .I3(GND_net), .O(n2597));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1764_3_lut (.I0(bit_ctr[10]), .I1(n2555[10]), .I2(n2522), 
            .I3(GND_net), .O(n2609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1747_3_lut (.I0(n2493), .I1(n2555[27]), .I2(n2522), 
            .I3(GND_net), .O(n2592));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1759_3_lut (.I0(n2505), .I1(n2555[15]), .I2(n2522), 
            .I3(GND_net), .O(n2604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1744_3_lut (.I0(n2490), .I1(n2555[30]), .I2(n2522), 
            .I3(GND_net), .O(n2589));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1760_3_lut (.I0(n2506), .I1(n2555[14]), .I2(n2522), 
            .I3(GND_net), .O(n2605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(n2605), .I1(n2588), .I2(n2589), .I3(n2604), 
            .O(n36));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2592), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_5154));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut (.I0(n2597), .I1(n2608), .I2(n2591), .I3(n2607), 
            .O(n34));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n25_adj_5154), .I1(n36), .I2(n2599), .I3(n2600), 
            .O(n40));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2595), .I1(n2601), .I2(n2606), .I3(n2598), 
            .O(n38));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2602), .I1(n34), .I2(n2594), .I3(GND_net), 
            .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut (.I0(n2590), .I1(n2593), .I2(n2596), .I3(n2603), 
            .O(n37));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n2621));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n1037), .I1(n4), .I2(VCC_net), .I3(n40584), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_736_7_lut (.I0(GND_net), .I1(n1005), .I2(VCC_net), 
            .I3(n40583), .O(n1070[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_7 (.CI(n40583), .I0(n1005), .I1(VCC_net), .CO(n40584));
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1692_3_lut (.I0(n2406), .I1(n2456[15]), .I2(n2423), 
            .I3(GND_net), .O(n2505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1683_3_lut (.I0(n2397), .I1(n2456[24]), .I2(n2423), 
            .I3(GND_net), .O(n2496));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1684_3_lut (.I0(n2398), .I1(n2456[23]), .I2(n2423), 
            .I3(GND_net), .O(n2497));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1694_3_lut (.I0(n2408), .I1(n2456[13]), .I2(n2423), 
            .I3(GND_net), .O(n2507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1687_3_lut (.I0(n2401), .I1(n2456[20]), .I2(n2423), 
            .I3(GND_net), .O(n2500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1690_3_lut (.I0(n2404), .I1(n2456[17]), .I2(n2423), 
            .I3(GND_net), .O(n2503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1691_3_lut (.I0(n2405), .I1(n2456[16]), .I2(n2423), 
            .I3(GND_net), .O(n2504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1695_3_lut (.I0(n2409), .I1(n2456[12]), .I2(n2423), 
            .I3(GND_net), .O(n2508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1686_3_lut (.I0(n2400), .I1(n2456[21]), .I2(n2423), 
            .I3(GND_net), .O(n2499));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1693_3_lut (.I0(n2407), .I1(n2456[14]), .I2(n2423), 
            .I3(GND_net), .O(n2506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1689_3_lut (.I0(n2403), .I1(n2456[18]), .I2(n2423), 
            .I3(GND_net), .O(n2502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1688_3_lut (.I0(n2402), .I1(n2456[19]), .I2(n2423), 
            .I3(GND_net), .O(n2501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1682_3_lut (.I0(n2396), .I1(n2456[25]), .I2(n2423), 
            .I3(GND_net), .O(n2495));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1677_3_lut (.I0(n2391), .I1(n2456[30]), .I2(n2423), 
            .I3(GND_net), .O(n2490));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1681_3_lut (.I0(n2395), .I1(n2456[26]), .I2(n2423), 
            .I3(GND_net), .O(n2494));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1679_3_lut (.I0(n2393), .I1(n2456[28]), .I2(n2423), 
            .I3(GND_net), .O(n2492));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1680_3_lut (.I0(n2394), .I1(n2456[27]), .I2(n2423), 
            .I3(GND_net), .O(n2493));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1678_3_lut (.I0(n2392), .I1(n2456[29]), .I2(n2423), 
            .I3(GND_net), .O(n2491));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1696_3_lut (.I0(bit_ctr[11]), .I1(n2456[11]), .I2(n2423), 
            .I3(GND_net), .O(n2509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1685_3_lut (.I0(n2399), .I1(n2456[22]), .I2(n2423), 
            .I3(GND_net), .O(n2498));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(n2498), .I1(bit_ctr[10]), .I2(n2509), .I3(GND_net), 
            .O(n26_adj_5155));
    defparam i5_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1529 (.I0(n2491), .I1(n2493), .I2(n2492), .I3(n2494), 
            .O(n33_adj_5156));
    defparam i12_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(n2490), .I1(n2489), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_5157));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut (.I0(n33_adj_5156), .I1(n2495), .I2(n26_adj_5155), 
            .I3(n2501), .O(n38_adj_5158));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1530 (.I0(n2502), .I1(n2506), .I2(n2499), .I3(n2508), 
            .O(n36_adj_5159));
    defparam i15_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1531 (.I0(n2504), .I1(n2503), .I2(n2500), .I3(n22_adj_5157), 
            .O(n37_adj_5160));
    defparam i16_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1532 (.I0(n2507), .I1(n2497), .I2(n2496), .I3(n2505), 
            .O(n35));
    defparam i14_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37_adj_5160), .I2(n36_adj_5159), 
            .I3(n38_adj_5158), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2188_add_4_14 (.CI(n41750), .I0(GND_net), .I1(timer[12]), 
            .CO(n41751));
    SB_LUT4 timer_2188_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n41749), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_6_lut (.I0(GND_net), .I1(n1006), .I2(VCC_net), 
            .I3(n40582), .O(n1070[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_13 (.CI(n41749), .I0(GND_net), .I1(timer[11]), 
            .CO(n41750));
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2188_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n41748), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24917_4_lut (.I0(n125), .I1(n75), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n132));   // verilog/neopixel.v(16[20:25])
    defparam i24917_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(n132), .I2(n45645), .I3(start), 
            .O(n2956));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2188_add_4_12 (.CI(n41748), .I0(GND_net), .I1(timer[10]), 
            .CO(n41749));
    SB_CARRY mod_5_add_736_6 (.CI(n40582), .I0(n1006), .I1(VCC_net), .CO(n40583));
    SB_LUT4 mod_5_add_736_5_lut (.I0(GND_net), .I1(n1007), .I2(VCC_net), 
            .I3(n40581), .O(n1070[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2188_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n41747), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_11 (.CI(n41747), .I0(GND_net), .I1(timer[9]), 
            .CO(n41748));
    SB_LUT4 timer_2188_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n41746), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_10 (.CI(n41746), .I0(GND_net), .I1(timer[8]), 
            .CO(n41747));
    SB_LUT4 mod_5_i1626_3_lut (.I0(n2308), .I1(n2357[14]), .I2(n2324), 
            .I3(GND_net), .O(n2407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1625_3_lut (.I0(n2307), .I1(n2357[15]), .I2(n2324), 
            .I3(GND_net), .O(n2406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1624_3_lut (.I0(n2306), .I1(n2357[16]), .I2(n2324), 
            .I3(GND_net), .O(n2405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n41745), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_9 (.CI(n41745), .I0(GND_net), .I1(timer[7]), 
            .CO(n41746));
    SB_CARRY mod_5_add_736_5 (.CI(n40581), .I0(n1007), .I1(VCC_net), .CO(n40582));
    SB_LUT4 timer_2188_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n41744), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1622_3_lut (.I0(n2304), .I1(n2357[18]), .I2(n2324), 
            .I3(GND_net), .O(n2403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1622_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_8 (.CI(n41744), .I0(GND_net), .I1(timer[6]), 
            .CO(n41745));
    SB_LUT4 mod_5_i1623_3_lut (.I0(n2305), .I1(n2357[17]), .I2(n2324), 
            .I3(GND_net), .O(n2404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1621_3_lut (.I0(n2303), .I1(n2357[19]), .I2(n2324), 
            .I3(GND_net), .O(n2402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1616_3_lut (.I0(n2298), .I1(n2357[24]), .I2(n2324), 
            .I3(GND_net), .O(n2397));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1614_3_lut (.I0(n2296), .I1(n2357[26]), .I2(n2324), 
            .I3(GND_net), .O(n2395));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1615_3_lut (.I0(n2297), .I1(n2357[25]), .I2(n2324), 
            .I3(GND_net), .O(n2396));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1613_3_lut (.I0(n2295), .I1(n2357[27]), .I2(n2324), 
            .I3(GND_net), .O(n2394));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1612_3_lut (.I0(n2294), .I1(n2357[28]), .I2(n2324), 
            .I3(GND_net), .O(n2393));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1611_3_lut (.I0(n2293), .I1(n2357[29]), .I2(n2324), 
            .I3(GND_net), .O(n2392));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1610_3_lut (.I0(n2292), .I1(n2357[30]), .I2(n2324), 
            .I3(GND_net), .O(n2391));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_736_4_lut (.I0(GND_net), .I1(n1008), .I2(VCC_net), 
            .I3(n40580), .O(n1070[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_4 (.CI(n40580), .I0(n1008), .I1(VCC_net), .CO(n40581));
    SB_LUT4 mod_5_i1619_3_lut (.I0(n2301), .I1(n2357[21]), .I2(n2324), 
            .I3(GND_net), .O(n2400));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n41743), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1618_3_lut (.I0(n2300), .I1(n2357[22]), .I2(n2324), 
            .I3(GND_net), .O(n2399));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_736_3_lut (.I0(GND_net), .I1(n1009), .I2(GND_net), 
            .I3(n40579), .O(n1070[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1620_3_lut (.I0(n2302), .I1(n2357[20]), .I2(n2324), 
            .I3(GND_net), .O(n2401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1620_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_7 (.CI(n41743), .I0(GND_net), .I1(timer[5]), 
            .CO(n41744));
    SB_LUT4 mod_5_i1617_3_lut (.I0(n2299), .I1(n2357[23]), .I2(n2324), 
            .I3(GND_net), .O(n2398));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n41742), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1628_3_lut (.I0(bit_ctr[12]), .I1(n2357[12]), .I2(n2324), 
            .I3(GND_net), .O(n2409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1627_3_lut (.I0(n2309), .I1(n2357[13]), .I2(n2324), 
            .I3(GND_net), .O(n2408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2408), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_5161));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut (.I0(n2398), .I1(n2401), .I2(n2399), .I3(n2400), 
            .O(n33_adj_5162));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1533 (.I0(n2394), .I1(n2396), .I2(n2395), .I3(n2397), 
            .O(n32_adj_5163));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2391), .I1(n2392), .I2(n2390), .I3(n2393), 
            .O(n31_adj_5164));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1534 (.I0(n2402), .I1(n2404), .I2(n2403), .I3(n2405), 
            .O(n35_adj_5165));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1535 (.I0(n33_adj_5162), .I1(n27_adj_5161), .I2(n2406), 
            .I3(n2407), .O(n37_adj_5166));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37_adj_5166), .I1(n35_adj_5165), .I2(n31_adj_5164), 
            .I3(n32_adj_5163), .O(n2423));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2188_add_4_6 (.CI(n41742), .I0(GND_net), .I1(timer[4]), 
            .CO(n41743));
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_736_3 (.CI(n40579), .I0(n1009), .I1(GND_net), .CO(n40580));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2188_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n41741), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36595_1_lut (.I0(n43736), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52230));   // verilog/neopixel.v(22[26:36])
    defparam i36595_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2188_add_4_5 (.CI(n41741), .I0(GND_net), .I1(timer[3]), 
            .CO(n41742));
    SB_LUT4 mod_5_i1555_3_lut (.I0(n2205), .I1(n2258[18]), .I2(n2225), 
            .I3(GND_net), .O(n2304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1558_3_lut (.I0(n2208), .I1(n2258[15]), .I2(n2225), 
            .I3(GND_net), .O(n2307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n41740), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1547_3_lut (.I0(n2197), .I1(n2258[26]), .I2(n2225), 
            .I3(GND_net), .O(n2296));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1551_3_lut (.I0(n2201), .I1(n2258[22]), .I2(n2225), 
            .I3(GND_net), .O(n2300));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1557_3_lut (.I0(n2207), .I1(n2258[16]), .I2(n2225), 
            .I3(GND_net), .O(n2306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1556_3_lut (.I0(n2206), .I1(n2258[17]), .I2(n2225), 
            .I3(GND_net), .O(n2305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1559_3_lut (.I0(n2209), .I1(n2258[14]), .I2(n2225), 
            .I3(GND_net), .O(n2308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1553_3_lut (.I0(n2203), .I1(n2258[20]), .I2(n2225), 
            .I3(GND_net), .O(n2302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1552_3_lut (.I0(n2202), .I1(n2258[21]), .I2(n2225), 
            .I3(GND_net), .O(n2301));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1550_3_lut (.I0(n2200), .I1(n2258[23]), .I2(n2225), 
            .I3(GND_net), .O(n2299));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1549_3_lut (.I0(n2199), .I1(n2258[24]), .I2(n2225), 
            .I3(GND_net), .O(n2298));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1543_3_lut (.I0(n2193), .I1(n2258[30]), .I2(n2225), 
            .I3(GND_net), .O(n2292));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1554_3_lut (.I0(n2204), .I1(n2258[19]), .I2(n2225), 
            .I3(GND_net), .O(n2303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1554_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_4 (.CI(n41740), .I0(GND_net), .I1(timer[2]), 
            .CO(n41741));
    SB_LUT4 mod_5_i1560_3_lut (.I0(bit_ctr[13]), .I1(n2258[13]), .I2(n2225), 
            .I3(GND_net), .O(n2309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1548_3_lut (.I0(n2198), .I1(n2258[25]), .I2(n2225), 
            .I3(GND_net), .O(n2297));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_736_2_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(VCC_net), .O(n1070[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1545_3_lut (.I0(n2195), .I1(n2258[28]), .I2(n2225), 
            .I3(GND_net), .O(n2294));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1546_3_lut (.I0(n2196), .I1(n2258[27]), .I2(n2225), 
            .I3(GND_net), .O(n2295));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1544_3_lut (.I0(n2194), .I1(n2258[29]), .I2(n2225), 
            .I3(GND_net), .O(n2293));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1536 (.I0(n2293), .I1(n2295), .I2(n2294), .I3(n2297), 
            .O(n30_adj_5168));
    defparam i11_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2188_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n41739), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22928_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n36610));
    defparam i22928_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut_adj_1537 (.I0(n2303), .I1(n30_adj_5168), .I2(n2292), 
            .I3(n2291), .O(n34_adj_5169));
    defparam i15_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(GND_net), 
            .CO(n40579));
    SB_LUT4 i13_4_lut_adj_1538 (.I0(n2308), .I1(n2305), .I2(n2306), .I3(n2300), 
            .O(n32_adj_5170));
    defparam i13_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1539 (.I0(n2298), .I1(n2299), .I2(n2301), .I3(n2302), 
            .O(n33_adj_5171));
    defparam i14_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1540 (.I0(n2296), .I1(n36610), .I2(n2307), .I3(n2304), 
            .O(n31_adj_5172));
    defparam i12_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n30251));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n30250));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n30249));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n30248));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i18_4_lut_adj_1541 (.I0(n31_adj_5172), .I1(n33_adj_5171), .I2(n32_adj_5170), 
            .I3(n34_adj_5169), .O(n2324));
    defparam i18_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n30247));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n30246));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n30245));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n30244));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n30243));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n30242));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_2188_add_4_3 (.CI(n41739), .I0(GND_net), .I1(timer[1]), 
            .CO(n41740));
    SB_LUT4 timer_2188_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n30241));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1482_3_lut (.I0(n2100), .I1(n2159[24]), .I2(n2126), 
            .I3(GND_net), .O(n2199));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1480_3_lut (.I0(n2098), .I1(n2159[26]), .I2(n2126), 
            .I3(GND_net), .O(n2197));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1481_3_lut (.I0(n2099), .I1(n2159[25]), .I2(n2126), 
            .I3(GND_net), .O(n2198));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1479_3_lut (.I0(n2097), .I1(n2159[27]), .I2(n2126), 
            .I3(GND_net), .O(n2196));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1490_3_lut (.I0(n2108), .I1(n2159[16]), .I2(n2126), 
            .I3(GND_net), .O(n2207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1485_3_lut (.I0(n2103), .I1(n2159[21]), .I2(n2126), 
            .I3(GND_net), .O(n2202));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1487_3_lut (.I0(n2105), .I1(n2159[19]), .I2(n2126), 
            .I3(GND_net), .O(n2204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1491_3_lut (.I0(n2109), .I1(n2159[15]), .I2(n2126), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1488_3_lut (.I0(n2106), .I1(n2159[18]), .I2(n2126), 
            .I3(GND_net), .O(n2205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1484_3_lut (.I0(n2102), .I1(n2159[22]), .I2(n2126), 
            .I3(GND_net), .O(n2201));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1483_3_lut (.I0(n2101), .I1(n2159[23]), .I2(n2126), 
            .I3(GND_net), .O(n2200));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1489_3_lut (.I0(n2107), .I1(n2159[17]), .I2(n2126), 
            .I3(GND_net), .O(n2206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1486_3_lut (.I0(n2104), .I1(n2159[20]), .I2(n2126), 
            .I3(GND_net), .O(n2203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1492_3_lut (.I0(bit_ctr[14]), .I1(n2159[14]), .I2(n2126), 
            .I3(GND_net), .O(n2209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1478_3_lut (.I0(n2096), .I1(n2159[28]), .I2(n2126), 
            .I3(GND_net), .O(n2195));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1477_3_lut (.I0(n2095), .I1(n2159[29]), .I2(n2126), 
            .I3(GND_net), .O(n2194));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1476_3_lut (.I0(n2094), .I1(n2159[30]), .I2(n2126), 
            .I3(GND_net), .O(n2193));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(n2193), .I1(n2194), .I2(n2192), .I3(n2195), 
            .O(n28_adj_5173));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22926_2_lut (.I0(bit_ctr[13]), .I1(n2209), .I2(GND_net), 
            .I3(GND_net), .O(n36608));
    defparam i22926_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_3_lut (.I0(n2203), .I1(n28_adj_5173), .I2(n2206), .I3(GND_net), 
            .O(n32_adj_5174));
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1542 (.I0(n2200), .I1(n2201), .I2(n2205), .I3(n36608), 
            .O(n30_adj_5175));
    defparam i12_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1543 (.I0(n2208), .I1(n2204), .I2(n2202), .I3(n2207), 
            .O(n31_adj_5176));
    defparam i13_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1544 (.I0(n2196), .I1(n2198), .I2(n2197), .I3(n2199), 
            .O(n29_adj_5177));
    defparam i11_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1545 (.I0(n29_adj_5177), .I1(n31_adj_5176), .I2(n30_adj_5175), 
            .I3(n32_adj_5174), .O(n2225));
    defparam i17_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1418_3_lut (.I0(n2004), .I1(n2060[21]), .I2(n2027), 
            .I3(GND_net), .O(n2103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1411_3_lut (.I0(n1997), .I1(n2060[28]), .I2(n2027), 
            .I3(GND_net), .O(n2096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1410_3_lut (.I0(n1996), .I1(n2060[29]), .I2(n2027), 
            .I3(GND_net), .O(n2095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1412_3_lut (.I0(n1998), .I1(n2060[27]), .I2(n2027), 
            .I3(GND_net), .O(n2097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1416_3_lut (.I0(n2002), .I1(n2060[23]), .I2(n2027), 
            .I3(GND_net), .O(n2101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1413_3_lut (.I0(n1999), .I1(n2060[26]), .I2(n2027), 
            .I3(GND_net), .O(n2098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1419_3_lut (.I0(n2005), .I1(n2060[20]), .I2(n2027), 
            .I3(GND_net), .O(n2104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1422_3_lut (.I0(n2008), .I1(n2060[17]), .I2(n2027), 
            .I3(GND_net), .O(n2107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1420_3_lut (.I0(n2006), .I1(n2060[19]), .I2(n2027), 
            .I3(GND_net), .O(n2105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1414_3_lut (.I0(n2000), .I1(n2060[25]), .I2(n2027), 
            .I3(GND_net), .O(n2099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1415_3_lut (.I0(n2001), .I1(n2060[24]), .I2(n2027), 
            .I3(GND_net), .O(n2100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1424_3_lut (.I0(bit_ctr[15]), .I1(n2060[15]), .I2(n2027), 
            .I3(GND_net), .O(n2109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1423_3_lut (.I0(n2009), .I1(n2060[16]), .I2(n2027), 
            .I3(GND_net), .O(n2108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1417_3_lut (.I0(n2003), .I1(n2060[22]), .I2(n2027), 
            .I3(GND_net), .O(n2102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1421_3_lut (.I0(n2007), .I1(n2060[18]), .I2(n2027), 
            .I3(GND_net), .O(n2106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1409_3_lut (.I0(n1995), .I1(n2060[30]), .I2(n2027), 
            .I3(GND_net), .O(n2094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1546 (.I0(n2094), .I1(n2093), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5178));
    defparam i1_2_lut_adj_1546.LUT_INIT = 16'heeee;
    SB_LUT4 i22924_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n36606));
    defparam i22924_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1547 (.I0(n2106), .I1(n2102), .I2(n2108), .I3(n18_adj_5178), 
            .O(n30_adj_5179));
    defparam i13_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1548 (.I0(n2100), .I1(n2099), .I2(n36606), .I3(n2105), 
            .O(n28_adj_5180));
    defparam i11_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1549 (.I0(n2107), .I1(n2104), .I2(n2098), .I3(n2101), 
            .O(n29_adj_5181));
    defparam i12_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1550 (.I0(n2097), .I1(n2095), .I2(n2096), .I3(n2103), 
            .O(n27_adj_5182));
    defparam i10_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2188_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n41739));
    SB_LUT4 i16_4_lut_adj_1551 (.I0(n27_adj_5182), .I1(n29_adj_5181), .I2(n28_adj_5180), 
            .I3(n30_adj_5179), .O(n2126));
    defparam i16_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n30240));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n30239));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1344_3_lut (.I0(n1898), .I1(n1961[28]), .I2(n1928), 
            .I3(GND_net), .O(n1997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1343_3_lut (.I0(n1897), .I1(n1961[29]), .I2(n1928), 
            .I3(GND_net), .O(n1996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1342_3_lut (.I0(n1896), .I1(n1961[30]), .I2(n1928), 
            .I3(GND_net), .O(n1995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1342_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n30238));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n30237));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n30236));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1348_3_lut (.I0(n1902), .I1(n1961[24]), .I2(n1928), 
            .I3(GND_net), .O(n2001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1346_3_lut (.I0(n1900), .I1(n1961[26]), .I2(n1928), 
            .I3(GND_net), .O(n1999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1346_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n30235));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n30234));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n30233));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n30232));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1347_3_lut (.I0(n1901), .I1(n1961[25]), .I2(n1928), 
            .I3(GND_net), .O(n2000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1347_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n30231));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n30230));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1345_3_lut (.I0(n1899), .I1(n1961[27]), .I2(n1928), 
            .I3(GND_net), .O(n1998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1345_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n30229));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n30228));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n30227));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n30226));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n30225));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n30224));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n30223));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n30222));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n30221));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1354_3_lut (.I0(n1908), .I1(n1961[18]), .I2(n1928), 
            .I3(GND_net), .O(n2007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1349_3_lut (.I0(n1903), .I1(n1961[23]), .I2(n1928), 
            .I3(GND_net), .O(n2002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1355_3_lut (.I0(n1909), .I1(n1961[17]), .I2(n1928), 
            .I3(GND_net), .O(n2008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1356_3_lut (.I0(bit_ctr[16]), .I1(n1961[16]), .I2(n1928), 
            .I3(GND_net), .O(n2009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1353_3_lut (.I0(n1907), .I1(n1961[19]), .I2(n1928), 
            .I3(GND_net), .O(n2006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1352_3_lut (.I0(n1906), .I1(n1961[20]), .I2(n1928), 
            .I3(GND_net), .O(n2005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1351_3_lut (.I0(n1905), .I1(n1961[21]), .I2(n1928), 
            .I3(GND_net), .O(n2004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1350_3_lut (.I0(n1904), .I1(n1961[22]), .I2(n1928), 
            .I3(GND_net), .O(n2003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22922_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n36604));
    defparam i22922_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1552 (.I0(n2003), .I1(n2004), .I2(n2005), .I3(n2006), 
            .O(n28_adj_5183));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1553 (.I0(n1998), .I1(n2000), .I2(n1999), .I3(n2001), 
            .O(n26_adj_5184));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1554 (.I0(n2008), .I1(n36604), .I2(n2002), .I3(n2007), 
            .O(n27_adj_5185));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1995), .I1(n1996), .I2(n1994), .I3(n1997), 
            .O(n25_adj_5186));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1555 (.I0(n25_adj_5186), .I1(n27_adj_5185), .I2(n26_adj_5184), 
            .I3(n28_adj_5183), .O(n2027));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i22920_2_lut (.I0(bit_ctr[16]), .I1(n1909), .I2(GND_net), 
            .I3(GND_net), .O(n36602));
    defparam i22920_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut_adj_1556 (.I0(n1902), .I1(n1903), .I2(n1900), .I3(n1907), 
            .O(n26_adj_5187));
    defparam i11_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1557 (.I0(n1897), .I1(n36602), .I2(n1898), .I3(n1906), 
            .O(n24_adj_5188));
    defparam i9_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1558 (.I0(n1899), .I1(n1904), .I2(n1905), .I3(n1901), 
            .O(n25_adj_5189));
    defparam i10_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(n1908), .I1(n1896), .I2(n1895), .I3(GND_net), 
            .O(n23_adj_5190));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut_adj_1559 (.I0(n23_adj_5190), .I1(n25_adj_5189), .I2(n24_adj_5188), 
            .I3(n26_adj_5187), .O(n1928));
    defparam i14_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n51038), .I1(state[1]), .I2(n38580), .I3(GND_net), 
            .O(n12_adj_5191));   // verilog/neopixel.v(16[20:25])
    defparam i26_4_lut.LUT_INIT = 16'h7474;
    SB_LUT4 i37094_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n52729));
    defparam i37094_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n40466), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n40465), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_32 (.CI(n40465), .I0(bit_ctr[30]), .I1(GND_net), .CO(n40466));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n40464), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n40464), .I0(bit_ctr[29]), .I1(GND_net), .CO(n40465));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1136), .I1(n1103), .I2(VCC_net), 
            .I3(n41731), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_803_8_lut (.I0(GND_net), .I1(n1104), .I2(VCC_net), 
            .I3(n41730), .O(n1169[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_8 (.CI(n41730), .I0(n1104), .I1(VCC_net), .CO(n41731));
    SB_LUT4 mod_5_add_803_7_lut (.I0(GND_net), .I1(n1105), .I2(VCC_net), 
            .I3(n41729), .O(n1169[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_7 (.CI(n41729), .I0(n1105), .I1(VCC_net), .CO(n41730));
    SB_LUT4 mod_5_add_803_6_lut (.I0(GND_net), .I1(n1106), .I2(VCC_net), 
            .I3(n41728), .O(n1169[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_6 (.CI(n41728), .I0(n1106), .I1(VCC_net), .CO(n41729));
    SB_LUT4 mod_5_add_803_5_lut (.I0(GND_net), .I1(n1107), .I2(VCC_net), 
            .I3(n41727), .O(n1169[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_5 (.CI(n41727), .I0(n1107), .I1(VCC_net), .CO(n41728));
    SB_LUT4 mod_5_add_803_4_lut (.I0(GND_net), .I1(n1108), .I2(VCC_net), 
            .I3(n41726), .O(n1169[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_4 (.CI(n41726), .I0(n1108), .I1(VCC_net), .CO(n41727));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n40463), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n40463), .I0(bit_ctr[28]), .I1(GND_net), .CO(n40464));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n40462), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n40462), .I0(bit_ctr[27]), .I1(GND_net), .CO(n40463));
    SB_LUT4 mod_5_add_803_3_lut (.I0(GND_net), .I1(n1109), .I2(GND_net), 
            .I3(n41725), .O(n1169[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_3 (.CI(n41725), .I0(n1109), .I1(GND_net), .CO(n41726));
    SB_LUT4 mod_5_add_803_2_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(VCC_net), .O(n1169[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(GND_net), 
            .CO(n41725));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1334), .I1(n1301), .I2(VCC_net), 
            .I3(n41724), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_10_lut (.I0(GND_net), .I1(n1302), .I2(VCC_net), 
            .I3(n41723), .O(n1367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n41723), .I0(n1302), .I1(VCC_net), 
            .CO(n41724));
    SB_LUT4 mod_5_add_937_9_lut (.I0(GND_net), .I1(n1303), .I2(VCC_net), 
            .I3(n41722), .O(n1367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_9 (.CI(n41722), .I0(n1303), .I1(VCC_net), .CO(n41723));
    SB_LUT4 mod_5_add_937_8_lut (.I0(GND_net), .I1(n1304), .I2(VCC_net), 
            .I3(n41721), .O(n1367[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_8 (.CI(n41721), .I0(n1304), .I1(VCC_net), .CO(n41722));
    SB_DFFESS state_i0 (.Q(state[0]), .C(CLK_c), .E(n7_adj_5192), .D(state_3__N_528[0]), 
            .S(n38562));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_7_lut (.I0(GND_net), .I1(n1305), .I2(VCC_net), 
            .I3(n41720), .O(n1367[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n40461), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_7 (.CI(n41720), .I0(n1305), .I1(VCC_net), .CO(n41721));
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n29590), .D(n255[0]), 
            .R(n30005));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_6_lut (.I0(GND_net), .I1(n1306), .I2(VCC_net), 
            .I3(n41719), .O(n1367[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_6 (.CI(n41719), .I0(n1306), .I1(VCC_net), .CO(n41720));
    SB_LUT4 mod_5_add_937_5_lut (.I0(GND_net), .I1(n1307), .I2(VCC_net), 
            .I3(n41718), .O(n1367[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_5 (.CI(n41718), .I0(n1307), .I1(VCC_net), .CO(n41719));
    SB_CARRY add_21_28 (.CI(n40461), .I0(bit_ctr[26]), .I1(GND_net), .CO(n40462));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n40460), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_4_lut (.I0(GND_net), .I1(n1308), .I2(VCC_net), 
            .I3(n41717), .O(n1367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n41717), .I0(n1308), .I1(VCC_net), .CO(n41718));
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_3_lut (.I0(GND_net), .I1(n1309), .I2(GND_net), 
            .I3(n41716), .O(n1367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n41716), .I0(n1309), .I1(GND_net), .CO(n41717));
    SB_LUT4 mod_5_add_937_2_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(VCC_net), .O(n1367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(GND_net), 
            .CO(n41716));
    SB_LUT4 i36538_2_lut (.I0(n43736), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i36538_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n49915), .I1(timer[31]), .I2(n1[31]), 
            .I3(n40630), .O(n28470)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_27 (.CI(n40460), .I0(bit_ctr[25]), .I1(GND_net), .CO(n40461));
    SB_LUT4 i36536_2_lut (.I0(n43736), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i36536_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n49913), .I1(timer[30]), .I2(n1[30]), 
            .I3(n40629), .O(n49915)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n40629), .I0(timer[30]), .I1(n1[30]), 
            .CO(n40630));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n49911), .I1(timer[29]), .I2(n1[29]), 
            .I3(n40628), .O(n49913)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1235), .I1(n1202), .I2(VCC_net), 
            .I3(n42258), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_870_9_lut (.I0(GND_net), .I1(n1203), .I2(VCC_net), 
            .I3(n42257), .O(n1268[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_9 (.CI(n42257), .I0(n1203), .I1(VCC_net), .CO(n42258));
    SB_LUT4 mod_5_add_870_8_lut (.I0(GND_net), .I1(n1204), .I2(VCC_net), 
            .I3(n42256), .O(n1268[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_8 (.CI(n42256), .I0(n1204), .I1(VCC_net), .CO(n42257));
    SB_LUT4 mod_5_add_870_7_lut (.I0(GND_net), .I1(n1205), .I2(VCC_net), 
            .I3(n42255), .O(n1268[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_7 (.CI(n42255), .I0(n1205), .I1(VCC_net), .CO(n42256));
    SB_LUT4 mod_5_add_870_6_lut (.I0(GND_net), .I1(n1206), .I2(VCC_net), 
            .I3(n42254), .O(n1268[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_6 (.CI(n42254), .I0(n1206), .I1(VCC_net), .CO(n42255));
    SB_LUT4 mod_5_add_870_5_lut (.I0(GND_net), .I1(n1207), .I2(VCC_net), 
            .I3(n42253), .O(n1268[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_5 (.CI(n42253), .I0(n1207), .I1(VCC_net), .CO(n42254));
    SB_LUT4 mod_5_add_870_4_lut (.I0(GND_net), .I1(n1208), .I2(VCC_net), 
            .I3(n42252), .O(n1268[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_4 (.CI(n42252), .I0(n1208), .I1(VCC_net), .CO(n42253));
    SB_LUT4 mod_5_add_870_3_lut (.I0(GND_net), .I1(n1209), .I2(GND_net), 
            .I3(n42251), .O(n1268[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_3 (.CI(n42251), .I0(n1209), .I1(GND_net), .CO(n42252));
    SB_LUT4 mod_5_add_870_2_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(VCC_net), .O(n1268[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_31 (.CI(n40628), .I0(timer[29]), .I1(n1[29]), 
            .CO(n40629));
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(GND_net), 
            .CO(n42251));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1631), .I1(n1598), .I2(VCC_net), 
            .I3(n42250), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(GND_net), .I1(n1599), .I2(VCC_net), 
            .I3(n42249), .O(n1664[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_13 (.CI(n42249), .I0(n1599), .I1(VCC_net), 
            .CO(n42250));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(GND_net), .I1(n1600), .I2(VCC_net), 
            .I3(n42248), .O(n1664[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_12 (.CI(n42248), .I0(n1600), .I1(VCC_net), 
            .CO(n42249));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(GND_net), .I1(n1601), .I2(VCC_net), 
            .I3(n42247), .O(n1664[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_11 (.CI(n42247), .I0(n1601), .I1(VCC_net), 
            .CO(n42248));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(GND_net), .I1(n1602), .I2(VCC_net), 
            .I3(n42246), .O(n1664[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_10 (.CI(n42246), .I0(n1602), .I1(VCC_net), 
            .CO(n42247));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(GND_net), .I1(n1603), .I2(VCC_net), 
            .I3(n42245), .O(n1664[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_9 (.CI(n42245), .I0(n1603), .I1(VCC_net), 
            .CO(n42246));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(GND_net), .I1(n1604), .I2(VCC_net), 
            .I3(n42244), .O(n1664[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_8 (.CI(n42244), .I0(n1604), .I1(VCC_net), 
            .CO(n42245));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(GND_net), .I1(n1605), .I2(VCC_net), 
            .I3(n42243), .O(n1664[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_7 (.CI(n42243), .I0(n1605), .I1(VCC_net), 
            .CO(n42244));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(GND_net), .I1(n1606), .I2(VCC_net), 
            .I3(n42242), .O(n1664[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_6 (.CI(n42242), .I0(n1606), .I1(VCC_net), 
            .CO(n42243));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(GND_net), .I1(n1607), .I2(VCC_net), 
            .I3(n42241), .O(n1664[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_5 (.CI(n42241), .I0(n1607), .I1(VCC_net), 
            .CO(n42242));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(GND_net), .I1(n1608), .I2(VCC_net), 
            .I3(n42240), .O(n1664[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_4 (.CI(n42240), .I0(n1608), .I1(VCC_net), 
            .CO(n42241));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(GND_net), .I1(n1609), .I2(GND_net), 
            .I3(n42239), .O(n1664[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_3 (.CI(n42239), .I0(n1609), .I1(GND_net), 
            .CO(n42240));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(VCC_net), .O(n1664[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(GND_net), 
            .CO(n42239));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1730), .I1(n1697), .I2(VCC_net), 
            .I3(n42238), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(GND_net), .I1(n1698), .I2(VCC_net), 
            .I3(n42237), .O(n1763[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_14 (.CI(n42237), .I0(n1698), .I1(VCC_net), 
            .CO(n42238));
    SB_LUT4 mod_5_i1217_3_lut (.I0(n1707), .I1(n1763[21]), .I2(n1730), 
            .I3(GND_net), .O(n1806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1210_3_lut (.I0(n1700), .I1(n1763[28]), .I2(n1730), 
            .I3(GND_net), .O(n1799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1219_3_lut (.I0(n1709), .I1(n1763[19]), .I2(n1730), 
            .I3(GND_net), .O(n1808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1218_3_lut (.I0(n1708), .I1(n1763[20]), .I2(n1730), 
            .I3(GND_net), .O(n1807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1209_3_lut (.I0(n1699), .I1(n1763[29]), .I2(n1730), 
            .I3(GND_net), .O(n1798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1208_3_lut (.I0(n1698), .I1(n1763[30]), .I2(n1730), 
            .I3(GND_net), .O(n1797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1214_3_lut (.I0(n1704), .I1(n1763[24]), .I2(n1730), 
            .I3(GND_net), .O(n1803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1212_3_lut (.I0(n1702), .I1(n1763[26]), .I2(n1730), 
            .I3(GND_net), .O(n1801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1205_13_lut (.I0(GND_net), .I1(n1699), .I2(VCC_net), 
            .I3(n42236), .O(n1763[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_13 (.CI(n42236), .I0(n1699), .I1(VCC_net), 
            .CO(n42237));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(GND_net), .I1(n1700), .I2(VCC_net), 
            .I3(n42235), .O(n1763[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_12 (.CI(n42235), .I0(n1700), .I1(VCC_net), 
            .CO(n42236));
    SB_LUT4 mod_5_i1220_3_lut (.I0(bit_ctr[18]), .I1(n1763[18]), .I2(n1730), 
            .I3(GND_net), .O(n1809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(GND_net), .I1(n1701), .I2(VCC_net), 
            .I3(n42234), .O(n1763[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_11 (.CI(n42234), .I0(n1701), .I1(VCC_net), 
            .CO(n42235));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(GND_net), .I1(n1702), .I2(VCC_net), 
            .I3(n42233), .O(n1763[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n42233), .I0(n1702), .I1(VCC_net), 
            .CO(n42234));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(GND_net), .I1(n1703), .I2(VCC_net), 
            .I3(n42232), .O(n1763[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_9 (.CI(n42232), .I0(n1703), .I1(VCC_net), 
            .CO(n42233));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(GND_net), .I1(n1704), .I2(VCC_net), 
            .I3(n42231), .O(n1763[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_8 (.CI(n42231), .I0(n1704), .I1(VCC_net), 
            .CO(n42232));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(GND_net), .I1(n1705), .I2(VCC_net), 
            .I3(n42230), .O(n1763[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_7 (.CI(n42230), .I0(n1705), .I1(VCC_net), 
            .CO(n42231));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(GND_net), .I1(n1706), .I2(VCC_net), 
            .I3(n42229), .O(n1763[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_6 (.CI(n42229), .I0(n1706), .I1(VCC_net), 
            .CO(n42230));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(GND_net), .I1(n1707), .I2(VCC_net), 
            .I3(n42228), .O(n1763[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_5 (.CI(n42228), .I0(n1707), .I1(VCC_net), 
            .CO(n42229));
    SB_LUT4 mod_5_i1211_3_lut (.I0(n1701), .I1(n1763[27]), .I2(n1730), 
            .I3(GND_net), .O(n1800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(GND_net), .I1(n1708), .I2(VCC_net), 
            .I3(n42227), .O(n1763[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_4 (.CI(n42227), .I0(n1708), .I1(VCC_net), 
            .CO(n42228));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(GND_net), .I1(n1709), .I2(GND_net), 
            .I3(n42226), .O(n1763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n42226), .I0(n1709), .I1(GND_net), 
            .CO(n42227));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(VCC_net), .O(n1763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(GND_net), 
            .CO(n42226));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n42225), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n42224), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n42224), .I0(n1797), .I1(n1829), .CO(n42225));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n42223), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i1215_3_lut (.I0(n1705), .I1(n1763[23]), .I2(n1730), 
            .I3(GND_net), .O(n1804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1272_14 (.CI(n42223), .I0(n1798), .I1(n1829), .CO(n42224));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n42222), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n42222), .I0(n1799), .I1(n1829), .CO(n42223));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n42221), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n42221), .I0(n1800), .I1(n1829), .CO(n42222));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n42220), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n42220), .I0(n1801), .I1(n1829), .CO(n42221));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n42219), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n42219), .I0(n1802), .I1(n1829), .CO(n42220));
    SB_LUT4 mod_5_i1213_3_lut (.I0(n1703), .I1(n1763[25]), .I2(n1730), 
            .I3(GND_net), .O(n1802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n42218), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n42218), .I0(n1803), .I1(n1829), .CO(n42219));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n42217), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i1216_3_lut (.I0(n1706), .I1(n1763[22]), .I2(n1730), 
            .I3(GND_net), .O(n1805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1560 (.I0(n1805), .I1(n1802), .I2(n1804), .I3(n1796), 
            .O(n24_adj_5194));
    defparam i10_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1561 (.I0(bit_ctr[17]), .I1(n1800), .I2(n1809), 
            .I3(GND_net), .O(n17_adj_5195));
    defparam i3_3_lut_adj_1561.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1272_8 (.CI(n42217), .I0(n1804), .I1(n1829), .CO(n42218));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n42216), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n42216), .I0(n1805), .I1(n1829), .CO(n42217));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n49909), .I1(timer[28]), .I2(n1[28]), 
            .I3(n40627), .O(n49911)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i8_4_lut (.I0(n1801), .I1(n1803), .I2(n1797), .I3(n1798), 
            .O(n22_adj_5196));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_30 (.CI(n40627), .I0(timer[28]), .I1(n1[28]), 
            .CO(n40628));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n49907), .I1(timer[27]), .I2(n1[27]), 
            .I3(n40626), .O(n49909)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_4_lut_adj_1562 (.I0(n17_adj_5195), .I1(n24_adj_5194), .I2(n1807), 
            .I3(n1808), .O(n26_adj_5197));
    defparam i12_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n42215), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n42215), .I0(n1806), .I1(n1829), .CO(n42216));
    SB_LUT4 i13_4_lut_adj_1563 (.I0(n1799), .I1(n26_adj_5197), .I2(n22_adj_5196), 
            .I3(n1806), .O(n1829));
    defparam i13_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n42214), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n42214), .I0(n1807), .I1(n1829), .CO(n42215));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n42213), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n42213), .I0(n1808), .I1(n1829), .CO(n42214));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n52729), 
            .I3(n42212), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n42212), .I0(n1809), .I1(n52729), .CO(n42213));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n52729), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_29 (.CI(n40626), .I0(timer[27]), .I1(n1[27]), 
            .CO(n40627));
    SB_DFFE state_i1 (.Q(state[1]), .C(CLK_c), .E(VCC_net), .D(n12_adj_5191));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_2188__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n52729), 
            .CO(n42212));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1928), .I1(n1895), .I2(VCC_net), 
            .I3(n42211), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(GND_net), .I1(n1896), .I2(VCC_net), 
            .I3(n42210), .O(n1961[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n42210), .I0(n1896), .I1(VCC_net), 
            .CO(n42211));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(GND_net), .I1(n1897), .I2(VCC_net), 
            .I3(n42209), .O(n1961[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n42209), .I0(n1897), .I1(VCC_net), 
            .CO(n42210));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(GND_net), .I1(n1898), .I2(VCC_net), 
            .I3(n42208), .O(n1961[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_14 (.CI(n42208), .I0(n1898), .I1(VCC_net), 
            .CO(n42209));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(GND_net), .I1(n1899), .I2(VCC_net), 
            .I3(n42207), .O(n1961[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_13 (.CI(n42207), .I0(n1899), .I1(VCC_net), 
            .CO(n42208));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(GND_net), .I1(n1900), .I2(VCC_net), 
            .I3(n42206), .O(n1961[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n42206), .I0(n1900), .I1(VCC_net), 
            .CO(n42207));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(GND_net), .I1(n1901), .I2(VCC_net), 
            .I3(n42205), .O(n1961[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n52930));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY mod_5_add_1339_11 (.CI(n42205), .I0(n1901), .I1(VCC_net), 
            .CO(n42206));
    SB_LUT4 n52930_bdd_4_lut (.I0(n52930), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n50183));
    defparam n52930_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(GND_net), .I1(n1902), .I2(VCC_net), 
            .I3(n42204), .O(n1961[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_10 (.CI(n42204), .I0(n1902), .I1(VCC_net), 
            .CO(n42205));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(GND_net), .I1(n1903), .I2(VCC_net), 
            .I3(n42203), .O(n1961[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_9 (.CI(n42203), .I0(n1903), .I1(VCC_net), 
            .CO(n42204));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(GND_net), .I1(n1904), .I2(VCC_net), 
            .I3(n42202), .O(n1961[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n42202), .I0(n1904), .I1(VCC_net), 
            .CO(n42203));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(GND_net), .I1(n1905), .I2(VCC_net), 
            .I3(n42201), .O(n1961[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_7 (.CI(n42201), .I0(n1905), .I1(VCC_net), 
            .CO(n42202));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(GND_net), .I1(n1906), .I2(VCC_net), 
            .I3(n42200), .O(n1961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_6 (.CI(n42200), .I0(n1906), .I1(VCC_net), 
            .CO(n42201));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(GND_net), .I1(n1907), .I2(VCC_net), 
            .I3(n42199), .O(n1961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_5 (.CI(n42199), .I0(n1907), .I1(VCC_net), 
            .CO(n42200));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(GND_net), .I1(n1908), .I2(VCC_net), 
            .I3(n42198), .O(n1961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_4 (.CI(n42198), .I0(n1908), .I1(VCC_net), 
            .CO(n42199));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(GND_net), .I1(n1909), .I2(GND_net), 
            .I3(n42197), .O(n1961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_3 (.CI(n42197), .I0(n1909), .I1(GND_net), 
            .CO(n42198));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(VCC_net), .O(n1961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(GND_net), 
            .CO(n42197));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n2027), .I1(n1994), .I2(VCC_net), 
            .I3(n42196), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 bit_ctr_0__bdd_4_lut_37257 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n52888));
    defparam bit_ctr_0__bdd_4_lut_37257.LUT_INIT = 16'he4aa;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(GND_net), .I1(n1995), .I2(VCC_net), 
            .I3(n42195), .O(n2060[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n52888_bdd_4_lut (.I0(n52888), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n50261));
    defparam n52888_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY mod_5_add_1406_17 (.CI(n42195), .I0(n1995), .I1(VCC_net), 
            .CO(n42196));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(GND_net), .I1(n1996), .I2(VCC_net), 
            .I3(n42194), .O(n2060[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n42194), .I0(n1996), .I1(VCC_net), 
            .CO(n42195));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(GND_net), .I1(n1997), .I2(VCC_net), 
            .I3(n42193), .O(n2060[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_15 (.CI(n42193), .I0(n1997), .I1(VCC_net), 
            .CO(n42194));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(GND_net), .I1(n1998), .I2(VCC_net), 
            .I3(n42192), .O(n2060[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n42192), .I0(n1998), .I1(VCC_net), 
            .CO(n42193));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(GND_net), .I1(n1999), .I2(VCC_net), 
            .I3(n42191), .O(n2060[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_13 (.CI(n42191), .I0(n1999), .I1(VCC_net), 
            .CO(n42192));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(GND_net), .I1(n2000), .I2(VCC_net), 
            .I3(n42190), .O(n2060[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n42190), .I0(n2000), .I1(VCC_net), 
            .CO(n42191));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(GND_net), .I1(n2001), .I2(VCC_net), 
            .I3(n42189), .O(n2060[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n42189), .I0(n2001), .I1(VCC_net), 
            .CO(n42190));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(GND_net), .I1(n2002), .I2(VCC_net), 
            .I3(n42188), .O(n2060[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_10 (.CI(n42188), .I0(n2002), .I1(VCC_net), 
            .CO(n42189));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(GND_net), .I1(n2003), .I2(VCC_net), 
            .I3(n42187), .O(n2060[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_9 (.CI(n42187), .I0(n2003), .I1(VCC_net), 
            .CO(n42188));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(GND_net), .I1(n2004), .I2(VCC_net), 
            .I3(n42186), .O(n2060[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_8 (.CI(n42186), .I0(n2004), .I1(VCC_net), 
            .CO(n42187));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(GND_net), .I1(n2005), .I2(VCC_net), 
            .I3(n42185), .O(n2060[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n42185), .I0(n2005), .I1(VCC_net), 
            .CO(n42186));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(GND_net), .I1(n2006), .I2(VCC_net), 
            .I3(n42184), .O(n2060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_6 (.CI(n42184), .I0(n2006), .I1(VCC_net), 
            .CO(n42185));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(GND_net), .I1(n2007), .I2(VCC_net), 
            .I3(n42183), .O(n2060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n42183), .I0(n2007), .I1(VCC_net), 
            .CO(n42184));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(GND_net), .I1(n2008), .I2(VCC_net), 
            .I3(n42182), .O(n2060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_4 (.CI(n42182), .I0(n2008), .I1(VCC_net), 
            .CO(n42183));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(GND_net), .I1(n2009), .I2(GND_net), 
            .I3(n42181), .O(n2060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_28_lut (.I0(n49905), .I1(timer[26]), .I2(n1[26]), 
            .I3(n40625), .O(n49907)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n40459), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_3 (.CI(n42181), .I0(n2009), .I1(GND_net), 
            .CO(n42182));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(VCC_net), .O(n2060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(GND_net), 
            .CO(n42181));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2126), .I1(n2093), .I2(VCC_net), 
            .I3(n42180), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(GND_net), .I1(n2094), .I2(VCC_net), 
            .I3(n42179), .O(n2159[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_18 (.CI(n42179), .I0(n2094), .I1(VCC_net), 
            .CO(n42180));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(GND_net), .I1(n2095), .I2(VCC_net), 
            .I3(n42178), .O(n2159[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_17 (.CI(n42178), .I0(n2095), .I1(VCC_net), 
            .CO(n42179));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(GND_net), .I1(n2096), .I2(VCC_net), 
            .I3(n42177), .O(n2159[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n42177), .I0(n2096), .I1(VCC_net), 
            .CO(n42178));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(GND_net), .I1(n2097), .I2(VCC_net), 
            .I3(n42176), .O(n2159[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n42176), .I0(n2097), .I1(VCC_net), 
            .CO(n42177));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(GND_net), .I1(n2098), .I2(VCC_net), 
            .I3(n42175), .O(n2159[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n42175), .I0(n2098), .I1(VCC_net), 
            .CO(n42176));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(GND_net), .I1(n2099), .I2(VCC_net), 
            .I3(n42174), .O(n2159[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n42174), .I0(n2099), .I1(VCC_net), 
            .CO(n42175));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(GND_net), .I1(n2100), .I2(VCC_net), 
            .I3(n42173), .O(n2159[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_12 (.CI(n42173), .I0(n2100), .I1(VCC_net), 
            .CO(n42174));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(GND_net), .I1(n2101), .I2(VCC_net), 
            .I3(n42172), .O(n2159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n42172), .I0(n2101), .I1(VCC_net), 
            .CO(n42173));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(GND_net), .I1(n2102), .I2(VCC_net), 
            .I3(n42171), .O(n2159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n42171), .I0(n2102), .I1(VCC_net), 
            .CO(n42172));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(GND_net), .I1(n2103), .I2(VCC_net), 
            .I3(n42170), .O(n2159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_9 (.CI(n42170), .I0(n2103), .I1(VCC_net), 
            .CO(n42171));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(GND_net), .I1(n2104), .I2(VCC_net), 
            .I3(n42169), .O(n2159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_8 (.CI(n42169), .I0(n2104), .I1(VCC_net), 
            .CO(n42170));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(GND_net), .I1(n2105), .I2(VCC_net), 
            .I3(n42168), .O(n2159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n42168), .I0(n2105), .I1(VCC_net), 
            .CO(n42169));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(GND_net), .I1(n2106), .I2(VCC_net), 
            .I3(n42167), .O(n2159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n40625), .I0(timer[26]), .I1(n1[26]), 
            .CO(n40626));
    SB_CARRY mod_5_add_1473_6 (.CI(n42167), .I0(n2106), .I1(VCC_net), 
            .CO(n42168));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(GND_net), .I1(n2107), .I2(VCC_net), 
            .I3(n42166), .O(n2159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_5 (.CI(n42166), .I0(n2107), .I1(VCC_net), 
            .CO(n42167));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(GND_net), .I1(n2108), .I2(VCC_net), 
            .I3(n42165), .O(n2159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_4 (.CI(n42165), .I0(n2108), .I1(VCC_net), 
            .CO(n42166));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(GND_net), .I1(n2109), .I2(GND_net), 
            .I3(n42164), .O(n2159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_3 (.CI(n42164), .I0(n2109), .I1(GND_net), 
            .CO(n42165));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(VCC_net), .O(n2159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(GND_net), 
            .CO(n42164));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2225), .I1(n2192), .I2(VCC_net), 
            .I3(n42163), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(GND_net), .I1(n2193), .I2(VCC_net), 
            .I3(n42162), .O(n2258[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_19 (.CI(n42162), .I0(n2193), .I1(VCC_net), 
            .CO(n42163));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(GND_net), .I1(n2194), .I2(VCC_net), 
            .I3(n42161), .O(n2258[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_18 (.CI(n42161), .I0(n2194), .I1(VCC_net), 
            .CO(n42162));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(GND_net), .I1(n2195), .I2(VCC_net), 
            .I3(n42160), .O(n2258[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_17 (.CI(n42160), .I0(n2195), .I1(VCC_net), 
            .CO(n42161));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(GND_net), .I1(n2196), .I2(VCC_net), 
            .I3(n42159), .O(n2258[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_16 (.CI(n42159), .I0(n2196), .I1(VCC_net), 
            .CO(n42160));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(GND_net), .I1(n2197), .I2(VCC_net), 
            .I3(n42158), .O(n2258[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_15 (.CI(n42158), .I0(n2197), .I1(VCC_net), 
            .CO(n42159));
    SB_LUT4 sub_14_add_2_27_lut (.I0(n49903), .I1(timer[25]), .I2(n1[25]), 
            .I3(n40624), .O(n49905)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i36398_4_lut (.I0(n807), .I1(n838), .I2(n12165), .I3(n46352), 
            .O(n50068));
    defparam i36398_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mod_5_i605_4_lut (.I0(n807), .I1(n46352), .I2(n838), .I3(n12165), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_4_lut.LUT_INIT = 16'haaa9;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(GND_net), .I1(n2198), .I2(VCC_net), 
            .I3(n42157), .O(n2258[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_14 (.CI(n42157), .I0(n2198), .I1(VCC_net), 
            .CO(n42158));
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n43736), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n43736), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(GND_net), .I1(n2199), .I2(VCC_net), 
            .I3(n42156), .O(n2258[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_13 (.CI(n42156), .I0(n2199), .I1(VCC_net), 
            .CO(n42157));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(GND_net), .I1(n2200), .I2(VCC_net), 
            .I3(n42155), .O(n2258[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_12 (.CI(n42155), .I0(n2200), .I1(VCC_net), 
            .CO(n42156));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(GND_net), .I1(n2201), .I2(VCC_net), 
            .I3(n42154), .O(n2258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_11 (.CI(n42154), .I0(n2201), .I1(VCC_net), 
            .CO(n42155));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(GND_net), .I1(n2202), .I2(VCC_net), 
            .I3(n42153), .O(n2258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i675_3_lut (.I0(n26840), .I1(n971[27]), .I2(n43736), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n26854));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i34471_4_lut (.I0(n36796), .I1(bit_ctr[29]), .I2(bit_ctr[28]), 
            .I3(n739), .O(n46352));   // verilog/neopixel.v(22[26:36])
    defparam i34471_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n46742), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[31]), .I2(bit_ctr[30]), 
            .I3(GND_net), .O(n13435));   // verilog/neopixel.v(22[26:36])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i22769_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i22769_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_1540_10 (.CI(n42153), .I0(n2202), .I1(VCC_net), 
            .CO(n42154));
    SB_LUT4 bit_ctr_0__bdd_4_lut_37223 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n52882));
    defparam bit_ctr_0__bdd_4_lut_37223.LUT_INIT = 16'he4aa;
    SB_CARRY sub_14_add_2_27 (.CI(n40624), .I0(timer[25]), .I1(n1[25]), 
            .CO(n40625));
    SB_LUT4 i30760_rep_4_3_lut (.I0(bit_ctr[28]), .I1(bit_ctr[29]), .I2(n36796), 
            .I3(GND_net), .O(n46742));
    defparam i30760_rep_4_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(GND_net), .I1(n2203), .I2(VCC_net), 
            .I3(n42152), .O(n2258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35781_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[29]), .I2(bit_ctr[31]), 
            .I3(n36796), .O(n708));
    defparam i35781_4_lut.LUT_INIT = 16'hc60a;
    SB_CARRY mod_5_add_1540_9 (.CI(n42152), .I0(n2203), .I1(VCC_net), 
            .CO(n42153));
    SB_LUT4 i1_4_lut_adj_1565 (.I0(n708), .I1(n46742), .I2(n608), .I3(n13435), 
            .O(n739));
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'h0111;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(n807), .I1(n46352), .I2(bit_ctr[27]), 
            .I3(n26854), .O(n838));
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'h1101;
    SB_LUT4 i1_2_lut_adj_1567 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n26840));
    defparam i1_2_lut_adj_1567.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(GND_net), .I1(n2204), .I2(VCC_net), 
            .I3(n42151), .O(n2258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n42151), .I0(n2204), .I1(VCC_net), 
            .CO(n42152));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n49901), .I1(timer[24]), .I2(n1[24]), 
            .I3(n40623), .O(n49903)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_26 (.CI(n40459), .I0(bit_ctr[24]), .I1(GND_net), .CO(n40460));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(GND_net), .I1(n2205), .I2(VCC_net), 
            .I3(n42150), .O(n2258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34372_4_lut (.I0(n739), .I1(bit_ctr[28]), .I2(bit_ctr[27]), 
            .I3(n838), .O(n29881));   // verilog/neopixel.v(22[26:36])
    defparam i34372_4_lut.LUT_INIT = 16'h9969;
    SB_CARRY mod_5_add_1540_7 (.CI(n42150), .I0(n2205), .I1(VCC_net), 
            .CO(n42151));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(GND_net), .I1(n2206), .I2(VCC_net), 
            .I3(n42149), .O(n2258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n42149), .I0(n2206), .I1(VCC_net), 
            .CO(n42150));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(GND_net), .I1(n2207), .I2(VCC_net), 
            .I3(n42148), .O(n2258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_5 (.CI(n42148), .I0(n2207), .I1(VCC_net), 
            .CO(n42149));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(GND_net), .I1(n2208), .I2(VCC_net), 
            .I3(n42147), .O(n2258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1568 (.I0(n50068), .I1(n46442), .I2(n906), .I3(n49527), 
            .O(n43736));
    defparam i1_4_lut_adj_1568.LUT_INIT = 16'h0100;
    SB_CARRY mod_5_add_1540_4 (.CI(n42147), .I0(n2208), .I1(VCC_net), 
            .CO(n42148));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(GND_net), .I1(n2209), .I2(GND_net), 
            .I3(n42146), .O(n2258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n40458), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n42146), .I0(n2209), .I1(GND_net), 
            .CO(n42147));
    SB_LUT4 i30870_3_lut (.I0(n43736), .I1(n971[28]), .I2(n971[29]), .I3(GND_net), 
            .O(n46437));
    defparam i30870_3_lut.LUT_INIT = 16'habab;
    SB_CARRY sub_14_add_2_26 (.CI(n40623), .I0(timer[24]), .I1(n1[24]), 
            .CO(n40624));
    SB_LUT4 i2_3_lut (.I0(n1005), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n7_adj_5198));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5198), .I1(n1008), .I2(n46437), .I3(n4), 
            .O(n1037));
    defparam i4_4_lut.LUT_INIT = 16'hffef;
    SB_CARRY add_21_25 (.CI(n40458), .I0(bit_ctr[23]), .I1(GND_net), .CO(n40459));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(VCC_net), .O(n2258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(GND_net), 
            .CO(n42146));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n49899), .I1(timer[23]), .I2(n1[23]), 
            .I3(n40622), .O(n49901)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2324), .I1(n2291), .I2(VCC_net), 
            .I3(n42145), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(GND_net), .I1(n2292), .I2(VCC_net), 
            .I3(n42144), .O(n2357[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n40457), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_25 (.CI(n40622), .I0(timer[23]), .I1(n1[23]), 
            .CO(n40623));
    SB_CARRY mod_5_add_1607_20 (.CI(n42144), .I0(n2292), .I1(VCC_net), 
            .CO(n42145));
    SB_LUT4 mod_5_add_669_7_lut (.I0(n52230), .I1(n50068), .I2(VCC_net), 
            .I3(n40704), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_19_lut (.I0(GND_net), .I1(n2293), .I2(VCC_net), 
            .I3(n42143), .O(n2357[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_19 (.CI(n42143), .I0(n2293), .I1(VCC_net), 
            .CO(n42144));
    SB_CARRY add_21_24 (.CI(n40457), .I0(bit_ctr[22]), .I1(GND_net), .CO(n40458));
    SB_LUT4 n52882_bdd_4_lut (.I0(n52882), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n50267));
    defparam n52882_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1607_18_lut (.I0(GND_net), .I1(n2294), .I2(VCC_net), 
            .I3(n42142), .O(n2357[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_18 (.CI(n42142), .I0(n2294), .I1(VCC_net), 
            .CO(n42143));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(GND_net), .I1(n2295), .I2(VCC_net), 
            .I3(n42141), .O(n2357[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n42141), .I0(n2295), .I1(VCC_net), 
            .CO(n42142));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(GND_net), .I1(n2296), .I2(VCC_net), 
            .I3(n42140), .O(n2357[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n42140), .I0(n2296), .I1(VCC_net), 
            .CO(n42141));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n40456), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(GND_net), .I1(n2297), .I2(VCC_net), 
            .I3(n42139), .O(n2357[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n40456), .I0(bit_ctr[21]), .I1(GND_net), .CO(n40457));
    SB_CARRY mod_5_add_1607_15 (.CI(n42139), .I0(n2297), .I1(VCC_net), 
            .CO(n42140));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(GND_net), .I1(n2298), .I2(VCC_net), 
            .I3(n42138), .O(n2357[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n42138), .I0(n2298), .I1(VCC_net), 
            .CO(n42139));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(GND_net), .I1(n2299), .I2(VCC_net), 
            .I3(n42137), .O(n2357[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_13 (.CI(n42137), .I0(n2299), .I1(VCC_net), 
            .CO(n42138));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n49897), .I1(timer[22]), .I2(n1[22]), 
            .I3(n40621), .O(n49899)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(GND_net), .I1(n2300), .I2(VCC_net), 
            .I3(n42136), .O(n2357[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_12 (.CI(n42136), .I0(n2300), .I1(VCC_net), 
            .CO(n42137));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(GND_net), .I1(n2301), .I2(VCC_net), 
            .I3(n42135), .O(n2357[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n42135), .I0(n2301), .I1(VCC_net), 
            .CO(n42136));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(GND_net), .I1(n2302), .I2(VCC_net), 
            .I3(n42134), .O(n2357[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n42134), .I0(n2302), .I1(VCC_net), 
            .CO(n42135));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(GND_net), .I1(n2303), .I2(VCC_net), 
            .I3(n42133), .O(n2357[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_9 (.CI(n42133), .I0(n2303), .I1(VCC_net), 
            .CO(n42134));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(GND_net), .I1(n2304), .I2(VCC_net), 
            .I3(n42132), .O(n2357[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n40455), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n40703), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n40703), .I0(n906), .I1(VCC_net), .CO(n40704));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n46442), .I2(VCC_net), 
            .I3(n40702), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n40702), .I0(n46442), .I1(VCC_net), 
            .CO(n40703));
    SB_CARRY mod_5_add_1607_8 (.CI(n42132), .I0(n2304), .I1(VCC_net), 
            .CO(n42133));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n29881), .I2(VCC_net), 
            .I3(n40701), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(GND_net), .I1(n2305), .I2(VCC_net), 
            .I3(n42131), .O(n2357[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_7 (.CI(n42131), .I0(n2305), .I1(VCC_net), 
            .CO(n42132));
    SB_CARRY mod_5_add_669_4 (.CI(n40701), .I0(n29881), .I1(VCC_net), 
            .CO(n40702));
    SB_CARRY sub_14_add_2_24 (.CI(n40621), .I0(timer[22]), .I1(n1[22]), 
            .CO(n40622));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n49895), .I1(timer[21]), .I2(n1[21]), 
            .I3(n40620), .O(n49897)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n26840), .I2(GND_net), 
            .I3(n40700), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_6_lut (.I0(GND_net), .I1(n2306), .I2(VCC_net), 
            .I3(n42130), .O(n2357[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_6 (.CI(n42130), .I0(n2306), .I1(VCC_net), 
            .CO(n42131));
    SB_CARRY sub_14_add_2_23 (.CI(n40620), .I0(timer[21]), .I1(n1[21]), 
            .CO(n40621));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(GND_net), .I1(n2307), .I2(VCC_net), 
            .I3(n42129), .O(n2357[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_5 (.CI(n42129), .I0(n2307), .I1(VCC_net), 
            .CO(n42130));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(GND_net), .I1(n2308), .I2(VCC_net), 
            .I3(n42128), .O(n2357[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n42128), .I0(n2308), .I1(VCC_net), 
            .CO(n42129));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(GND_net), .I1(n2309), .I2(GND_net), 
            .I3(n42127), .O(n2357[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_22_lut (.I0(n49893), .I1(timer[20]), .I2(n1[20]), 
            .I3(n40619), .O(n49895)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1607_3 (.CI(n42127), .I0(n2309), .I1(GND_net), 
            .CO(n42128));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(VCC_net), .O(n2357[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_22 (.CI(n40619), .I0(timer[20]), .I1(n1[20]), 
            .CO(n40620));
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(GND_net), 
            .CO(n42127));
    SB_LUT4 sub_14_add_2_21_lut (.I0(n49891), .I1(timer[19]), .I2(n1[19]), 
            .I3(n40618), .O(n49893)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_22 (.CI(n40455), .I0(bit_ctr[20]), .I1(GND_net), .CO(n40456));
    SB_CARRY mod_5_add_669_3 (.CI(n40700), .I0(n26840), .I1(GND_net), 
            .CO(n40701));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2423), .I1(n2390), .I2(VCC_net), 
            .I3(n42126), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(GND_net), .I1(n2391), .I2(VCC_net), 
            .I3(n42125), .O(n2456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n42125), .I0(n2391), .I1(VCC_net), 
            .CO(n42126));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(GND_net), .I1(n2392), .I2(VCC_net), 
            .I3(n42124), .O(n2456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n42124), .I0(n2392), .I1(VCC_net), 
            .CO(n42125));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n40454), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_19_lut (.I0(GND_net), .I1(n2393), .I2(VCC_net), 
            .I3(n42123), .O(n2456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_19 (.CI(n42123), .I0(n2393), .I1(VCC_net), 
            .CO(n42124));
    SB_CARRY sub_14_add_2_21 (.CI(n40618), .I0(timer[19]), .I1(n1[19]), 
            .CO(n40619));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(GND_net), .I1(n2394), .I2(VCC_net), 
            .I3(n42122), .O(n2456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_21 (.CI(n40454), .I0(bit_ctr[19]), .I1(GND_net), .CO(n40455));
    SB_CARRY mod_5_add_1674_18 (.CI(n42122), .I0(n2394), .I1(VCC_net), 
            .CO(n42123));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(GND_net), .I1(n2395), .I2(VCC_net), 
            .I3(n42121), .O(n2456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_17 (.CI(n42121), .I0(n2395), .I1(VCC_net), 
            .CO(n42122));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(GND_net), .I1(n2396), .I2(VCC_net), 
            .I3(n42120), .O(n2456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n42120), .I0(n2396), .I1(VCC_net), 
            .CO(n42121));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(GND_net), .I1(n2397), .I2(VCC_net), 
            .I3(n42119), .O(n2456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_15 (.CI(n42119), .I0(n2397), .I1(VCC_net), 
            .CO(n42120));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_14_lut (.I0(GND_net), .I1(n2398), .I2(VCC_net), 
            .I3(n42118), .O(n2456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n40700));
    SB_CARRY mod_5_add_1674_14 (.CI(n42118), .I0(n2398), .I1(VCC_net), 
            .CO(n42119));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n49889), .I1(timer[18]), .I2(n1[18]), 
            .I3(n40617), .O(n49891)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_13_lut (.I0(GND_net), .I1(n2399), .I2(VCC_net), 
            .I3(n42117), .O(n2456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n40453), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n42117), .I0(n2399), .I1(VCC_net), 
            .CO(n42118));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(GND_net), .I1(n2400), .I2(VCC_net), 
            .I3(n42116), .O(n2456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n40617), .I0(timer[18]), .I1(n1[18]), 
            .CO(n40618));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n49887), .I1(timer[17]), .I2(n1[17]), 
            .I3(n40616), .O(n49889)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1674_12 (.CI(n42116), .I0(n2400), .I1(VCC_net), 
            .CO(n42117));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(GND_net), .I1(n2401), .I2(VCC_net), 
            .I3(n42115), .O(n2456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n40453), .I0(bit_ctr[18]), .I1(GND_net), .CO(n40454));
    SB_CARRY mod_5_add_1674_11 (.CI(n42115), .I0(n2401), .I1(VCC_net), 
            .CO(n42116));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(GND_net), .I1(n2402), .I2(VCC_net), 
            .I3(n42114), .O(n2456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n40452), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_10 (.CI(n42114), .I0(n2402), .I1(VCC_net), 
            .CO(n42115));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(GND_net), .I1(n2403), .I2(VCC_net), 
            .I3(n42113), .O(n2456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n42113), .I0(n2403), .I1(VCC_net), 
            .CO(n42114));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(GND_net), .I1(n2404), .I2(VCC_net), 
            .I3(n42112), .O(n2456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_19 (.CI(n40616), .I0(timer[17]), .I1(n1[17]), 
            .CO(n40617));
    SB_CARRY mod_5_add_1674_8 (.CI(n42112), .I0(n2404), .I1(VCC_net), 
            .CO(n42113));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(GND_net), .I1(n2405), .I2(VCC_net), 
            .I3(n42111), .O(n2456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_7 (.CI(n42111), .I0(n2405), .I1(VCC_net), 
            .CO(n42112));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(GND_net), .I1(n2406), .I2(VCC_net), 
            .I3(n42110), .O(n2456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_6 (.CI(n42110), .I0(n2406), .I1(VCC_net), 
            .CO(n42111));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(GND_net), .I1(n2407), .I2(VCC_net), 
            .I3(n42109), .O(n2456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_5 (.CI(n42109), .I0(n2407), .I1(VCC_net), 
            .CO(n42110));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n49885), .I1(timer[16]), .I2(n1[16]), 
            .I3(n40615), .O(n49887)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(GND_net), .I1(n2408), .I2(VCC_net), 
            .I3(n42108), .O(n2456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_4 (.CI(n42108), .I0(n2408), .I1(VCC_net), 
            .CO(n42109));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(GND_net), .I1(n2409), .I2(GND_net), 
            .I3(n42107), .O(n2456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_3 (.CI(n42107), .I0(n2409), .I1(GND_net), 
            .CO(n42108));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(VCC_net), .O(n2456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(GND_net), 
            .CO(n42107));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2522), .I1(n2489), .I2(VCC_net), 
            .I3(n42106), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(GND_net), .I1(n2490), .I2(VCC_net), 
            .I3(n42105), .O(n2555[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_22 (.CI(n42105), .I0(n2490), .I1(VCC_net), 
            .CO(n42106));
    SB_CARRY sub_14_add_2_18 (.CI(n40615), .I0(timer[16]), .I1(n1[16]), 
            .CO(n40616));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(GND_net), .I1(n2491), .I2(VCC_net), 
            .I3(n42104), .O(n2555[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_17_lut (.I0(n49883), .I1(timer[15]), .I2(n1[15]), 
            .I3(n40614), .O(n49885)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_17 (.CI(n40614), .I0(timer[15]), .I1(n1[15]), 
            .CO(n40615));
    SB_CARRY mod_5_add_1741_21 (.CI(n42104), .I0(n2491), .I1(VCC_net), 
            .CO(n42105));
    SB_LUT4 sub_14_add_2_16_lut (.I0(n49881), .I1(timer[14]), .I2(n1[14]), 
            .I3(n40613), .O(n49883)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(GND_net), .I1(n2492), .I2(VCC_net), 
            .I3(n42103), .O(n2555[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_20 (.CI(n42103), .I0(n2492), .I1(VCC_net), 
            .CO(n42104));
    SB_CARRY sub_14_add_2_16 (.CI(n40613), .I0(timer[14]), .I1(n1[14]), 
            .CO(n40614));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(GND_net), .I1(n2493), .I2(VCC_net), 
            .I3(n42102), .O(n2555[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n40452), .I0(bit_ctr[17]), .I1(GND_net), .CO(n40453));
    SB_CARRY mod_5_add_1741_19 (.CI(n42102), .I0(n2493), .I1(VCC_net), 
            .CO(n42103));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(GND_net), .I1(n2494), .I2(VCC_net), 
            .I3(n42101), .O(n2555[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_18 (.CI(n42101), .I0(n2494), .I1(VCC_net), 
            .CO(n42102));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(GND_net), .I1(n2495), .I2(VCC_net), 
            .I3(n42100), .O(n2555[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_17 (.CI(n42100), .I0(n2495), .I1(VCC_net), 
            .CO(n42101));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(GND_net), .I1(n2496), .I2(VCC_net), 
            .I3(n42099), .O(n2555[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n42099), .I0(n2496), .I1(VCC_net), 
            .CO(n42100));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(GND_net), .I1(n2497), .I2(VCC_net), 
            .I3(n42098), .O(n2555[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_15 (.CI(n42098), .I0(n2497), .I1(VCC_net), 
            .CO(n42099));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(GND_net), .I1(n2498), .I2(VCC_net), 
            .I3(n42097), .O(n2555[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_14 (.CI(n42097), .I0(n2498), .I1(VCC_net), 
            .CO(n42098));
    SB_LUT4 mod_5_i1146_3_lut (.I0(n1604), .I1(n1664[25]), .I2(n1631), 
            .I3(GND_net), .O(n1703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1147_3_lut (.I0(n1605), .I1(n1664[24]), .I2(n1631), 
            .I3(GND_net), .O(n1704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1148_3_lut (.I0(n1606), .I1(n1664[23]), .I2(n1631), 
            .I3(GND_net), .O(n1705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_15_lut (.I0(n49879), .I1(timer[13]), .I2(n1[13]), 
            .I3(n40612), .O(n49881)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1151_3_lut (.I0(n1609), .I1(n1664[20]), .I2(n1631), 
            .I3(GND_net), .O(n1708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_13_lut (.I0(GND_net), .I1(n2499), .I2(VCC_net), 
            .I3(n42096), .O(n2555[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1141_3_lut (.I0(n1599), .I1(n1664[30]), .I2(n1631), 
            .I3(GND_net), .O(n1698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_13 (.CI(n42096), .I0(n2499), .I1(VCC_net), 
            .CO(n42097));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(GND_net), .I1(n2500), .I2(VCC_net), 
            .I3(n42095), .O(n2555[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_12 (.CI(n42095), .I0(n2500), .I1(VCC_net), 
            .CO(n42096));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(GND_net), .I1(n2501), .I2(VCC_net), 
            .I3(n42094), .O(n2555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1150_3_lut (.I0(n1608), .I1(n1664[21]), .I2(n1631), 
            .I3(GND_net), .O(n1707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1150_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_11 (.CI(n42094), .I0(n2501), .I1(VCC_net), 
            .CO(n42095));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(GND_net), .I1(n2502), .I2(VCC_net), 
            .I3(n42093), .O(n2555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_10 (.CI(n42093), .I0(n2502), .I1(VCC_net), 
            .CO(n42094));
    SB_LUT4 mod_5_i1143_3_lut (.I0(n1601), .I1(n1664[28]), .I2(n1631), 
            .I3(GND_net), .O(n1700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(GND_net), .I1(n2503), .I2(VCC_net), 
            .I3(n42092), .O(n2555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1142_3_lut (.I0(n1600), .I1(n1664[29]), .I2(n1631), 
            .I3(GND_net), .O(n1699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_9 (.CI(n42092), .I0(n2503), .I1(VCC_net), 
            .CO(n42093));
    SB_CARRY sub_14_add_2_15 (.CI(n40612), .I0(timer[13]), .I1(n1[13]), 
            .CO(n40613));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(GND_net), .I1(n2504), .I2(VCC_net), 
            .I3(n42091), .O(n2555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n42091), .I0(n2504), .I1(VCC_net), 
            .CO(n42092));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(GND_net), .I1(n2505), .I2(VCC_net), 
            .I3(n42090), .O(n2555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1145_3_lut (.I0(n1603), .I1(n1664[26]), .I2(n1631), 
            .I3(GND_net), .O(n1702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1149_3_lut (.I0(n1607), .I1(n1664[22]), .I2(n1631), 
            .I3(GND_net), .O(n1706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n40451), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n42090), .I0(n2505), .I1(VCC_net), 
            .CO(n42091));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(GND_net), .I1(n2506), .I2(VCC_net), 
            .I3(n42089), .O(n2555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n42089), .I0(n2506), .I1(VCC_net), 
            .CO(n42090));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(GND_net), .I1(n2507), .I2(VCC_net), 
            .I3(n42088), .O(n2555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1152_3_lut (.I0(bit_ctr[19]), .I1(n1664[19]), .I2(n1631), 
            .I3(GND_net), .O(n1709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1144_3_lut (.I0(n1602), .I1(n1664[27]), .I2(n1631), 
            .I3(GND_net), .O(n1701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1569 (.I0(bit_ctr[18]), .I1(n1701), .I2(n1709), 
            .I3(GND_net), .O(n18_adj_5199));
    defparam i5_3_lut_adj_1569.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1741_5 (.CI(n42088), .I0(n2507), .I1(VCC_net), 
            .CO(n42089));
    SB_LUT4 i8_4_lut_adj_1570 (.I0(n1706), .I1(n1702), .I2(n1699), .I3(n1700), 
            .O(n21_adj_5200));
    defparam i8_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1571 (.I0(n1707), .I1(n1698), .I2(n1697), .I3(GND_net), 
            .O(n20_adj_5201));
    defparam i7_3_lut_adj_1571.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(GND_net), .I1(n2508), .I2(VCC_net), 
            .I3(n42087), .O(n2555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut_adj_1572 (.I0(n21_adj_5200), .I1(n1708), .I2(n18_adj_5199), 
            .I3(n1705), .O(n24_adj_5202));
    defparam i11_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1573 (.I0(n1704), .I1(n24_adj_5202), .I2(n20_adj_5201), 
            .I3(n1703), .O(n1730));
    defparam i12_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_679[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n40611), .O(n49879)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_4 (.CI(n42087), .I0(n2508), .I1(VCC_net), 
            .CO(n42088));
    SB_CARRY sub_14_add_2_14 (.CI(n40611), .I0(timer[12]), .I1(n1[12]), 
            .CO(n40612));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(GND_net), .I1(n2509), .I2(GND_net), 
            .I3(n42086), .O(n2555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n42086), .I0(n2509), .I1(GND_net), 
            .CO(n42087));
    SB_CARRY add_21_18 (.CI(n40451), .I0(bit_ctr[16]), .I1(GND_net), .CO(n40452));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(VCC_net), .O(n2555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(GND_net), 
            .CO(n42086));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n40610), .O(one_wire_N_679[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n42085), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n42084), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n42084), .I0(n2589), .I1(n2621), .CO(n42085));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n42083), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n42083), .I0(n2590), .I1(n2621), .CO(n42084));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n42082), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n42082), .I0(n2591), .I1(n2621), .CO(n42083));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n42081), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n42081), .I0(n2592), .I1(n2621), .CO(n42082));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n42080), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n42080), .I0(n2593), .I1(n2621), .CO(n42081));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n42079), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n40450), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_17 (.CI(n40450), .I0(bit_ctr[15]), .I1(GND_net), .CO(n40451));
    SB_CARRY sub_14_add_2_13 (.CI(n40610), .I0(timer[11]), .I1(n1[11]), 
            .CO(n40611));
    SB_LUT4 mod_5_i1079_3_lut (.I0(n1505), .I1(n1565[25]), .I2(n1532), 
            .I3(GND_net), .O(n1604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1083_3_lut (.I0(n1509), .I1(n1565[21]), .I2(n1532), 
            .I3(GND_net), .O(n1608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1808_18 (.CI(n42079), .I0(n2594), .I1(n2621), .CO(n42080));
    SB_LUT4 mod_5_i1082_3_lut (.I0(n1508), .I1(n1565[22]), .I2(n1532), 
            .I3(GND_net), .O(n1607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1077_3_lut (.I0(n1503), .I1(n1565[27]), .I2(n1532), 
            .I3(GND_net), .O(n1602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n42078), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n40449), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n42078), .I0(n2595), .I1(n2621), .CO(n42079));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n42077), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n42077), .I0(n2596), .I1(n2621), .CO(n42078));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n42076), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n42076), .I0(n2597), .I1(n2621), .CO(n42077));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n42075), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n42075), .I0(n2598), .I1(n2621), .CO(n42076));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n42074), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n42074), .I0(n2599), .I1(n2621), .CO(n42075));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n42073), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n42073), .I0(n2600), .I1(n2621), .CO(n42074));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n42072), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n40609), .O(one_wire_N_679[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n42072), .I0(n2601), .I1(n2621), .CO(n42073));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n42071), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n42071), .I0(n2602), .I1(n2621), .CO(n42072));
    SB_CARRY sub_14_add_2_12 (.CI(n40609), .I0(timer[10]), .I1(n1[10]), 
            .CO(n40610));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n42070), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n40449), .I0(bit_ctr[14]), .I1(GND_net), .CO(n40450));
    SB_CARRY mod_5_add_1808_9 (.CI(n42070), .I0(n2603), .I1(n2621), .CO(n42071));
    SB_LUT4 i15_3_lut_4_lut (.I0(state[0]), .I1(n38636), .I2(state[1]), 
            .I3(n38580), .O(n7_adj_5192));
    defparam i15_3_lut_4_lut.LUT_INIT = 16'hefe0;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n42069), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n42069), .I0(n2604), .I1(n2621), .CO(n42070));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n42068), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n42068), .I0(n2605), .I1(n2621), .CO(n42069));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n42067), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n42067), .I0(n2606), .I1(n2621), .CO(n42068));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n42066), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n42066), .I0(n2607), .I1(n2621), .CO(n42067));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n42065), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n42065), .I0(n2608), .I1(n2621), .CO(n42066));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n52730), 
            .I3(n42064), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n42064), .I0(n2609), .I1(n52730), .CO(n42065));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n52730), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n52730), 
            .CO(n42064));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n40448), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2720), .I1(n2687), .I2(VCC_net), 
            .I3(n42063), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(GND_net), .I1(n2688), .I2(VCC_net), 
            .I3(n42062), .O(n2753[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1076_3_lut (.I0(n1502), .I1(n1565[28]), .I2(n1532), 
            .I3(GND_net), .O(n1601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1075_3_lut (.I0(n1501), .I1(n1565[29]), .I2(n1532), 
            .I3(GND_net), .O(n1600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1075_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_15 (.CI(n40448), .I0(bit_ctr[13]), .I1(GND_net), .CO(n40449));
    SB_LUT4 mod_5_i1074_3_lut (.I0(n1500), .I1(n1565[30]), .I2(n1532), 
            .I3(GND_net), .O(n1599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n40608), .O(one_wire_N_679[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_24 (.CI(n42062), .I0(n2688), .I1(VCC_net), 
            .CO(n42063));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(GND_net), .I1(n2689), .I2(VCC_net), 
            .I3(n42061), .O(n2753[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_23 (.CI(n42061), .I0(n2689), .I1(VCC_net), 
            .CO(n42062));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(GND_net), .I1(n2690), .I2(VCC_net), 
            .I3(n42060), .O(n2753[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_22 (.CI(n42060), .I0(n2690), .I1(VCC_net), 
            .CO(n42061));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(GND_net), .I1(n2691), .I2(VCC_net), 
            .I3(n42059), .O(n2753[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_21 (.CI(n42059), .I0(n2691), .I1(VCC_net), 
            .CO(n42060));
    SB_LUT4 mod_5_i1080_3_lut (.I0(n1506), .I1(n1565[24]), .I2(n1532), 
            .I3(GND_net), .O(n1605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(GND_net), .I1(n2692), .I2(VCC_net), 
            .I3(n42058), .O(n2753[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_20 (.CI(n42058), .I0(n2692), .I1(VCC_net), 
            .CO(n42059));
    SB_LUT4 mod_5_i1081_3_lut (.I0(n1507), .I1(n1565[23]), .I2(n1532), 
            .I3(GND_net), .O(n1606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_19_lut (.I0(GND_net), .I1(n2693), .I2(VCC_net), 
            .I3(n42057), .O(n2753[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_19 (.CI(n42057), .I0(n2693), .I1(VCC_net), 
            .CO(n42058));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(GND_net), .I1(n2694), .I2(VCC_net), 
            .I3(n42056), .O(n2753[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_18 (.CI(n42056), .I0(n2694), .I1(VCC_net), 
            .CO(n42057));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(GND_net), .I1(n2695), .I2(VCC_net), 
            .I3(n42055), .O(n2753[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_17 (.CI(n42055), .I0(n2695), .I1(VCC_net), 
            .CO(n42056));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(GND_net), .I1(n2696), .I2(VCC_net), 
            .I3(n42054), .O(n2753[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1013_3_lut (.I0(n1407), .I1(n1466[24]), .I2(n1433), 
            .I3(GND_net), .O(n1506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n40447), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1433), .I1(n1400), .I2(VCC_net), 
            .I3(n41084), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_14 (.CI(n40447), .I0(bit_ctr[12]), .I1(GND_net), .CO(n40448));
    SB_CARRY mod_5_add_1875_16 (.CI(n42054), .I0(n2696), .I1(VCC_net), 
            .CO(n42055));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(GND_net), .I1(n2697), .I2(VCC_net), 
            .I3(n42053), .O(n2753[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n42053), .I0(n2697), .I1(VCC_net), 
            .CO(n42054));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(GND_net), .I1(n2698), .I2(VCC_net), 
            .I3(n42052), .O(n2753[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_14 (.CI(n42052), .I0(n2698), .I1(VCC_net), 
            .CO(n42053));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(GND_net), .I1(n2699), .I2(VCC_net), 
            .I3(n42051), .O(n2753[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_13 (.CI(n42051), .I0(n2699), .I1(VCC_net), 
            .CO(n42052));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(GND_net), .I1(n1401), .I2(VCC_net), 
            .I3(n41083), .O(n1466[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_12_lut (.I0(GND_net), .I1(n2700), .I2(VCC_net), 
            .I3(n42050), .O(n2753[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_12 (.CI(n42050), .I0(n2700), .I1(VCC_net), 
            .CO(n42051));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(GND_net), .I1(n2701), .I2(VCC_net), 
            .I3(n42049), .O(n2753[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n41083), .I0(n1401), .I1(VCC_net), 
            .CO(n41084));
    SB_CARRY mod_5_add_1875_11 (.CI(n42049), .I0(n2701), .I1(VCC_net), 
            .CO(n42050));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(GND_net), .I1(n2702), .I2(VCC_net), 
            .I3(n42048), .O(n2753[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_10 (.CI(n42048), .I0(n2702), .I1(VCC_net), 
            .CO(n42049));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(GND_net), .I1(n2703), .I2(VCC_net), 
            .I3(n42047), .O(n2753[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_10_lut (.I0(GND_net), .I1(n1402), .I2(VCC_net), 
            .I3(n41082), .O(n1466[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_9 (.CI(n42047), .I0(n2703), .I1(VCC_net), 
            .CO(n42048));
    SB_CARRY sub_14_add_2_11 (.CI(n40608), .I0(timer[9]), .I1(n1[9]), 
            .CO(n40609));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(GND_net), .I1(n2704), .I2(VCC_net), 
            .I3(n42046), .O(n2753[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n42046), .I0(n2704), .I1(VCC_net), 
            .CO(n42047));
    SB_CARRY mod_5_add_1004_10 (.CI(n41082), .I0(n1402), .I1(VCC_net), 
            .CO(n41083));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n40607), .O(one_wire_N_679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(GND_net), .I1(n1403), .I2(VCC_net), 
            .I3(n41081), .O(n1466[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_9 (.CI(n41081), .I0(n1403), .I1(VCC_net), 
            .CO(n41082));
    SB_CARRY sub_14_add_2_10 (.CI(n40607), .I0(timer[8]), .I1(n1[8]), 
            .CO(n40608));
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n50217), .I2(n50218), 
            .I3(bit_ctr[2]), .O(n52810));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n52810_bdd_4_lut (.I0(n52810), .I1(n50212), .I2(n50211), .I3(bit_ctr[2]), 
            .O(n52813));
    defparam n52810_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(GND_net), .I1(n2705), .I2(VCC_net), 
            .I3(n42045), .O(n2753[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(GND_net), .I1(n1404), .I2(VCC_net), 
            .I3(n41080), .O(n1466[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_7 (.CI(n42045), .I0(n2705), .I1(VCC_net), 
            .CO(n42046));
    SB_CARRY mod_5_add_1004_8 (.CI(n41080), .I0(n1404), .I1(VCC_net), 
            .CO(n41081));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(GND_net), .I1(n2706), .I2(VCC_net), 
            .I3(n42044), .O(n2753[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_6 (.CI(n42044), .I0(n2706), .I1(VCC_net), 
            .CO(n42045));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(GND_net), .I1(n2707), .I2(VCC_net), 
            .I3(n42043), .O(n2753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_5 (.CI(n42043), .I0(n2707), .I1(VCC_net), 
            .CO(n42044));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(GND_net), .I1(n2708), .I2(VCC_net), 
            .I3(n42042), .O(n2753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n42042), .I0(n2708), .I1(VCC_net), 
            .CO(n42043));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(GND_net), .I1(n2709), .I2(GND_net), 
            .I3(n42041), .O(n2753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n42041), .I0(n2709), .I1(GND_net), 
            .CO(n42042));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(VCC_net), .O(n2753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n40446), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(GND_net), 
            .CO(n42041));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2819), .I1(n2786), .I2(VCC_net), 
            .I3(n42040), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(GND_net), .I1(n1405), .I2(VCC_net), 
            .I3(n41079), .O(n1466[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(GND_net), .I1(n2787), .I2(VCC_net), 
            .I3(n42039), .O(n2852[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n41079), .I0(n1405), .I1(VCC_net), 
            .CO(n41080));
    SB_CARRY mod_5_add_1942_25 (.CI(n42039), .I0(n2787), .I1(VCC_net), 
            .CO(n42040));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(GND_net), .I1(n2788), .I2(VCC_net), 
            .I3(n42038), .O(n2852[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_24 (.CI(n42038), .I0(n2788), .I1(VCC_net), 
            .CO(n42039));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(GND_net), .I1(n2789), .I2(VCC_net), 
            .I3(n42037), .O(n2852[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_6_lut (.I0(GND_net), .I1(n1406), .I2(VCC_net), 
            .I3(n41078), .O(n1466[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_9_lut (.I0(n49871), .I1(timer[7]), .I2(n1[7]), 
            .I3(n40606), .O(n49873)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_13 (.CI(n40446), .I0(bit_ctr[11]), .I1(GND_net), .CO(n40447));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n40445), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_23 (.CI(n42037), .I0(n2789), .I1(VCC_net), 
            .CO(n42038));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(GND_net), .I1(n2790), .I2(VCC_net), 
            .I3(n42036), .O(n2852[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n40606), .I0(timer[7]), .I1(n1[7]), .CO(n40607));
    SB_CARRY mod_5_add_1942_22 (.CI(n42036), .I0(n2790), .I1(VCC_net), 
            .CO(n42037));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(GND_net), .I1(n2791), .I2(VCC_net), 
            .I3(n42035), .O(n2852[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_6 (.CI(n41078), .I0(n1406), .I1(VCC_net), 
            .CO(n41079));
    SB_CARRY mod_5_add_1942_21 (.CI(n42035), .I0(n2791), .I1(VCC_net), 
            .CO(n42036));
    SB_LUT4 mod_5_i1014_3_lut (.I0(n1408), .I1(n1466[23]), .I2(n1433), 
            .I3(GND_net), .O(n1507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(GND_net), .I1(n2792), .I2(VCC_net), 
            .I3(n42034), .O(n2852[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_20 (.CI(n42034), .I0(n2792), .I1(VCC_net), 
            .CO(n42035));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(GND_net), .I1(n2793), .I2(VCC_net), 
            .I3(n42033), .O(n2852[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_19 (.CI(n42033), .I0(n2793), .I1(VCC_net), 
            .CO(n42034));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(GND_net), .I1(n2794), .I2(VCC_net), 
            .I3(n42032), .O(n2852[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_18 (.CI(n42032), .I0(n2794), .I1(VCC_net), 
            .CO(n42033));
    SB_LUT4 mod_5_i1007_3_lut (.I0(n1401), .I1(n1466[30]), .I2(n1433), 
            .I3(GND_net), .O(n1500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1942_17_lut (.I0(GND_net), .I1(n2795), .I2(VCC_net), 
            .I3(n42031), .O(n2852[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_17 (.CI(n42031), .I0(n2795), .I1(VCC_net), 
            .CO(n42032));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(GND_net), .I1(n2796), .I2(VCC_net), 
            .I3(n42030), .O(n2852[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1012_3_lut (.I0(n1406), .I1(n1466[25]), .I2(n1433), 
            .I3(GND_net), .O(n1505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1012_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1942_16 (.CI(n42030), .I0(n2796), .I1(VCC_net), 
            .CO(n42031));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(GND_net), .I1(n2797), .I2(VCC_net), 
            .I3(n42029), .O(n2852[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1016_3_lut (.I0(bit_ctr[21]), .I1(n1466[21]), .I2(n1433), 
            .I3(GND_net), .O(n1509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1942_15 (.CI(n42029), .I0(n2797), .I1(VCC_net), 
            .CO(n42030));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(GND_net), .I1(n2798), .I2(VCC_net), 
            .I3(n42028), .O(n2852[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(GND_net), .I1(n1407), .I2(VCC_net), 
            .I3(n41077), .O(n1466[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_12 (.CI(n40445), .I0(bit_ctr[10]), .I1(GND_net), .CO(n40446));
    SB_LUT4 mod_5_i1010_3_lut (.I0(n1404), .I1(n1466[27]), .I2(n1433), 
            .I3(GND_net), .O(n1503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1010_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1004_5 (.CI(n41077), .I0(n1407), .I1(VCC_net), 
            .CO(n41078));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(GND_net), .I1(n1408), .I2(VCC_net), 
            .I3(n41076), .O(n1466[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_14 (.CI(n42028), .I0(n2798), .I1(VCC_net), 
            .CO(n42029));
    SB_CARRY mod_5_add_1004_4 (.CI(n41076), .I0(n1408), .I1(VCC_net), 
            .CO(n41077));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(GND_net), .I1(n2799), .I2(VCC_net), 
            .I3(n42027), .O(n2852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_3_lut (.I0(GND_net), .I1(n1409), .I2(GND_net), 
            .I3(n41075), .O(n1466[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_13 (.CI(n42027), .I0(n2799), .I1(VCC_net), 
            .CO(n42028));
    SB_LUT4 sub_14_add_2_8_lut (.I0(n49869), .I1(timer[6]), .I2(n1[6]), 
            .I3(n40605), .O(n49871)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(GND_net), .I1(n2800), .I2(VCC_net), 
            .I3(n42026), .O(n2852[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_3 (.CI(n41075), .I0(n1409), .I1(GND_net), 
            .CO(n41076));
    SB_CARRY mod_5_add_1942_12 (.CI(n42026), .I0(n2800), .I1(VCC_net), 
            .CO(n42027));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(GND_net), .I1(n2801), .I2(VCC_net), 
            .I3(n42025), .O(n2852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_11 (.CI(n42025), .I0(n2801), .I1(VCC_net), 
            .CO(n42026));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(GND_net), .I1(n2802), .I2(VCC_net), 
            .I3(n42024), .O(n2852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n40605), .I0(timer[6]), .I1(n1[6]), .CO(n40606));
    SB_LUT4 mod_5_i1011_3_lut (.I0(n1405), .I1(n1466[26]), .I2(n1433), 
            .I3(GND_net), .O(n1504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(VCC_net), .O(n1466[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i946_3_lut (.I0(n1308), .I1(n1367[24]), .I2(n1334), 
            .I3(GND_net), .O(n1407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i944_3_lut (.I0(n1306), .I1(n1367[26]), .I2(n1334), 
            .I3(GND_net), .O(n1405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1942_10 (.CI(n42024), .I0(n2802), .I1(VCC_net), 
            .CO(n42025));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(GND_net), .I1(n2803), .I2(VCC_net), 
            .I3(n42023), .O(n2852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i943_3_lut (.I0(n1305), .I1(n1367[27]), .I2(n1334), 
            .I3(GND_net), .O(n1404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i942_3_lut (.I0(n1304), .I1(n1367[28]), .I2(n1334), 
            .I3(GND_net), .O(n1403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i941_3_lut (.I0(n1303), .I1(n1367[29]), .I2(n1334), 
            .I3(GND_net), .O(n1402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i940_3_lut (.I0(n1302), .I1(n1367[30]), .I2(n1334), 
            .I3(GND_net), .O(n1401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i940_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1942_9 (.CI(n42023), .I0(n2803), .I1(VCC_net), 
            .CO(n42024));
    SB_LUT4 sub_14_add_2_7_lut (.I0(one_wire_N_679[4]), .I1(timer[5]), .I2(n1[5]), 
            .I3(n40604), .O(n49869)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(GND_net), 
            .CO(n41075));
    SB_LUT4 mod_5_i947_3_lut (.I0(n1309), .I1(n1367[23]), .I2(n1334), 
            .I3(GND_net), .O(n1408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(GND_net), .I1(n2804), .I2(VCC_net), 
            .I3(n42022), .O(n2852[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i945_3_lut (.I0(n1307), .I1(n1367[25]), .I2(n1334), 
            .I3(GND_net), .O(n1406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1942_8 (.CI(n42022), .I0(n2804), .I1(VCC_net), 
            .CO(n42023));
    SB_LUT4 i6_4_lut (.I0(n1401), .I1(n1402), .I2(n1400), .I3(n1403), 
            .O(n16_adj_5203));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut_adj_1574 (.I0(n1406), .I1(n16_adj_5203), .I2(n1408), 
            .I3(GND_net), .O(n18_adj_5204));   // verilog/neopixel.v(22[26:36])
    defparam i8_3_lut_adj_1574.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut_adj_1575 (.I0(bit_ctr[21]), .I1(n1404), .I2(n1409), 
            .I3(GND_net), .O(n13_adj_5205));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1575.LUT_INIT = 16'hecec;
    SB_LUT4 i9_4_lut_adj_1576 (.I0(n13_adj_5205), .I1(n18_adj_5204), .I2(n1405), 
            .I3(n1407), .O(n1433));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i948_3_lut (.I0(bit_ctr[22]), .I1(n1367[22]), .I2(n1334), 
            .I3(GND_net), .O(n1409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1015_3_lut (.I0(n1409), .I1(n1466[22]), .I2(n1433), 
            .I3(GND_net), .O(n1508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1009_3_lut (.I0(n1403), .I1(n1466[28]), .I2(n1433), 
            .I3(GND_net), .O(n1502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1008_3_lut (.I0(n1402), .I1(n1466[29]), .I2(n1433), 
            .I3(GND_net), .O(n1501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1008_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_7 (.CI(n40604), .I0(timer[5]), .I1(n1[5]), .CO(n40605));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(GND_net), .I1(n2805), .I2(VCC_net), 
            .I3(n42021), .O(n2852[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_7 (.CI(n42021), .I0(n2805), .I1(VCC_net), 
            .CO(n42022));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(GND_net), .I1(n2806), .I2(VCC_net), 
            .I3(n42020), .O(n2852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n42020), .I0(n2806), .I1(VCC_net), 
            .CO(n42021));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n40444), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(GND_net), .I1(n2807), .I2(VCC_net), 
            .I3(n42019), .O(n2852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_5 (.CI(n42019), .I0(n2807), .I1(VCC_net), 
            .CO(n42020));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(GND_net), .I1(n2808), .I2(VCC_net), 
            .I3(n42018), .O(n2852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_4 (.CI(n42018), .I0(n2808), .I1(VCC_net), 
            .CO(n42019));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(GND_net), .I1(n2809), .I2(GND_net), 
            .I3(n42017), .O(n2852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_3 (.CI(n42017), .I0(n2809), .I1(GND_net), 
            .CO(n42018));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(VCC_net), .O(n2852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(GND_net), 
            .CO(n42017));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2918), .I1(n2885), .I2(VCC_net), 
            .I3(n42016), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(GND_net), .I1(n2886), .I2(VCC_net), 
            .I3(n42015), .O(n2951[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n42015), .I0(n2886), .I1(VCC_net), 
            .CO(n42016));
    SB_LUT4 i22954_2_lut (.I0(bit_ctr[20]), .I1(n1509), .I2(GND_net), 
            .I3(GND_net), .O(n36636));
    defparam i22954_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut (.I0(n1501), .I1(n1502), .I2(n36636), .I3(n1508), 
            .O(n18_adj_5206));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(GND_net), .I1(n2887), .I2(VCC_net), 
            .I3(n42014), .O(n2951[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_2_lut (.I0(n1504), .I1(n1503), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5207));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1577 (.I0(n1505), .I1(n18_adj_5206), .I2(n1500), 
            .I3(n1499), .O(n20_adj_5208));
    defparam i9_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1578 (.I0(n1507), .I1(n20_adj_5208), .I2(n16_adj_5207), 
            .I3(n1506), .O(n1532));
    defparam i10_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1084_3_lut (.I0(bit_ctr[20]), .I1(n1565[20]), .I2(n1532), 
            .I3(GND_net), .O(n1609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1084_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_25 (.CI(n42014), .I0(n2887), .I1(VCC_net), 
            .CO(n42015));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(GND_net), .I1(n2888), .I2(VCC_net), 
            .I3(n42013), .O(n2951[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1078_3_lut (.I0(n1504), .I1(n1565[26]), .I2(n1532), 
            .I3(GND_net), .O(n1603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_3_lut (.I0(n1603), .I1(bit_ctr[19]), .I2(n1609), .I3(GND_net), 
            .O(n16_adj_5209));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_2009_24 (.CI(n42013), .I0(n2888), .I1(VCC_net), 
            .CO(n42014));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n40603), .O(one_wire_N_679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut_adj_1579 (.I0(n1599), .I1(n1600), .I2(n1598), .I3(n1601), 
            .O(n19_adj_5210));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1606), .I1(n1605), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5211));   // verilog/neopixel.v(22[26:36])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(GND_net), .I1(n2889), .I2(VCC_net), 
            .I3(n42012), .O(n2951[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_23 (.CI(n42012), .I0(n2889), .I1(VCC_net), 
            .CO(n42013));
    SB_LUT4 i10_4_lut_adj_1580 (.I0(n19_adj_5210), .I1(n1602), .I2(n16_adj_5209), 
            .I3(n1607), .O(n22_adj_5213));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1581 (.I0(n1608), .I1(n22_adj_5213), .I2(n18_adj_5211), 
            .I3(n1604), .O(n1631));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_22_lut (.I0(GND_net), .I1(n2890), .I2(VCC_net), 
            .I3(n42011), .O(n2951[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n42011), .I0(n2890), .I1(VCC_net), 
            .CO(n42012));
    SB_CARRY sub_14_add_2_6 (.CI(n40603), .I0(timer[4]), .I1(n1[4]), .CO(n40604));
    SB_LUT4 i1_4_lut_adj_1582 (.I0(\neo_pixel_transmitter.done ), .I1(n38574), 
            .I2(n98), .I3(state[0]), .O(n38580));   // verilog/neopixel.v(16[20:25])
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'h0a88;
    SB_LUT4 i19_4_lut_adj_1583 (.I0(bit_ctr[16]), .I1(bit_ctr[25]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[22]), .O(n46));
    defparam i19_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1584 (.I0(bit_ctr[24]), .I1(bit_ctr[26]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i17_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1585 (.I0(bit_ctr[19]), .I1(bit_ctr[23]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[20]), .O(n45));
    defparam i18_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1586 (.I0(bit_ctr[30]), .I1(bit_ctr[21]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[14]), .O(n43));
    defparam i16_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1587 (.I0(bit_ctr[7]), .I1(bit_ctr[17]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[18]), .O(n42));
    defparam i15_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_3_lut_adj_1588 (.I0(bit_ctr[10]), .I1(bit_ctr[12]), .I2(bit_ctr[9]), 
            .I3(GND_net), .O(n41));
    defparam i14_3_lut_adj_1588.LUT_INIT = 16'hfefe;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1589 (.I0(bit_ctr[31]), .I1(bit_ctr[8]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[5]), .O(n47));
    defparam i20_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1590 (.I0(n47), .I1(n52), .I2(n41), .I3(n42), 
            .O(n43659));
    defparam i26_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(bit_ctr[3]), .I1(n42573), .I2(GND_net), 
            .I3(GND_net), .O(n42886));
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_add_2009_21_lut (.I0(GND_net), .I1(n2891), .I2(VCC_net), 
            .I3(n42010), .O(n2951[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_21 (.CI(n42010), .I0(n2891), .I1(VCC_net), 
            .CO(n42011));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n40602), .O(one_wire_N_679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(GND_net), .I1(n2892), .I2(VCC_net), 
            .I3(n42009), .O(n2951[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_20 (.CI(n42009), .I0(n2892), .I1(VCC_net), 
            .CO(n42010));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(GND_net), .I1(n2893), .I2(VCC_net), 
            .I3(n42008), .O(n2951[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n42008), .I0(n2893), .I1(VCC_net), 
            .CO(n42009));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(GND_net), .I1(n2894), .I2(VCC_net), 
            .I3(n42007), .O(n2951[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35561_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(state[1]), .I3(GND_net), .O(n51058));   // verilog/neopixel.v(35[12] 117[6])
    defparam i35561_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i24_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n51058), .I2(state[0]), 
            .I3(n38574), .O(n18_adj_5214));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_4_lut.LUT_INIT = 16'hc5cf;
    SB_CARRY mod_5_add_2009_18 (.CI(n42007), .I0(n2894), .I1(VCC_net), 
            .CO(n42008));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(GND_net), .I1(n2895), .I2(VCC_net), 
            .I3(n42006), .O(n2951[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n40602), .I0(timer[3]), .I1(n1[3]), .CO(n40603));
    SB_CARRY add_21_11 (.CI(n40444), .I0(bit_ctr[9]), .I1(GND_net), .CO(n40445));
    SB_LUT4 i24910_4_lut (.I0(n38580), .I1(n51053), .I2(state[1]), .I3(state[0]), 
            .O(n29590));   // verilog/neopixel.v(16[20:25])
    defparam i24910_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n40601), .O(one_wire_N_679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n40601), .I0(timer[2]), .I1(n1[2]), .CO(n40602));
    SB_CARRY mod_5_add_2009_17 (.CI(n42006), .I0(n2895), .I1(VCC_net), 
            .CO(n42007));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_679[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n40600), .O(n4_adj_5215)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_3 (.CI(n40600), .I0(timer[1]), .I1(n1[1]), .CO(n40601));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(GND_net), .I1(n2896), .I2(VCC_net), 
            .I3(n42005), .O(n2951[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n42005), .I0(n2896), .I1(VCC_net), 
            .CO(n42006));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(GND_net), .I1(n2897), .I2(VCC_net), 
            .I3(n42004), .O(n2951[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n40443), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_15 (.CI(n42004), .I0(n2897), .I1(VCC_net), 
            .CO(n42005));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(GND_net), .I1(n2898), .I2(VCC_net), 
            .I3(n42003), .O(n2951[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_14 (.CI(n42003), .I0(n2898), .I1(VCC_net), 
            .CO(n42004));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(GND_net), .I1(n2899), .I2(VCC_net), 
            .I3(n42002), .O(n2951[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_13 (.CI(n42002), .I0(n2899), .I1(VCC_net), 
            .CO(n42003));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(GND_net), .I1(n2900), .I2(VCC_net), 
            .I3(n42001), .O(n2951[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n42001), .I0(n2900), .I1(VCC_net), 
            .CO(n42002));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(GND_net), .I1(n2901), .I2(VCC_net), 
            .I3(n42000), .O(n2951[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_11 (.CI(n42000), .I0(n2901), .I1(VCC_net), 
            .CO(n42001));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(GND_net), .I1(n2902), .I2(VCC_net), 
            .I3(n41999), .O(n2951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_10 (.CI(n41999), .I0(n2902), .I1(VCC_net), 
            .CO(n42000));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(GND_net), .I1(n2903), .I2(VCC_net), 
            .I3(n41998), .O(n2951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_10 (.CI(n40443), .I0(bit_ctr[8]), .I1(GND_net), .CO(n40444));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n40442), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n40600));
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_9 (.CI(n41998), .I0(n2903), .I1(VCC_net), 
            .CO(n41999));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1532), .I1(n1499), .I2(VCC_net), 
            .I3(n41044), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(GND_net), .I1(n2904), .I2(VCC_net), 
            .I3(n41997), .O(n2951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_8 (.CI(n41997), .I0(n2904), .I1(VCC_net), 
            .CO(n41998));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(GND_net), .I1(n2905), .I2(VCC_net), 
            .I3(n41996), .O(n2951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_7 (.CI(n41996), .I0(n2905), .I1(VCC_net), 
            .CO(n41997));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(GND_net), .I1(n2906), .I2(VCC_net), 
            .I3(n41995), .O(n2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_6 (.CI(n41995), .I0(n2906), .I1(VCC_net), 
            .CO(n41996));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(GND_net), .I1(n2907), .I2(VCC_net), 
            .I3(n41994), .O(n2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(GND_net), .I1(n1500), .I2(VCC_net), 
            .I3(n41043), .O(n1565[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_12 (.CI(n41043), .I0(n1500), .I1(VCC_net), 
            .CO(n41044));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(GND_net), .I1(n1501), .I2(VCC_net), 
            .I3(n41042), .O(n1565[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n41042), .I0(n1501), .I1(VCC_net), 
            .CO(n41043));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(GND_net), .I1(n1502), .I2(VCC_net), 
            .I3(n41041), .O(n1565[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_10 (.CI(n41041), .I0(n1502), .I1(VCC_net), 
            .CO(n41042));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(GND_net), .I1(n1503), .I2(VCC_net), 
            .I3(n41040), .O(n1565[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_9 (.CI(n41040), .I0(n1503), .I1(VCC_net), 
            .CO(n41041));
    SB_CARRY mod_5_add_2009_5 (.CI(n41994), .I0(n2907), .I1(VCC_net), 
            .CO(n41995));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(GND_net), .I1(n1504), .I2(VCC_net), 
            .I3(n41039), .O(n1565[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_8 (.CI(n41039), .I0(n1504), .I1(VCC_net), 
            .CO(n41040));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(GND_net), .I1(n1505), .I2(VCC_net), 
            .I3(n41038), .O(n1565[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_7 (.CI(n41038), .I0(n1505), .I1(VCC_net), 
            .CO(n41039));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(GND_net), .I1(n2908), .I2(VCC_net), 
            .I3(n41993), .O(n2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(GND_net), .I1(n1506), .I2(VCC_net), 
            .I3(n41037), .O(n1565[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_6 (.CI(n41037), .I0(n1506), .I1(VCC_net), 
            .CO(n41038));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(GND_net), .I1(n1507), .I2(VCC_net), 
            .I3(n41036), .O(n1565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_5 (.CI(n41036), .I0(n1507), .I1(VCC_net), 
            .CO(n41037));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(GND_net), .I1(n1508), .I2(VCC_net), 
            .I3(n41035), .O(n1565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_4 (.CI(n41035), .I0(n1508), .I1(VCC_net), 
            .CO(n41036));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(GND_net), .I1(n1509), .I2(GND_net), 
            .I3(n41034), .O(n1565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_3 (.CI(n41034), .I0(n1509), .I1(GND_net), 
            .CO(n41035));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(VCC_net), .O(n1565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(GND_net), 
            .CO(n41034));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n46516), .D(\neo_pixel_transmitter.done_N_742 ), 
            .R(n48388));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_4 (.CI(n41993), .I0(n2908), .I1(VCC_net), 
            .CO(n41994));
    SB_LUT4 i54_3_lut_4_lut (.I0(one_wire_N_679[2]), .I1(n4_adj_5215), .I2(one_wire_N_679[3]), 
            .I3(state[0]), .O(n55));
    defparam i54_3_lut_4_lut.LUT_INIT = 16'hfa88;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(one_wire_N_679[10]), .I1(n121), .I2(GND_net), 
            .I3(GND_net), .O(n45645));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1593 (.I0(one_wire_N_679[10]), .I1(n28470), .I2(one_wire_N_679[8]), 
            .I3(one_wire_N_679[9]), .O(n38635));   // verilog/neopixel.v(6[16:24])
    defparam i1_4_lut_adj_1593.LUT_INIT = 16'heeec;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(\neo_pixel_transmitter.done ), .I1(n38635), 
            .I2(GND_net), .I3(GND_net), .O(n38636));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'h4444;
    SB_LUT4 i30919_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n55), .I3(n45645), .O(n46488));
    defparam i30919_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i35537_2_lut_4_lut (.I0(LED_c), .I1(bit_ctr[4]), .I2(bit_ctr[3]), 
            .I3(n43659), .O(n51053));   // verilog/neopixel.v(16[20:25])
    defparam i35537_2_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 i31_4_lut (.I0(n46488), .I1(n38636), .I2(state[1]), .I3(state[0]), 
            .O(n14));
    defparam i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36601_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_727));   // verilog/neopixel.v(36[4] 116[11])
    defparam i36601_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut_4_lut (.I0(start), .I1(one_wire_N_679[2]), .I2(n4_adj_5215), 
            .I3(n45645), .O(n38574));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h5540;
    SB_LUT4 i1_2_lut_adj_1595 (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/neopixel.v(53[15:25])
    defparam i1_2_lut_adj_1595.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_679[2]), .I1(n4_adj_5215), .I2(GND_net), 
            .I3(GND_net), .O(n75));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(one_wire_N_679[9]), .I1(n28470), .I2(one_wire_N_679[8]), 
            .I3(n49873), .O(n121));   // verilog/neopixel.v(6[16:24])
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(state[1]), .I1(n125), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n8_adj_5216));
    defparam i2_4_lut.LUT_INIT = 16'heaae;
    SB_LUT4 i1_4_lut_adj_1597 (.I0(n121), .I1(n75), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n7_adj_5217));
    defparam i1_4_lut_adj_1597.LUT_INIT = 16'haeea;
    SB_LUT4 i5_4_lut (.I0(start), .I1(n7_adj_5217), .I2(one_wire_N_679[10]), 
            .I3(n8_adj_5216), .O(n52965));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24969_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(16[20:25])
    defparam i24969_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_9 (.CI(n40442), .I0(bit_ctr[7]), .I1(GND_net), .CO(n40443));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n40441), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(GND_net), .I1(n2909), .I2(GND_net), 
            .I3(n41992), .O(n2951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_8 (.CI(n40441), .I0(bit_ctr[6]), .I1(GND_net), .CO(n40442));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n40440), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n41992), .I0(n2909), .I1(GND_net), 
            .CO(n41993));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(VCC_net), .O(n2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(GND_net), 
            .CO(n41992));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n3017), .I1(n2984), .I2(VCC_net), 
            .I3(n41991), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(GND_net), .I1(n2985), .I2(VCC_net), 
            .I3(n41990), .O(n3050[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_27 (.CI(n41990), .I0(n2985), .I1(VCC_net), 
            .CO(n41991));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(GND_net), .I1(n2986), .I2(VCC_net), 
            .I3(n41989), .O(n3050[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_26 (.CI(n41989), .I0(n2986), .I1(VCC_net), 
            .CO(n41990));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(GND_net), .I1(n2987), .I2(VCC_net), 
            .I3(n41988), .O(n3050[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_25 (.CI(n41988), .I0(n2987), .I1(VCC_net), 
            .CO(n41989));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(GND_net), .I1(n2988), .I2(VCC_net), 
            .I3(n41987), .O(n3050[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_24 (.CI(n41987), .I0(n2988), .I1(VCC_net), 
            .CO(n41988));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(GND_net), .I1(n2989), .I2(VCC_net), 
            .I3(n41986), .O(n3050[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_23 (.CI(n41986), .I0(n2989), .I1(VCC_net), 
            .CO(n41987));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(GND_net), .I1(n2990), .I2(VCC_net), 
            .I3(n41985), .O(n3050[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_22 (.CI(n41985), .I0(n2990), .I1(VCC_net), 
            .CO(n41986));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(GND_net), .I1(n2991), .I2(VCC_net), 
            .I3(n41984), .O(n3050[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_21 (.CI(n41984), .I0(n2991), .I1(VCC_net), 
            .CO(n41985));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(GND_net), .I1(n2992), .I2(VCC_net), 
            .I3(n41983), .O(n3050[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_20 (.CI(n41983), .I0(n2992), .I1(VCC_net), 
            .CO(n41984));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(GND_net), .I1(n2993), .I2(VCC_net), 
            .I3(n41982), .O(n3050[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_19 (.CI(n41982), .I0(n2993), .I1(VCC_net), 
            .CO(n41983));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(GND_net), .I1(n2994), .I2(VCC_net), 
            .I3(n41981), .O(n3050[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_18 (.CI(n41981), .I0(n2994), .I1(VCC_net), 
            .CO(n41982));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(GND_net), .I1(n2995), .I2(VCC_net), 
            .I3(n41980), .O(n3050[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_17 (.CI(n41980), .I0(n2995), .I1(VCC_net), 
            .CO(n41981));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(GND_net), .I1(n2996), .I2(VCC_net), 
            .I3(n41979), .O(n3050[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_16 (.CI(n41979), .I0(n2996), .I1(VCC_net), 
            .CO(n41980));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(GND_net), .I1(n2997), .I2(VCC_net), 
            .I3(n41978), .O(n3050[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_15 (.CI(n41978), .I0(n2997), .I1(VCC_net), 
            .CO(n41979));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(GND_net), .I1(n2998), .I2(VCC_net), 
            .I3(n41977), .O(n3050[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_14 (.CI(n41977), .I0(n2998), .I1(VCC_net), 
            .CO(n41978));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(GND_net), .I1(n2999), .I2(VCC_net), 
            .I3(n41976), .O(n3050[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_13 (.CI(n41976), .I0(n2999), .I1(VCC_net), 
            .CO(n41977));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(GND_net), .I1(n3000), .I2(VCC_net), 
            .I3(n41975), .O(n3050[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_12 (.CI(n41975), .I0(n3000), .I1(VCC_net), 
            .CO(n41976));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(GND_net), .I1(n3001), .I2(VCC_net), 
            .I3(n41974), .O(n3050[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_11 (.CI(n41974), .I0(n3001), .I1(VCC_net), 
            .CO(n41975));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(GND_net), .I1(n3002), .I2(VCC_net), 
            .I3(n41973), .O(n3050[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_10 (.CI(n41973), .I0(n3002), .I1(VCC_net), 
            .CO(n41974));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(GND_net), .I1(n3003), .I2(VCC_net), 
            .I3(n41972), .O(n3050[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_9 (.CI(n41972), .I0(n3003), .I1(VCC_net), 
            .CO(n41973));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(GND_net), .I1(n3004), .I2(VCC_net), 
            .I3(n41971), .O(n3050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_8 (.CI(n41971), .I0(n3004), .I1(VCC_net), 
            .CO(n41972));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(GND_net), .I1(n3005), .I2(VCC_net), 
            .I3(n41970), .O(n3050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_7 (.CI(n41970), .I0(n3005), .I1(VCC_net), 
            .CO(n41971));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(GND_net), .I1(n3006), .I2(VCC_net), 
            .I3(n41969), .O(n3050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_6 (.CI(n41969), .I0(n3006), .I1(VCC_net), 
            .CO(n41970));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(GND_net), .I1(n3007), .I2(VCC_net), 
            .I3(n41968), .O(n3050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_5 (.CI(n41968), .I0(n3007), .I1(VCC_net), 
            .CO(n41969));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(GND_net), .I1(n3008), .I2(VCC_net), 
            .I3(n41967), .O(n3050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_4 (.CI(n41967), .I0(n3008), .I1(VCC_net), 
            .CO(n41968));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(GND_net), .I1(n3009), .I2(GND_net), 
            .I3(n41966), .O(n3050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_3 (.CI(n41966), .I0(n3009), .I1(GND_net), 
            .CO(n41967));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(VCC_net), .O(n3050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(GND_net), 
            .CO(n41966));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3116), .I1(n3083), .I2(VCC_net), 
            .I3(n41965), .O(n50010)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(GND_net), .I1(n3084), .I2(VCC_net), 
            .I3(n41964), .O(n3149[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_28 (.CI(n41964), .I0(n3084), .I1(VCC_net), 
            .CO(n41965));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(GND_net), .I1(n3085), .I2(VCC_net), 
            .I3(n41963), .O(n3149[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n41963), .I0(n3085), .I1(VCC_net), 
            .CO(n41964));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(GND_net), .I1(n3086), .I2(VCC_net), 
            .I3(n41962), .O(n3149[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_26 (.CI(n41962), .I0(n3086), .I1(VCC_net), 
            .CO(n41963));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(GND_net), .I1(n3087), .I2(VCC_net), 
            .I3(n41961), .O(n3149[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_25 (.CI(n41961), .I0(n3087), .I1(VCC_net), 
            .CO(n41962));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(GND_net), .I1(n3088), .I2(VCC_net), 
            .I3(n41960), .O(n3149[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_24 (.CI(n41960), .I0(n3088), .I1(VCC_net), 
            .CO(n41961));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(GND_net), .I1(n3089), .I2(VCC_net), 
            .I3(n41959), .O(n3149[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_23 (.CI(n41959), .I0(n3089), .I1(VCC_net), 
            .CO(n41960));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(GND_net), .I1(n3090), .I2(VCC_net), 
            .I3(n41958), .O(n3149[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n41958), .I0(n3090), .I1(VCC_net), 
            .CO(n41959));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(GND_net), .I1(n3091), .I2(VCC_net), 
            .I3(n41957), .O(n3149[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_21 (.CI(n41957), .I0(n3091), .I1(VCC_net), 
            .CO(n41958));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(GND_net), .I1(n3092), .I2(VCC_net), 
            .I3(n41956), .O(n3149[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_20 (.CI(n41956), .I0(n3092), .I1(VCC_net), 
            .CO(n41957));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(GND_net), .I1(n3093), .I2(VCC_net), 
            .I3(n41955), .O(n3149[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_19 (.CI(n41955), .I0(n3093), .I1(VCC_net), 
            .CO(n41956));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(GND_net), .I1(n3094), .I2(VCC_net), 
            .I3(n41954), .O(n3149[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_18 (.CI(n41954), .I0(n3094), .I1(VCC_net), 
            .CO(n41955));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(GND_net), .I1(n3095), .I2(VCC_net), 
            .I3(n41953), .O(n3149[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_17 (.CI(n41953), .I0(n3095), .I1(VCC_net), 
            .CO(n41954));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(GND_net), .I1(n3096), .I2(VCC_net), 
            .I3(n41952), .O(n3149[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_16 (.CI(n41952), .I0(n3096), .I1(VCC_net), 
            .CO(n41953));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(GND_net), .I1(n3097), .I2(VCC_net), 
            .I3(n41951), .O(n3149[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_15 (.CI(n41951), .I0(n3097), .I1(VCC_net), 
            .CO(n41952));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(GND_net), .I1(n3098), .I2(VCC_net), 
            .I3(n41950), .O(n3149[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_14 (.CI(n41950), .I0(n3098), .I1(VCC_net), 
            .CO(n41951));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(GND_net), .I1(n3099), .I2(VCC_net), 
            .I3(n41949), .O(n3149[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n41949), .I0(n3099), .I1(VCC_net), 
            .CO(n41950));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(GND_net), .I1(n3100), .I2(VCC_net), 
            .I3(n41948), .O(n3149[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_12 (.CI(n41948), .I0(n3100), .I1(VCC_net), 
            .CO(n41949));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(GND_net), .I1(n3101), .I2(VCC_net), 
            .I3(n41947), .O(n3149[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_11 (.CI(n41947), .I0(n3101), .I1(VCC_net), 
            .CO(n41948));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(GND_net), .I1(n3102), .I2(VCC_net), 
            .I3(n41946), .O(n3149[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_10 (.CI(n41946), .I0(n3102), .I1(VCC_net), 
            .CO(n41947));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(GND_net), .I1(n3103), .I2(VCC_net), 
            .I3(n41945), .O(n3149[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_9 (.CI(n41945), .I0(n3103), .I1(VCC_net), 
            .CO(n41946));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(GND_net), .I1(n3104), .I2(VCC_net), 
            .I3(n41944), .O(n3149[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_8 (.CI(n41944), .I0(n3104), .I1(VCC_net), 
            .CO(n41945));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(GND_net), .I1(n3105), .I2(VCC_net), 
            .I3(n41943), .O(n3149[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_7 (.CI(n41943), .I0(n3105), .I1(VCC_net), 
            .CO(n41944));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(GND_net), .I1(n3106), .I2(VCC_net), 
            .I3(n41942), .O(n3149[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_6 (.CI(n41942), .I0(n3106), .I1(VCC_net), 
            .CO(n41943));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(GND_net), .I1(n3107), .I2(VCC_net), 
            .I3(n41941), .O(n3149[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_5 (.CI(n41941), .I0(n3107), .I1(VCC_net), 
            .CO(n41942));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(GND_net), .I1(n3108), .I2(VCC_net), 
            .I3(n41940), .O(n3149[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_4 (.CI(n41940), .I0(n3108), .I1(VCC_net), 
            .CO(n41941));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(GND_net), .I1(n3109), .I2(GND_net), 
            .I3(n41939), .O(n3149[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_3 (.CI(n41939), .I0(n3109), .I1(GND_net), 
            .CO(n41940));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(VCC_net), .O(n3149[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(GND_net), 
            .CO(n41939));
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n50261), .I2(n50267), 
            .I3(n42886), .O(n52768));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF timer_2188__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2188__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i1_3_lut_4_lut_adj_1598 (.I0(n29881), .I1(bit_ctr[26]), .I2(bit_ctr[27]), 
            .I3(n838), .O(n49527));
    defparam i1_3_lut_4_lut_adj_1598.LUT_INIT = 16'h1551;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n30122));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_7 (.CI(n40440), .I0(bit_ctr[5]), .I1(GND_net), .CO(n40441));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n40439), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23109_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[31]), .I2(bit_ctr[30]), 
            .I3(GND_net), .O(n36796));
    defparam i23109_2_lut_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i5702_2_lut_3_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(GND_net), .O(n12165));   // verilog/neopixel.v(22[26:36])
    defparam i5702_2_lut_3_lut.LUT_INIT = 16'h9090;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n46352), .I1(n26854), .I2(bit_ctr[27]), 
            .I3(n838), .O(n46442));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'haa65;
    SB_CARRY add_21_6 (.CI(n40439), .I0(bit_ctr[4]), .I1(GND_net), .CO(n40440));
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n40438), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n52768_bdd_4_lut (.I0(n52768), .I1(n52735), .I2(n50183), .I3(n42886), 
            .O(n52771));
    defparam n52768_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_21_5 (.CI(n40438), .I0(bit_ctr[3]), .I1(GND_net), .CO(n40439));
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n40437), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n40437), .I0(bit_ctr[2]), .I1(GND_net), .CO(n40438));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n40436), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2188_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n41769), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2188_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n41768), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_32 (.CI(n41768), .I0(GND_net), .I1(timer[30]), 
            .CO(n41769));
    SB_LUT4 timer_2188_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n41767), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_31 (.CI(n41767), .I0(GND_net), .I1(timer[29]), 
            .CO(n41768));
    SB_LUT4 timer_2188_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n41766), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_30 (.CI(n41766), .I0(GND_net), .I1(timer[28]), 
            .CO(n41767));
    SB_LUT4 timer_2188_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n41765), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_29 (.CI(n41765), .I0(GND_net), .I1(timer[27]), 
            .CO(n41766));
    SB_LUT4 timer_2188_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n41764), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_28 (.CI(n41764), .I0(GND_net), .I1(timer[26]), 
            .CO(n41765));
    SB_LUT4 timer_2188_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n41763), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n40436), .I0(bit_ctr[1]), .I1(GND_net), .CO(n40437));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_27 (.CI(n41763), .I0(GND_net), .I1(timer[25]), 
            .CO(n41764));
    SB_LUT4 timer_2188_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n41762), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_26 (.CI(n41762), .I0(GND_net), .I1(timer[24]), 
            .CO(n41763));
    SB_LUT4 mod_5_i2087_3_lut (.I0(n2993), .I1(n3050[22]), .I2(n3017), 
            .I3(GND_net), .O(n3092));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2087_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n40436));
    SB_LUT4 timer_2188_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n41761), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_25 (.CI(n41761), .I0(GND_net), .I1(timer[23]), 
            .CO(n41762));
    SB_LUT4 mod_5_i2100_3_lut (.I0(n3006), .I1(n3050[9]), .I2(n3017), 
            .I3(GND_net), .O(n3105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n41760), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i2093_3_lut (.I0(n2999), .I1(n3050[16]), .I2(n3017), 
            .I3(GND_net), .O(n3098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2097_3_lut (.I0(n3003), .I1(n3050[12]), .I2(n3017), 
            .I3(GND_net), .O(n3102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2096_3_lut (.I0(n3002), .I1(n3050[13]), .I2(n3017), 
            .I3(GND_net), .O(n3101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2102_3_lut (.I0(n3008), .I1(n3050[7]), .I2(n3017), 
            .I3(GND_net), .O(n3107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2092_3_lut (.I0(n2998), .I1(n3050[17]), .I2(n3017), 
            .I3(GND_net), .O(n3097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2090_3_lut (.I0(n2996), .I1(n3050[19]), .I2(n3017), 
            .I3(GND_net), .O(n3095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2090_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_24 (.CI(n41760), .I0(GND_net), .I1(timer[22]), 
            .CO(n41761));
    SB_LUT4 timer_2188_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n41759), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2188_add_4_23 (.CI(n41759), .I0(GND_net), .I1(timer[21]), 
            .CO(n41760));
    SB_LUT4 timer_2188_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n41758), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i2079_3_lut (.I0(n2985), .I1(n3050[30]), .I2(n3017), 
            .I3(GND_net), .O(n3084));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_22 (.CI(n41758), .I0(GND_net), .I1(timer[20]), 
            .CO(n41759));
    SB_LUT4 mod_5_i2103_3_lut (.I0(n3009), .I1(n3050[6]), .I2(n3017), 
            .I3(GND_net), .O(n3108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2104_3_lut (.I0(bit_ctr[5]), .I1(n3050[5]), .I2(n3017), 
            .I3(GND_net), .O(n3109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2188_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n41757), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2188_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i2094_3_lut (.I0(n3000), .I1(n3050[15]), .I2(n3017), 
            .I3(GND_net), .O(n3099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2099_3_lut (.I0(n3005), .I1(n3050[10]), .I2(n3017), 
            .I3(GND_net), .O(n3104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2085_3_lut (.I0(n2991), .I1(n3050[24]), .I2(n3017), 
            .I3(GND_net), .O(n3090));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2086_3_lut (.I0(n2992), .I1(n3050[23]), .I2(n3017), 
            .I3(GND_net), .O(n3091));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2084_3_lut (.I0(n2990), .I1(n3050[25]), .I2(n3017), 
            .I3(GND_net), .O(n3089));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2083_3_lut (.I0(n2989), .I1(n3050[26]), .I2(n3017), 
            .I3(GND_net), .O(n3088));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2188_add_4_21 (.CI(n41757), .I0(GND_net), .I1(timer[19]), 
            .CO(n41758));
    SB_LUT4 mod_5_i2081_3_lut (.I0(n2987), .I1(n3050[28]), .I2(n3017), 
            .I3(GND_net), .O(n3086));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2082_3_lut (.I0(n2988), .I1(n3050[27]), .I2(n3017), 
            .I3(GND_net), .O(n3087));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2080_3_lut (.I0(n2986), .I1(n3050[29]), .I2(n3017), 
            .I3(GND_net), .O(n3085));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2098_3_lut (.I0(n3004), .I1(n3050[11]), .I2(n3017), 
            .I3(GND_net), .O(n3103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2089_3_lut (.I0(n2995), .I1(n3050[20]), .I2(n3017), 
            .I3(GND_net), .O(n3094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2033_3_lut (.I0(n2907), .I1(n2951[9]), .I2(n2918), 
            .I3(GND_net), .O(n3006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2034_3_lut (.I0(n2908), .I1(n2951[8]), .I2(n2918), 
            .I3(GND_net), .O(n3007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2023_3_lut (.I0(n2897), .I1(n2951[19]), .I2(n2918), 
            .I3(GND_net), .O(n2996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2018_3_lut (.I0(n2892), .I1(n2951[24]), .I2(n2918), 
            .I3(GND_net), .O(n2991));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2016_3_lut (.I0(n2890), .I1(n2951[26]), .I2(n2918), 
            .I3(GND_net), .O(n2989));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2017_3_lut (.I0(n2891), .I1(n2951[25]), .I2(n2918), 
            .I3(GND_net), .O(n2990));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2015_3_lut (.I0(n2889), .I1(n2951[27]), .I2(n2918), 
            .I3(GND_net), .O(n2988));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2022_3_lut (.I0(n2896), .I1(n2951[20]), .I2(n2918), 
            .I3(GND_net), .O(n2995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2020_3_lut (.I0(n2894), .I1(n2951[22]), .I2(n2918), 
            .I3(GND_net), .O(n2993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2021_3_lut (.I0(n2895), .I1(n2951[21]), .I2(n2918), 
            .I3(GND_net), .O(n2994));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2019_3_lut (.I0(n2893), .I1(n2951[23]), .I2(n2918), 
            .I3(GND_net), .O(n2992));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2014_3_lut (.I0(n2888), .I1(n2951[28]), .I2(n2918), 
            .I3(GND_net), .O(n2987));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2013_3_lut (.I0(n2887), .I1(n2951[29]), .I2(n2918), 
            .I3(GND_net), .O(n2986));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2012_3_lut (.I0(n2886), .I1(n2951[30]), .I2(n2918), 
            .I3(GND_net), .O(n2985));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2032_3_lut (.I0(n2906), .I1(n2951[10]), .I2(n2918), 
            .I3(GND_net), .O(n3005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2031_3_lut (.I0(n2905), .I1(n2951[11]), .I2(n2918), 
            .I3(GND_net), .O(n3004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2027_3_lut (.I0(n2901), .I1(n2951[15]), .I2(n2918), 
            .I3(GND_net), .O(n3000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2029_3_lut (.I0(n2903), .I1(n2951[13]), .I2(n2918), 
            .I3(GND_net), .O(n3002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2028_3_lut (.I0(n2902), .I1(n2951[14]), .I2(n2918), 
            .I3(GND_net), .O(n3001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2035_3_lut (.I0(n2909), .I1(n2951[7]), .I2(n2918), 
            .I3(GND_net), .O(n3008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2026_3_lut (.I0(n2900), .I1(n2951[16]), .I2(n2918), 
            .I3(GND_net), .O(n2999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2030_3_lut (.I0(n2904), .I1(n2951[12]), .I2(n2918), 
            .I3(GND_net), .O(n3003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1953_3_lut (.I0(n2795), .I1(n2852[22]), .I2(n2819), 
            .I3(GND_net), .O(n2894));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1961_3_lut (.I0(n2803), .I1(n2852[14]), .I2(n2819), 
            .I3(GND_net), .O(n2902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1951_3_lut (.I0(n2793), .I1(n2852[24]), .I2(n2819), 
            .I3(GND_net), .O(n2892));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1950_3_lut (.I0(n2792), .I1(n2852[25]), .I2(n2819), 
            .I3(GND_net), .O(n2891));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1967_3_lut (.I0(n2809), .I1(n2852[8]), .I2(n2819), 
            .I3(GND_net), .O(n2908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1965_3_lut (.I0(n2807), .I1(n2852[10]), .I2(n2819), 
            .I3(GND_net), .O(n2906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1956_3_lut (.I0(n2798), .I1(n2852[19]), .I2(n2819), 
            .I3(GND_net), .O(n2897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1952_3_lut (.I0(n2794), .I1(n2852[23]), .I2(n2819), 
            .I3(GND_net), .O(n2893));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1960_3_lut (.I0(n2802), .I1(n2852[15]), .I2(n2819), 
            .I3(GND_net), .O(n2901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1954_3_lut (.I0(n2796), .I1(n2852[21]), .I2(n2819), 
            .I3(GND_net), .O(n2895));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1962_3_lut (.I0(n2804), .I1(n2852[13]), .I2(n2819), 
            .I3(GND_net), .O(n2903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1966_3_lut (.I0(n2808), .I1(n2852[9]), .I2(n2819), 
            .I3(GND_net), .O(n2907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1949_3_lut (.I0(n2791), .I1(n2852[26]), .I2(n2819), 
            .I3(GND_net), .O(n2890));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1947_3_lut (.I0(n2789), .I1(n2852[28]), .I2(n2819), 
            .I3(GND_net), .O(n2888));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1948_3_lut (.I0(n2790), .I1(n2852[27]), .I2(n2819), 
            .I3(GND_net), .O(n2889));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1946_3_lut (.I0(n2788), .I1(n2852[29]), .I2(n2819), 
            .I3(GND_net), .O(n2887));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1957_3_lut (.I0(n2799), .I1(n2852[18]), .I2(n2819), 
            .I3(GND_net), .O(n2898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(n125), .I1(n45645), .I2(start), .I3(GND_net), 
            .O(n98));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf1f1;
    SB_LUT4 mod_5_i1955_3_lut (.I0(n2797), .I1(n2852[20]), .I2(n2819), 
            .I3(GND_net), .O(n2896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1963_3_lut (.I0(n2805), .I1(n2852[12]), .I2(n2819), 
            .I3(GND_net), .O(n2904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1964_3_lut (.I0(n2806), .I1(n2852[11]), .I2(n2819), 
            .I3(GND_net), .O(n2905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1896_3_lut (.I0(n2706), .I1(n2753[12]), .I2(n2720), 
            .I3(GND_net), .O(n2805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1892_3_lut (.I0(n2702), .I1(n2753[16]), .I2(n2720), 
            .I3(GND_net), .O(n2801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1895_3_lut (.I0(n2705), .I1(n2753[13]), .I2(n2720), 
            .I3(GND_net), .O(n2804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1891_3_lut (.I0(n2701), .I1(n2753[17]), .I2(n2720), 
            .I3(GND_net), .O(n2800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1890_3_lut (.I0(n2700), .I1(n2753[18]), .I2(n2720), 
            .I3(GND_net), .O(n2799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1599 (.I0(n125), .I1(n45645), .I2(n18_adj_5214), 
            .I3(n29590), .O(n30005));
    defparam i1_3_lut_4_lut_adj_1599.LUT_INIT = 16'hf100;
    SB_LUT4 mod_5_i1889_3_lut (.I0(n2699), .I1(n2753[19]), .I2(n2720), 
            .I3(GND_net), .O(n2798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1884_3_lut (.I0(n2694), .I1(n2753[24]), .I2(n2720), 
            .I3(GND_net), .O(n2793));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1882_3_lut (.I0(n2692), .I1(n2753[26]), .I2(n2720), 
            .I3(GND_net), .O(n2791));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1883_3_lut (.I0(n2693), .I1(n2753[25]), .I2(n2720), 
            .I3(GND_net), .O(n2792));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1881_3_lut (.I0(n2691), .I1(n2753[27]), .I2(n2720), 
            .I3(GND_net), .O(n2790));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1899_3_lut (.I0(n2709), .I1(n2753[9]), .I2(n2720), 
            .I3(GND_net), .O(n2808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1898_3_lut (.I0(n2708), .I1(n2753[10]), .I2(n2720), 
            .I3(GND_net), .O(n2807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35522_3_lut_4_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(state[0]), 
            .I3(n43659), .O(n51038));
    defparam i35522_3_lut_4_lut.LUT_INIT = 16'h0070;
    SB_LUT4 mod_5_i1897_3_lut (.I0(n2707), .I1(n2753[11]), .I2(n2720), 
            .I3(GND_net), .O(n2806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1894_3_lut (.I0(n2704), .I1(n2753[14]), .I2(n2720), 
            .I3(GND_net), .O(n2803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1600 (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n43659), 
            .I3(GND_net), .O(n128));
    defparam i1_2_lut_3_lut_adj_1600.LUT_INIT = 16'hf8f8;
    SB_LUT4 mod_5_i1880_3_lut (.I0(n2690), .I1(n2753[28]), .I2(n2720), 
            .I3(GND_net), .O(n2789));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1879_3_lut (.I0(n2689), .I1(n2753[29]), .I2(n2720), 
            .I3(GND_net), .O(n2788));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1601 (.I0(n2703), .I1(bit_ctr[8]), .I2(n2709), 
            .I3(GND_net), .O(n28_adj_5218));
    defparam i5_3_lut_adj_1601.LUT_INIT = 16'heaea;
    SB_LUT4 i15_4_lut_adj_1602 (.I0(n2702), .I1(n2700), .I2(n2695), .I3(n2705), 
            .O(n38_adj_5219));
    defparam i15_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1603 (.I0(n2689), .I1(n2691), .I2(n2690), .I3(n2692), 
            .O(n36_adj_5220));
    defparam i13_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1604 (.I0(n2693), .I1(n38_adj_5219), .I2(n28_adj_5218), 
            .I3(n2697), .O(n42_adj_5221));
    defparam i19_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1605 (.I0(n2708), .I1(n2698), .I2(n2706), .I3(n2707), 
            .O(n40_adj_5222));
    defparam i17_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1606 (.I0(n2704), .I1(n36_adj_5220), .I2(n2688), 
            .I3(n2687), .O(n41_adj_5223));
    defparam i18_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1607 (.I0(n2696), .I1(n2694), .I2(n2701), .I3(n2699), 
            .O(n39_adj_5224));
    defparam i16_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_5224), .I1(n41_adj_5223), .I2(n40_adj_5222), 
            .I3(n42_adj_5221), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1888_3_lut (.I0(n2698), .I1(n2753[20]), .I2(n2720), 
            .I3(GND_net), .O(n2797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1886_3_lut (.I0(n2696), .I1(n2753[22]), .I2(n2720), 
            .I3(GND_net), .O(n2795));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1887_3_lut (.I0(n2697), .I1(n2753[21]), .I2(n2720), 
            .I3(GND_net), .O(n2796));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1885_3_lut (.I0(n2695), .I1(n2753[23]), .I2(n2720), 
            .I3(GND_net), .O(n2794));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1900_3_lut (.I0(bit_ctr[8]), .I1(n2753[8]), .I2(n2720), 
            .I3(GND_net), .O(n2809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1893_3_lut (.I0(n2703), .I1(n2753[15]), .I2(n2720), 
            .I3(GND_net), .O(n2802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_3_lut_adj_1608 (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), 
            .I3(GND_net), .O(n32_adj_5225));   // verilog/neopixel.v(22[26:36])
    defparam i8_3_lut_adj_1608.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1609 (.I0(n2794), .I1(n2796), .I2(n2795), .I3(n2797), 
            .O(n39_adj_5226));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1610 (.I0(n2788), .I1(n2789), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_5227));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut_adj_1610.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1611 (.I0(n2790), .I1(n2792), .I2(n2791), .I3(n2793), 
            .O(n38_adj_5228));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1612 (.I0(n39_adj_5226), .I1(n2798), .I2(n32_adj_5225), 
            .I3(n2799), .O(n44_adj_5229));   // verilog/neopixel.v(22[26:36])
    defparam i20_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1613 (.I0(n2800), .I1(n2804), .I2(n2801), .I3(n2805), 
            .O(n42_adj_5230));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1614 (.I0(n2787), .I1(n38_adj_5228), .I2(n26_adj_5227), 
            .I3(n2786), .O(n43_adj_5231));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1615 (.I0(n2803), .I1(n2806), .I2(n2807), .I3(n2808), 
            .O(n41_adj_5232));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_5232), .I1(n43_adj_5231), .I2(n42_adj_5230), 
            .I3(n44_adj_5229), .O(n2819));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1878_3_lut (.I0(n2688), .I1(n2753[30]), .I2(n2720), 
            .I3(GND_net), .O(n2787));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1945_3_lut (.I0(n2787), .I1(n2852[30]), .I2(n2819), 
            .I3(GND_net), .O(n2886));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1958_3_lut (.I0(n2800), .I1(n2852[17]), .I2(n2819), 
            .I3(GND_net), .O(n2899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1968_3_lut (.I0(bit_ctr[7]), .I1(n2852[7]), .I2(n2819), 
            .I3(GND_net), .O(n2909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1959_3_lut (.I0(n2801), .I1(n2852[16]), .I2(n2819), 
            .I3(GND_net), .O(n2900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1616 (.I0(n2900), .I1(bit_ctr[6]), .I2(n2909), 
            .I3(GND_net), .O(n30_adj_5233));
    defparam i5_3_lut_adj_1616.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1617 (.I0(n2887), .I1(n2889), .I2(n2888), .I3(n2890), 
            .O(n39_adj_5234));
    defparam i14_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2899), .I1(n2886), .I2(n2885), .I3(GND_net), 
            .O(n38_adj_5235));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1618 (.I0(n2905), .I1(n2904), .I2(n2896), .I3(n2898), 
            .O(n43_adj_5236));
    defparam i18_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1619 (.I0(n2907), .I1(n2903), .I2(n2895), .I3(n2901), 
            .O(n42_adj_5237));
    defparam i17_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1620 (.I0(n2893), .I1(n2897), .I2(n2906), .I3(n2908), 
            .O(n41_adj_5238));
    defparam i16_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1621 (.I0(n39_adj_5234), .I1(n2891), .I2(n30_adj_5233), 
            .I3(n2892), .O(n45_adj_5239));
    defparam i20_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1622 (.I0(n43_adj_5236), .I1(n2902), .I2(n38_adj_5235), 
            .I3(n2894), .O(n47_adj_5240));
    defparam i22_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1623 (.I0(n47_adj_5240), .I1(n45_adj_5239), .I2(n41_adj_5238), 
            .I3(n42_adj_5237), .O(n2918));
    defparam i24_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2036_3_lut (.I0(bit_ctr[6]), .I1(n2951[6]), .I2(n2918), 
            .I3(GND_net), .O(n3009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2025_3_lut (.I0(n2899), .I1(n2951[17]), .I2(n2918), 
            .I3(GND_net), .O(n2998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_3_lut_adj_1624 (.I0(n2998), .I1(bit_ctr[5]), .I2(n3009), 
            .I3(GND_net), .O(n34_adj_5241));   // verilog/neopixel.v(22[26:36])
    defparam i8_3_lut_adj_1624.LUT_INIT = 16'heaea;
    SB_LUT4 i18_4_lut_adj_1625 (.I0(n3003), .I1(n2999), .I2(n3008), .I3(n3001), 
            .O(n44_adj_5242));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1626 (.I0(n2985), .I1(n2986), .I2(n2984), .I3(n2987), 
            .O(n40_adj_5243));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1627 (.I0(n3002), .I1(n3000), .I2(n3004), .I3(n3005), 
            .O(n45_adj_5244));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1628 (.I0(n2992), .I1(n2994), .I2(n2993), .I3(n2995), 
            .O(n42_adj_5245));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1629 (.I0(n2996), .I1(n44_adj_5242), .I2(n34_adj_5241), 
            .I3(n2997), .O(n48));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1630 (.I0(n2988), .I1(n2990), .I2(n2989), .I3(n2991), 
            .O(n41_adj_5246));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1631 (.I0(n45_adj_5244), .I1(n3007), .I2(n40_adj_5243), 
            .I3(n3006), .O(n49));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1632 (.I0(n49), .I1(n41_adj_5246), .I2(n48), 
            .I3(n42_adj_5245), .O(n3017));   // verilog/neopixel.v(22[26:36])
    defparam i25_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2024_3_lut (.I0(n2898), .I1(n2951[18]), .I2(n2918), 
            .I3(GND_net), .O(n2997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2088_3_lut (.I0(n2994), .I1(n3050[21]), .I2(n3017), 
            .I3(GND_net), .O(n3093));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2091_3_lut (.I0(n2997), .I1(n3050[18]), .I2(n3017), 
            .I3(GND_net), .O(n3096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2095_3_lut (.I0(n3001), .I1(n3050[14]), .I2(n3017), 
            .I3(GND_net), .O(n3100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_2_lut (.I0(n3094), .I1(n3103), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_5247));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1633 (.I0(n3100), .I1(n3106), .I2(n3096), .I3(n3093), 
            .O(n46_adj_5248));
    defparam i19_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1634 (.I0(n3085), .I1(n3087), .I2(n3086), .I3(n3088), 
            .O(n42_adj_5249));
    defparam i15_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[4]), .I1(n3099), .I2(n3109), .I3(GND_net), 
            .O(n33_adj_5250));
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1635 (.I0(n3089), .I1(n3091), .I2(n3090), .I3(n3104), 
            .O(n43_adj_5251));
    defparam i16_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1636 (.I0(n3095), .I1(n46_adj_5248), .I2(n36_adj_5247), 
            .I3(n3097), .O(n50));
    defparam i23_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1637 (.I0(n3108), .I1(n42_adj_5249), .I2(n3084), 
            .I3(n3083), .O(n48_adj_5252));
    defparam i21_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1638 (.I0(n43_adj_5251), .I1(n33_adj_5250), .I2(n3105), 
            .I3(n3092), .O(n49_adj_5253));
    defparam i22_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1639 (.I0(n3107), .I1(n3101), .I2(n3102), .I3(n3098), 
            .O(n47_adj_5254));
    defparam i20_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1640 (.I0(n47_adj_5254), .I1(n49_adj_5253), .I2(n48_adj_5252), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2101_3_lut (.I0(n3007), .I1(n3050[8]), .I2(n3017), 
            .I3(GND_net), .O(n3106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2166_3_lut (.I0(n3104), .I1(n3149[10]), .I2(n3116), 
            .I3(GND_net), .O(n21_adj_5255));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2164_3_lut (.I0(n3102), .I1(n3149[12]), .I2(n3116), 
            .I3(GND_net), .O(n25_adj_5256));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2171_3_lut (.I0(n3109), .I1(n3149[5]), .I2(n3116), 
            .I3(GND_net), .O(n11_adj_5257));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1641 (.I0(n3106), .I1(n11_adj_5257), .I2(n3149[8]), 
            .I3(n3116), .O(n49309));
    defparam i1_4_lut_adj_1641.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2169_3_lut (.I0(n3107), .I1(n3149[7]), .I2(n3116), 
            .I3(GND_net), .O(n15_adj_5258));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2162_3_lut (.I0(n3100), .I1(n3149[14]), .I2(n3116), 
            .I3(GND_net), .O(n29_adj_5259));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(n3103), .I1(n29_adj_5259), .I2(n3149[11]), 
            .I3(n3116), .O(n49313));
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(n3101), .I1(n15_adj_5258), .I2(n3149[13]), 
            .I3(n3116), .O(n49315));
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1644 (.I0(n3108), .I1(n21_adj_5255), .I2(n3149[6]), 
            .I3(n3116), .O(n49317));
    defparam i1_4_lut_adj_1644.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(n3105), .I1(n25_adj_5256), .I2(n3149[9]), 
            .I3(n3116), .O(n49311));
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n49309), .I1(n3099), .I2(n3149[15]), 
            .I3(n3116), .O(n49319));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hfaee;
    SB_LUT4 mod_5_i2160_3_lut (.I0(n3098), .I1(n3149[16]), .I2(n3116), 
            .I3(GND_net), .O(n33_adj_5260));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(bit_ctr[3]), .I1(n49315), .I2(n3209), 
            .I3(n49313), .O(n49327));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'hffec;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n33_adj_5260), .I1(n49319), .I2(n49311), 
            .I3(n49317), .O(n49329));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2159_3_lut (.I0(n3097), .I1(n3149[17]), .I2(n3116), 
            .I3(GND_net), .O(n35_adj_5261));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2158_3_lut (.I0(n3096), .I1(n3149[18]), .I2(n3116), 
            .I3(GND_net), .O(n37_adj_5262));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n37_adj_5262), .I1(n35_adj_5261), .I2(n49329), 
            .I3(n49327), .O(n49335));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n3095), .I1(n49335), .I2(n3149[19]), 
            .I3(n3116), .O(n49337));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n3094), .I1(n49337), .I2(n3149[20]), 
            .I3(n3116), .O(n49339));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n3093), .I1(n49339), .I2(n3149[21]), 
            .I3(n3116), .O(n49341));
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n3092), .I1(n49341), .I2(n3149[22]), 
            .I3(n3116), .O(n49343));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n3091), .I1(n49343), .I2(n3149[23]), 
            .I3(n3116), .O(n49345));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n3090), .I1(n49345), .I2(n3149[24]), 
            .I3(n3116), .O(n49347));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1656 (.I0(n3089), .I1(n49347), .I2(n3149[25]), 
            .I3(n3116), .O(n49349));
    defparam i1_4_lut_adj_1656.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n3088), .I1(n49349), .I2(n3149[26]), 
            .I3(n3116), .O(n49351));
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1658 (.I0(n3087), .I1(n49351), .I2(n3149[27]), 
            .I3(n3116), .O(n49353));
    defparam i1_4_lut_adj_1658.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n3086), .I1(n49353), .I2(n3149[28]), 
            .I3(n3116), .O(n49355));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2147_3_lut (.I0(n3085), .I1(n3149[29]), .I2(n3116), 
            .I3(GND_net), .O(n59));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2146_3_lut (.I0(n3084), .I1(n3149[30]), .I2(n3116), 
            .I3(GND_net), .O(n61));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1660 (.I0(n61), .I1(n50010), .I2(n59), .I3(n49355), 
            .O(n42573));
    defparam i1_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2172_3_lut (.I0(bit_ctr[4]), .I1(n3149[4]), .I2(n3116), 
            .I3(GND_net), .O(n3209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35579_2_lut (.I0(state[1]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n51034));   // verilog/neopixel.v(16[20:25])
    defparam i35579_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24_4_lut_adj_1661 (.I0(n38635), .I1(n38574), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[1]), .O(n10_adj_5263));   // verilog/neopixel.v(16[20:25])
    defparam i24_4_lut_adj_1661.LUT_INIT = 16'h0ac0;
    SB_LUT4 i23_4_lut_adj_1662 (.I0(n10_adj_5263), .I1(n51034), .I2(state[0]), 
            .I3(n98), .O(n38562));   // verilog/neopixel.v(16[20:25])
    defparam i23_4_lut_adj_1662.LUT_INIT = 16'h0aca;
    SB_LUT4 i35773_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n42573), .I3(GND_net), 
            .O(color_bit_N_722[4]));
    defparam i35773_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i35946_3_lut (.I0(n52813), .I1(bit_ctr[3]), .I2(n42573), .I3(GND_net), 
            .O(n51115));
    defparam i35946_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i36428_4_lut (.I0(n52771), .I1(n128), .I2(n51115), .I3(color_bit_N_722[4]), 
            .O(state_3__N_528[0]));   // verilog/neopixel.v(18[12:19])
    defparam i36428_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mod_5_i875_3_lut (.I0(n1205), .I1(n1268[28]), .I2(n1235), 
            .I3(GND_net), .O(n1304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i876_3_lut (.I0(n1206), .I1(n1268[27]), .I2(n1235), 
            .I3(GND_net), .O(n1305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i873_3_lut (.I0(n1203), .I1(n1268[30]), .I2(n1235), 
            .I3(GND_net), .O(n1302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i880_3_lut (.I0(bit_ctr[23]), .I1(n1268[23]), .I2(n1235), 
            .I3(GND_net), .O(n1309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i874_3_lut (.I0(n1204), .I1(n1268[29]), .I2(n1235), 
            .I3(GND_net), .O(n1303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i808_3_lut (.I0(n1106), .I1(n1169[28]), .I2(n1136), 
            .I3(GND_net), .O(n1205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i807_3_lut (.I0(n1105), .I1(n1169[29]), .I2(n1136), 
            .I3(GND_net), .O(n1204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i806_3_lut (.I0(n1104), .I1(n1169[30]), .I2(n1136), 
            .I3(GND_net), .O(n1203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i811_3_lut (.I0(n1109), .I1(n1169[25]), .I2(n1136), 
            .I3(GND_net), .O(n1208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i809_3_lut (.I0(n1107), .I1(n1169[27]), .I2(n1136), 
            .I3(GND_net), .O(n1206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i810_3_lut (.I0(n1108), .I1(n1169[26]), .I2(n1136), 
            .I3(GND_net), .O(n1207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_1663 (.I0(bit_ctr[23]), .I1(n1207), .I2(n1209), 
            .I3(GND_net), .O(n11_adj_5264));
    defparam i3_3_lut_adj_1663.LUT_INIT = 16'hecec;
    SB_LUT4 i5_4_lut_adj_1664 (.I0(n1203), .I1(n1204), .I2(n1202), .I3(n1205), 
            .O(n13_adj_5265));
    defparam i5_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1665 (.I0(n13_adj_5265), .I1(n11_adj_5264), .I2(n1206), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i812_3_lut (.I0(bit_ctr[24]), .I1(n1169[24]), .I2(n1136), 
            .I3(GND_net), .O(n1209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i879_3_lut (.I0(n1209), .I1(n1268[24]), .I2(n1235), 
            .I3(GND_net), .O(n1308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i878_3_lut (.I0(n1208), .I1(n1268[25]), .I2(n1235), 
            .I3(GND_net), .O(n1307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i877_3_lut (.I0(n1207), .I1(n1268[26]), .I2(n1235), 
            .I3(GND_net), .O(n1306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1666 (.I0(n1302), .I1(n1301), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5266));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_adj_1666.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1667 (.I0(n1306), .I1(n1307), .I2(n1308), .I3(n10_adj_5266), 
            .O(n16_adj_5267));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1668 (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), 
            .I3(GND_net), .O(n11_adj_5268));   // verilog/neopixel.v(22[26:36])
    defparam i2_3_lut_adj_1668.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1669 (.I0(n11_adj_5268), .I1(n16_adj_5267), .I2(n1305), 
            .I3(n1304), .O(n1334));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n38635), .I1(state[1]), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n48388));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i30876_2_lut_3_lut (.I0(start), .I1(one_wire_N_679[10]), .I2(n121), 
            .I3(GND_net), .O(n46444));
    defparam i30876_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_i741_3_lut (.I0(n1007), .I1(n1070[28]), .I2(n1037), 
            .I3(GND_net), .O(n1106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i742_3_lut (.I0(n1008), .I1(n1070[27]), .I2(n1037), 
            .I3(GND_net), .O(n1107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i743_3_lut (.I0(n1009), .I1(n1070[26]), .I2(n1037), 
            .I3(GND_net), .O(n1108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i740_3_lut (.I0(n1006), .I1(n1070[29]), .I2(n1037), 
            .I3(GND_net), .O(n1105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i744_3_lut (.I0(bit_ctr[25]), .I1(n1070[25]), .I2(n1037), 
            .I3(GND_net), .O(n1109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i739_3_lut (.I0(n1005), .I1(n1070[30]), .I2(n1037), 
            .I3(GND_net), .O(n1104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(n1105), .I1(n1108), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5269));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1670 (.I0(bit_ctr[24]), .I1(n10_adj_5269), .I2(n1104), 
            .I3(n1109), .O(n12_adj_5270));
    defparam i5_4_lut_adj_1670.LUT_INIT = 16'hfefc;
    SB_LUT4 i6_4_lut_adj_1671 (.I0(n1107), .I1(n12_adj_5270), .I2(n1106), 
            .I3(n1103), .O(n1136));
    defparam i6_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_37218 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n52732));
    defparam bit_ctr_0__bdd_4_lut_37218.LUT_INIT = 16'he4aa;
    SB_LUT4 n52732_bdd_4_lut (.I0(n52732), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n52735));
    defparam n52732_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Ki[2] , \Ki[0] , \Ki[1] , \Ki[3] , 
            PWMLimit, \Ki[6] , \Ki[4] , \Ki[5] , \Kp[5] , \Kp[1] , 
            \Kp[0] , \Kp[2] , \Kp[3] , \Kp[4] , \Kp[6] , \Kp[7] , 
            \Kp[8] , \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , 
            \Kp[14] , \Kp[15] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , 
            \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , IntegralLimit, 
            VCC_net, setpoint, motor_state, duty, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Ki[2] ;
    input \Ki[0] ;
    input \Ki[1] ;
    input \Ki[3] ;
    input [23:0]PWMLimit;
    input \Ki[6] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Kp[5] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]IntegralLimit;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output [23:0]duty;
    input clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [14:0]n17673;
    wire [13:0]n18153;
    
    wire n974, n40851, n40852;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3672 ;
    
    wire n204;
    wire [1:0]n20377;
    
    wire n901, n40850, n828, n40849, n131, n62, n40657;
    wire [23:0]n1;
    
    wire n40658, n4;
    wire [2:0]n20353;
    wire [3:0]n20313;
    
    wire n40747;
    wire [7:0]n19913;
    
    wire n262, n40748;
    wire [23:0]n1_adj_5153;
    
    wire n490, n12, n6, n8, n11, n6_adj_4731, n7, n40656;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n40134, n18, n13, n4_adj_4732, n47913, n755, n40848;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n40528;
    wire [8:0]n19733;
    
    wire n189, n40746;
    wire [23:0]n34;
    
    wire n414, n80, n11_adj_4733, n153, n226, n299, n372, n122, 
        n53, n445, n518, n591, n664, n737, n810, n883, n956, 
        n1029, n1102, n487, \PID_CONTROLLER.integral_23__N_3720 ;
    wire [23:0]n4230;
    
    wire n560, n195, n101, n32, n74, n268, n5, n147, n220, 
        n293, n366, n439, n512, n585, n174, n247, n658, n731, 
        n804, n877, n950, n1023, n40225, n4_adj_4736, n1096, n341, 
        n320, n414_adj_4737, n393, n466, n682, n40847, n77, n8_adj_4738, 
        n150, n223, n296, n369, n442, n539, n515, n588, n661, 
        n734, n487_adj_4739, n807, n880, n953, n1026, n612, n1099, 
        n560_adj_4741, n17, n9, n11_adj_4742, n51218, n51215;
    wire [4:0]n20253;
    
    wire n53201, n51694, n51503, n53183, n51498, n51496, n53176, 
        n27, n15, n13_adj_4743, n11_adj_4744, n51147, n21_adj_4745, 
        n19, n17_adj_4746, n9_adj_4747, n51154, n43, n16, n51430, 
        n8_adj_4748, n45, n24_adj_4749, n5_adj_4750, n51166, n51469, 
        n51465, n25_adj_4751, n23_adj_4752, n51858, n31, n29, n51670, 
        n37, n35, n33, n51912, n51515, n53170, n47, n116, n51489, 
        n53164, n12_adj_4754, n51184, n53188, n10_adj_4756, n30, 
        n609, n40846, n51792, n51196, n53168, n51688, n53194, 
        n51864, n53159, n51953, n53156, n16_adj_4759, n51169, n40655, 
        n110, n24_adj_4762, n6_adj_4763, n41, n51878, n51879, n51172, 
        n8_adj_4765, n53154, n51804, n51799;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3723 ;
    
    wire n3, n4_adj_4766, n51866, n51867, n12_adj_4767, n51448, 
        n10_adj_4768, n30_adj_4769, n51140, n536, n40845, n51939, 
        n28, n51967, n51968, n39, n51942, n6_adj_4770, n51868, 
        n183, n51869, n256, n51432, n329, n51810, n51807, n41_adj_4774, 
        n51434, n51924, n51526, n51926, n402, n4_adj_4775, n51872, 
        n475, n51873, n51186, n548, n51951, n51801, n51983, n51984, 
        n51964, n51174, n51882, n463, n40844, n40, \PID_CONTROLLER.integral_23__N_3722 , 
        n51884;
    wire [23:0]duty_23__N_3772;
    wire [23:0]n257;
    
    wire n51387, n40654, n621, n694, n390, n40843, n6_adj_4783, 
        n767;
    wire [6:0]n20057;
    
    wire n630, n40745, n51428, n557, n40744, n840, n6_adj_4786, 
        n125, n56, n198, n271, n317, n40842, n74_adj_4790, n344, 
        n5_adj_4791, n417, n119, n50, n147_adj_4792, n220_adj_4793, 
        n293_adj_4794, n685, n366_adj_4795, n192, n137;
    wire [1:0]n20385;
    
    wire n40268;
    wire [2:0]n20368;
    
    wire n439_adj_4796, n4_adj_4797;
    wire [3:0]n20337;
    
    wire n490_adj_4799, n4_adj_4800, n40653, n6_adj_4801, n8_adj_4802, 
        n14_adj_4803, n12_adj_4804, n11_adj_4805, n484, n40743, n15_adj_4806, 
        n244, n40841, n40652, n17_adj_4807;
    wire [23:0]duty_23__N_3648;
    
    wire n48333, n171, n40840, n29_adj_4808, n98, n107, n38, n40651;
    wire [12:0]n18573;
    
    wire n1050, n40839, n411, n40742, n977, n40838, n904, n40837, 
        n180, n253, n338, n40741;
    wire [0:0]n10669;
    wire [21:0]n11176;
    
    wire n41502, n41501, n41500, n40650, n512_adj_4810, n41499, 
        n585_adj_4812, n265, n40740, n41498, n41497, n326, n399, 
        n41496, n658_adj_4816, n731_adj_4817, n804_adj_4818, n41495, 
        n831, n40836, n877_adj_4819, n1096_adj_4820, n41494, n1023_adj_4821, 
        n41493, n758, n950_adj_4822, n41492, n40835, n41491, n41490, 
        n41489, n41488, n41487, n41486, n41485, n40739, n41484, 
        n40834, n41483, n41482, n41481, n40649, n472;
    wire [20:0]n13140;
    
    wire n41480, n41479, n40578, n41478, n40648, n41477, n41476, 
        n41475, n545, n41474;
    wire [5:0]n20169;
    
    wire n40738, n41473, n40577, n40833, n41472, n41471, n41470, 
        n41469, n618, n40737, n41468, n41467, n41466, n40647, 
        n41465, n40832, n41464, n41463, n691, n110_adj_4830, n41_adj_4832, 
        n183_adj_4833, n256_adj_4834, n329_adj_4835, n402_adj_4836, 
        n41462, n41461, n41460, n40646, n475_adj_4838, n764, n548_adj_4839, 
        n621_adj_4840, n40645, n40831, n40830, n40736, n694_adj_4842, 
        n767_adj_4843, n840_adj_4844, n40829, n40735, n40576, n40828, 
        n40827, n40644, n40734, n40733, n40643;
    wire [6:0]n20120;
    wire [5:0]n20217;
    
    wire n40826, n40575, n40825;
    wire [19:0]n14671;
    
    wire n41436, n41435, n335, n41434, n41433, n41432, n408, n41431, 
        n41430, n1047, n41429, n41428, n41427, n41426, n41425, 
        n41424, n41423, n1120, n41422, n41421, n481, n41420, n41419, 
        n119_adj_4848, n50_adj_4849, n41418, n41417, n40642;
    wire [18:0]n15472;
    
    wire n41416, n41415, n41414, n40824, n41413, n41412, n40732, 
        n1105, n41411, n417_adj_4852, n40731, n341_adj_4853, n40823, 
        n1032, n41410, n192_adj_4854, n268_adj_4855, n40822, n959, 
        n41409, n40574, n886, n41408, n265_adj_4856, n338_adj_4858, 
        n411_adj_4859, n484_adj_4860, n557_adj_4862, n813, n41407, 
        n630_adj_4863, n740, n41406, n667, n41405, n344_adj_4864, 
        n40730, n95, n594, n41404, n26_adj_4865, n521, n41403, 
        n168, n241, n448, n41402, n375, n41401, n302, n41400, 
        n314, n40573, n229, n41399, n271_adj_4866, n40729, n387, 
        n156, n41398, n460, n14_adj_4867, n83, n533;
    wire [17:0]n16193;
    
    wire n41397, n41396, n40641, n41395, n554, n606, n41394, n1108, 
        n41393, n40572, n1035, n41392, n679, n40640, n962, n41391, 
        n889, n41390, n752, n816, n41389, n825, n898, n627, 
        n971, n743, n41388, n1044, n670, n41387, n700, n597, 
        n41386, n524, n41385, n451, n41384, n378, n41383, n1117, 
        n305, n41382, n92, n23_adj_4869, n232, n41381, n113, n159, 
        n41380, n44, n165, n238, n195_adj_4871, n40821, n311, 
        n384, n17_adj_4872, n86;
    wire [16:0]n16840;
    
    wire n41379, n198_adj_4873, n40728, n41378, n457, n40571, n41377, 
        n1111, n41376, n1038, n41375, n965, n41374, n530, n892, 
        n41373, n603, n676, n819, n41372, n749, n822, n895, 
        n968, n1041, n746, n41371, n186, n1114, n116_adj_4876, 
        n673, n41370, n47_adj_4877, n600, n41369, n189_adj_4878, 
        n527, n41368, n262_adj_4880, n335_adj_4881, n454, n41367, 
        n381, n41366, n408_adj_4882, n308, n41365, n40639, n481_adj_4883, 
        n235, n41364, n554_adj_4884, n162, n41363, n627_adj_4885, 
        n56_adj_4886, n125_adj_4887, n53_adj_4888, n122_adj_4889, n700_adj_4890, 
        n20_adj_4891, n89, n89_adj_4892;
    wire [15:0]n17417;
    
    wire n41362, n40638, n41361, n20_adj_4893, n162_adj_4894, n259, 
        n1114_adj_4895, n41360, n1041_adj_4896, n41359, n968_adj_4897, 
        n41358, n895_adj_4898, n41357, n822_adj_4899, n41356, n235_adj_4900, 
        n749_adj_4901, n41355, n676_adj_4902, n41354, n603_adj_4903, 
        n41353, n530_adj_4905, n41352, n457_adj_4906, n41351, n308_adj_4907, 
        n381_adj_4908, n384_adj_4909, n41350, n311_adj_4910, n41349, 
        n454_adj_4912, n527_adj_4913, n238_adj_4914, n41348, n165_adj_4915, 
        n41347, n332, n23_adj_4916, n92_adj_4917, n40637, n40636;
    wire [14:0]n17928;
    
    wire n41346, n40570, n1117_adj_4918, n41345, n40635, n1044_adj_4919, 
        n41344, n600_adj_4920, n673_adj_4921, n971_adj_4922, n41343, 
        n898_adj_4923, n41342, n825_adj_4924, n41341, n40634, n746_adj_4925, 
        n819_adj_4926, n892_adj_4927, n405, n965_adj_4929, n1038_adj_4930, 
        n478, n1111_adj_4931, n86_adj_4932, n17_adj_4933, n551, n159_adj_4934, 
        n232_adj_4936, n41_adj_4937, n39_adj_4938, n305_adj_4939, n45_adj_4940, 
        n43_adj_4941, n23_adj_4942, n25_adj_4943, n37_adj_4944, n752_adj_4945, 
        n41340, n378_adj_4946, n29_adj_4947, n31_adj_4948, n35_adj_4949, 
        n679_adj_4950, n41339, n451_adj_4951, n524_adj_4952, n11_adj_4953, 
        n13_adj_4954, n15_adj_4955, n27_adj_4956, n597_adj_4958, n670_adj_4959, 
        n743_adj_4960, n606_adj_4961, n41338, n816_adj_4962, n33_adj_4963, 
        n9_adj_4964, n17_adj_4965, n19_adj_4966, n533_adj_4967, n41337, 
        n460_adj_4968, n41336, n21_adj_4969, n51418, n889_adj_4970, 
        n624, n387_adj_4971, n41335, n40633, n51411, n962_adj_4972, 
        n12_adj_4973, n314_adj_4974, n41334, n10_adj_4975, n30_adj_4976, 
        n241_adj_4977, n41333, n51652, n51648, n51910, n51764, n51947, 
        n697, n1035_adj_4978, n1108_adj_4979, n168_adj_4980, n41332, 
        n26_adj_4981, n95_adj_4982, n16_adj_4983, n51834, n51835, 
        n8_adj_4984, n24_adj_4985, n51392, n770, n51389, n51812, 
        n51528, n113_adj_4986, n44_adj_4987, n186_adj_4988, n4_adj_4989, 
        n51832, n51833, n51405, n259_adj_4990, n51402, n51914, n51530, 
        n51981, n51982, n332_adj_4991, n405_adj_4992, n51970, n51394, 
        n51928, n51536, n51930, duty_23__N_3771, n39_adj_4994, n41_adj_4995, 
        n478_adj_4996, n551_adj_4997, n624_adj_4999, n45_adj_5001, n43_adj_5002, 
        n697_adj_5004, n770_adj_5005, n83_adj_5007, n23_adj_5008, n40632, 
        n25_adj_5009, n37_adj_5010, n29_adj_5011, n31_adj_5012, n35_adj_5013, 
        n33_adj_5015, n14_adj_5016, n11_adj_5017, n13_adj_5018, n156_adj_5019, 
        n15_adj_5020, n27_adj_5022, n9_adj_5023, n17_adj_5024, n19_adj_5025, 
        n21_adj_5027, n229_adj_5028, n40569, n51377, n51371, n12_adj_5030, 
        n302_adj_5031, n375_adj_5033, n10_adj_5034, n837, n30_adj_5035, 
        n51620, n51616, n51904, n910, n51746, n51945, n16_adj_5036, 
        n107_adj_5037, n38_adj_5038, n51828, n51829, n8_adj_5039, 
        n24_adj_5040, n51354, n51352, n51814, n51538, n104, n4_adj_5041, 
        n40631, n35_adj_5042, n51826, n51827, n51367, n51365, n51916, 
        n51540, n51961, n51962, n51960, n51357, n51932, n51546, 
        n51934, n256_adj_5043;
    wire [23:0]duty_23__N_3747;
    
    wire n40568;
    wire [11:0]n18937;
    
    wire n980, n40813;
    wire [13:0]n18377;
    
    wire n1120_adj_5044, n41309, n907, n40812, n1047_adj_5045, n41308, 
        n974_adj_5046, n41307, n901_adj_5047, n41306, n834, n40811, 
        n828_adj_5048, n41305, n755_adj_5049, n41304, n682_adj_5050, 
        n41303, n609_adj_5051, n41302, n536_adj_5052, n41301, n463_adj_5053, 
        n41300, n390_adj_5054, n41299, n317_adj_5055, n41298, n244_adj_5056, 
        n41297, n171_adj_5057, n41296, n761, n40810, n29_adj_5058, 
        n98_adj_5059, n688, n40809;
    wire [12:0]n18768;
    
    wire n1050_adj_5060, n41295, n977_adj_5061, n41294, n904_adj_5062, 
        n41293, n831_adj_5063, n41292, n758_adj_5064, n41291, n685_adj_5065, 
        n41290, n612_adj_5066, n41289, n539_adj_5067, n41288, n615, 
        n40808, n466_adj_5068, n41287, n393_adj_5069, n41286, n40567, 
        n320_adj_5070, n41285, n247_adj_5071, n41284, n542, n40807, 
        n174_adj_5072, n41283, n32_adj_5073, n101_adj_5074;
    wire [11:0]n19105;
    
    wire n980_adj_5075, n41282, n907_adj_5076, n41281, n469, n40806, 
        n834_adj_5077, n41280, n761_adj_5078, n41279, n688_adj_5079, 
        n41278, n615_adj_5080, n41277, n542_adj_5081, n41276, n469_adj_5082, 
        n41275, n396, n41274, n323, n41273, n250, n41272, n177, 
        n41271, n35_adj_5083, n104_adj_5084;
    wire [10:0]n19392;
    
    wire n910_adj_5085, n41270, n396_adj_5086, n40805, n837_adj_5087, 
        n41269, n764_adj_5088, n41268, n691_adj_5089, n41267, n618_adj_5090, 
        n41266, n545_adj_5091, n41265, n472_adj_5092, n41264, n323_adj_5093, 
        n40804, n399_adj_5094, n41263, n326_adj_5095, n41262, n250_adj_5096, 
        n40803, n253_adj_5097, n41261, n177_adj_5098, n40802, n180_adj_5099, 
        n41260;
    wire [10:0]n19249;
    
    wire n40801, n40800;
    wire [9:0]n19633;
    
    wire n41238, n41237, n41236, n41235, n41234, n40799, n41233, 
        n40566, n41232, n41231, n41230, n41229, n40798, n40797, 
        n40565, n40796, n40564, n40563, n40795, n40562, n40794, 
        n40561, n40793, n40560, n40792, n40791, n40559, n40558, 
        n40557, n40790;
    wire [4:0]n20288;
    
    wire n40789, n40699, n40788, n40698, n40556, n40787, n40786;
    wire [9:0]n19513;
    
    wire n40785, n40784, n40697, n40696, n40783, n40695, n40150, 
        n40782, n40694, n40693, n40781;
    wire [0:0]n10138;
    
    wire n40550, n40692, n40780, n40549, n40779, n40778, n40691, 
        n40690, n40548, n40777, n40689, n40776, n40547, n40688, 
        n40687, n40686, n40685, n40546, n40684, n448_adj_5101, n521_adj_5103, 
        n40683, n40545, n40544, n594_adj_5105, n40682, n40543, n40542, 
        n40541, n40540;
    wire [21:0]n10645;
    
    wire n41033, n41032, n41031, n41030, n41029, n41028, n41027, 
        n41026, n41025, n41024, n41023, n41022, n41021, n41020, 
        n41019, n41018, n41017, n41016, n41015, n41014, n41013, 
        n41012, n40681, n40539, n40538;
    wire [20:0]n12653;
    
    wire n41003, n41002, n41001, n40680, n40679, n40537, n41000, 
        n40999, n40998, n40997, n1099_adj_5112, n40996, n1026_adj_5113, 
        n40995, n953_adj_5114, n40994, n880_adj_5115, n40993, n807_adj_5116, 
        n40992, n734_adj_5117, n40991, n661_adj_5118, n40990, n588_adj_5119, 
        n40989, n515_adj_5120, n40988, n442_adj_5121, n40987, n369_adj_5122, 
        n40986, n296_adj_5123, n40985, n223_adj_5124, n40984, n150_adj_5125, 
        n40983, n8_adj_5126, n77_adj_5127;
    wire [19:0]n14231;
    
    wire n40982, n40981, n40980, n40979, n40978, n40977, n1102_adj_5128, 
        n40976, n1029_adj_5129, n40975, n956_adj_5130, n40974, n883_adj_5131, 
        n40973, n810_adj_5132, n40972, n737_adj_5133, n40971, n664_adj_5134, 
        n40970, n591_adj_5135, n40969, n518_adj_5136, n40968, n445_adj_5137, 
        n40967, n372_adj_5138, n40966, n299_adj_5139, n40965, n226_adj_5140, 
        n40964, n153_adj_5141, n40963, n11_adj_5142, n80_adj_5143;
    wire [18:0]n15073;
    
    wire n40962, n40961, n40960, n40959, n40958, n1105_adj_5144, 
        n40957, n1032_adj_5145, n40956, n959_adj_5146, n40955, n886_adj_5147, 
        n40954, n813_adj_5148, n40953, n740_adj_5149, n40952, n667_adj_5150, 
        n40951, n40950, n40949, n40678, n40948, n40947, n40677, 
        n40946, n40945, n40944, n40536, n40676;
    wire [8:0]n19832;
    
    wire n40943, n40942, n40675, n40941, n40535, n40674, n40940, 
        n40939, n40938, n40937, n40936, n40935;
    wire [17:0]n15833;
    
    wire n40934, n40933, n40762, n40932, n40931, n40930, n40929, 
        n40761, n40534, n40928, n40760, n40927, n40926, n40925, 
        n40924, n40923, n40673, n40922, n40921, n40920, n40919, 
        n40533, n40918, n40672, n40917, n40759;
    wire [16:0]n16517;
    
    wire n40916, n40915, n40914, n40913, n40758, n40912, n40532, 
        n40911, n40671, n40757, n40910, n40909, n40908, n40907, 
        n40906, n40756, n40905, n40904, n40670, n40903, n40902, 
        n40669, n40901, n40755, n40900;
    wire [7:0]n19993;
    
    wire n40899, n40898, n40897, n40896, n40895, n40894, n40893, 
        n40668, n40892;
    wire [15:0]n17129;
    
    wire n40891, n40890, n40889, n40754, n40888, n40887, n40886, 
        n40885, n40884, n40883, n40882, n40667, n40881, n40666, 
        n40880, n40879, n40878, n40877, n40876, n40665, n40875, 
        n40874, n40753, n40873, n40872, n40752, n40871, n40664, 
        n40870, n40869, n40868, n40867, n40751, n40531, n40866, 
        n40530, n40865, n40864, n40863, n40529, n40862, n40861, 
        n40860, n40859, n40663, n40858, n40857, n40856, n40662, 
        n40855, n40854, n40661, n40660, n40750, n40659, n40853, 
        n40749, n6_adj_5151, n4_adj_5152, n40293, n40327;
    
    SB_LUT4 add_6621_14_lut (.I0(GND_net), .I1(n18153[11]), .I2(n974), 
            .I3(n40851), .O(n17673[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6621_14 (.CI(n40851), .I0(n18153[11]), .I1(n974), .CO(n40852));
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26472_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n20377[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26472_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_6621_13_lut (.I0(GND_net), .I1(n18153[10]), .I2(n901), 
            .I3(n40850), .O(n17673[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6621_13 (.CI(n40850), .I0(n18153[10]), .I1(n901), .CO(n40851));
    SB_LUT4 add_6621_12_lut (.I0(GND_net), .I1(n18153[9]), .I2(n828), 
            .I3(n40849), .O(n17673[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n40657), .I0(GND_net), .I1(n1[4]), 
            .CO(n40658));
    SB_LUT4 i2_4_lut (.I0(n4), .I1(\Ki[3] ), .I2(n20353[1]), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n20313[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_CARRY add_6765_4 (.CI(n40747), .I0(n19913[1]), .I1(n262), .CO(n40748));
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6621_12 (.CI(n40849), .I0(n18153[9]), .I1(n828), .CO(n40850));
    SB_LUT4 i2_4_lut_adj_1515 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [20]), .O(n12));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1515.LUT_INIT = 16'h9c50;
    SB_LUT4 i26585_4_lut (.I0(n20313[2]), .I1(\Ki[4] ), .I2(n6), .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .O(n8));   // verilog/motorControl.v(34[25:36])
    defparam i26585_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n11));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i26546_4_lut (.I0(n20353[1]), .I1(\Ki[3] ), .I2(n4), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n6_adj_4731));   // verilog/motorControl.v(34[25:36])
    defparam i26546_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n40656), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26474_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n40134));   // verilog/motorControl.v(34[25:36])
    defparam i26474_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4731), .I1(n11), .I2(n8), .I3(n12), 
            .O(n18));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [22]), .O(n13));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n40134), .I3(n4_adj_4732), 
            .O(n47913));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6621_11_lut (.I0(GND_net), .I1(n18153[8]), .I2(n755), 
            .I3(n40848), .O(n17673[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6621_11 (.CI(n40848), .I0(n18153[8]), .I1(n755), .CO(n40849));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n40656), .I0(GND_net), .I1(n1[3]), 
            .CO(n40657));
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n40528));
    SB_LUT4 add_6765_3_lut (.I0(GND_net), .I1(n19913[0]), .I2(n189), .I3(n40746), 
            .O(n19733[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4733));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22142_2_lut (.I0(n34[20]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22141_2_lut (.I0(n34[21]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22141_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26569_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n40225), .I3(n20313[0]), .O(n4_adj_4736));   // verilog/motorControl.v(34[25:36])
    defparam i26569_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6765_3 (.CI(n40746), .I0(n19913[0]), .I1(n189), .CO(n40747));
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6621_10_lut (.I0(GND_net), .I1(n18153[7]), .I2(n682), 
            .I3(n40847), .O(n17673[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n34[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4738));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4739));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22140_2_lut (.I0(n34[22]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4741));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4742));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35584_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n51218));
    defparam i35584_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i35581_3_lut (.I0(n11_adj_4742), .I1(n9), .I2(n51218), .I3(GND_net), 
            .O(n51215));
    defparam i35581_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i26556_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n20253[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26556_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i26558_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n40225));   // verilog/motorControl.v(34[25:36])
    defparam i26558_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_224_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n53201));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_224_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36059_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n53201), 
            .I2(IntegralLimit[7]), .I3(n51215), .O(n51694));
    defparam i36059_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35868_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n51694), .O(n51503));
    defparam i35868_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_206_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n53183));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_206_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35863_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n9), .O(n51498));
    defparam i35863_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35861_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n53183), 
            .I2(IntegralLimit[11]), .I3(n51498), .O(n51496));
    defparam i35861_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_199_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n53176));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_199_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35513_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_4743), .I3(n11_adj_4744), 
            .O(n51147));
    defparam i35513_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35520_4_lut (.I0(n21_adj_4745), .I1(n19), .I2(n17_adj_4746), 
            .I3(n9_adj_4747), .O(n51154));
    defparam i35520_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35796_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n51430));
    defparam i35796_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4746), .I3(GND_net), 
            .O(n8_adj_4748));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_4749));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35532_2_lut (.I0(n7), .I1(n5_adj_4750), .I2(GND_net), .I3(GND_net), 
            .O(n51166));
    defparam i35532_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35835_4_lut (.I0(n13_adj_4743), .I1(n11_adj_4744), .I2(n9_adj_4747), 
            .I3(n51166), .O(n51469));
    defparam i35835_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35831_4_lut (.I0(n19), .I1(n17_adj_4746), .I2(n15), .I3(n51469), 
            .O(n51465));
    defparam i35831_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36223_4_lut (.I0(n25_adj_4751), .I1(n23_adj_4752), .I2(n21_adj_4745), 
            .I3(n51465), .O(n51858));
    defparam i36223_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36035_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n51858), 
            .O(n51670));
    defparam i36035_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36277_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n51670), 
            .O(n51912));
    defparam i36277_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35880_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n53201), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4742), .O(n51515));
    defparam i35880_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_193_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n53170));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_193_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6621_10 (.CI(n40847), .I0(n18153[7]), .I1(n682), .CO(n40848));
    SB_LUT4 add_6765_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19733[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35854_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n53170), 
            .I2(IntegralLimit[14]), .I3(n51515), .O(n51489));
    defparam i35854_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_187_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n53164));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_187_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4754));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35550_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n51184));
    defparam i35550_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_211_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n53188));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_211_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4756));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4754), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6621_9_lut (.I0(GND_net), .I1(n18153[6]), .I2(n609), .I3(n40846), 
            .O(n17673[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36157_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n53183), 
            .I2(IntegralLimit[11]), .I3(n51503), .O(n51792));
    defparam i36157_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35562_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n53176), 
            .I2(IntegralLimit[13]), .I3(n51792), .O(n51196));
    defparam i35562_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_191_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n53168));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_191_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36053_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n53168), 
            .I2(IntegralLimit[15]), .I3(n51196), .O(n51688));
    defparam i36053_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_217_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n53194));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_217_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36229_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n53194), 
            .I2(IntegralLimit[17]), .I3(n51688), .O(n51864));
    defparam i36229_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_182_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n53159));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_182_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36318_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n53159), 
            .I2(IntegralLimit[19]), .I3(n51864), .O(n51953));
    defparam i36318_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_179_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n53156));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_179_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4759));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35535_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n51169));
    defparam i35535_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6765_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n40746));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n40655), .O(n5_adj_4750)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4759), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4762));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4763));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36243_3_lut (.I0(n6_adj_4763), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n51878));   // verilog/motorControl.v(31[10:34])
    defparam i36243_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36244_3_lut (.I0(n51878), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n51879));   // verilog/motorControl.v(31[10:34])
    defparam i36244_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6621_9 (.CI(n40846), .I0(n18153[6]), .I1(n609), .CO(n40847));
    SB_LUT4 i35538_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n53176), 
            .I2(IntegralLimit[21]), .I3(n51496), .O(n51172));
    defparam i35538_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i36169_4_lut (.I0(n24_adj_4762), .I1(n8_adj_4765), .I2(n53154), 
            .I3(n51169), .O(n51804));   // verilog/motorControl.v(31[10:34])
    defparam i36169_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36164_3_lut (.I0(n51879), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n51799));   // verilog/motorControl.v(31[10:34])
    defparam i36164_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3723 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4766));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i36231_3_lut (.I0(n4_adj_4766), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n51866));   // verilog/motorControl.v(31[38:63])
    defparam i36231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36232_3_lut (.I0(n51866), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n51867));   // verilog/motorControl.v(31[38:63])
    defparam i36232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4767));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35814_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n51448));
    defparam i35814_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4743), .I3(GND_net), 
            .O(n10_adj_4768));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4767), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_4769));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35506_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n51147), 
            .O(n51140));
    defparam i35506_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6621_8_lut (.I0(GND_net), .I1(n18153[5]), .I2(n536), .I3(n40845), 
            .O(n17673[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n40655), .I0(GND_net), .I1(n1[2]), 
            .CO(n40656));
    SB_LUT4 i36304_4_lut (.I0(n30_adj_4769), .I1(n10_adj_4768), .I2(n35), 
            .I3(n51448), .O(n51939));   // verilog/motorControl.v(31[38:63])
    defparam i36304_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36174_3_lut (.I0(n51867), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n28));   // verilog/motorControl.v(31[38:63])
    defparam i36174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36332_4_lut (.I0(n28), .I1(n51939), .I2(n35), .I3(n51140), 
            .O(n51967));   // verilog/motorControl.v(31[38:63])
    defparam i36332_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36333_3_lut (.I0(n51967), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n51968));   // verilog/motorControl.v(31[38:63])
    defparam i36333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36307_3_lut (.I0(n51968), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n51942));   // verilog/motorControl.v(31[38:63])
    defparam i36307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7), .I3(GND_net), 
            .O(n6_adj_4770));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36233_3_lut (.I0(n6_adj_4770), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4745), .I3(GND_net), .O(n51868));   // verilog/motorControl.v(31[38:63])
    defparam i36233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36234_3_lut (.I0(n51868), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4752), .I3(GND_net), .O(n51869));   // verilog/motorControl.v(31[38:63])
    defparam i36234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35798_4_lut (.I0(n43), .I1(n25_adj_4751), .I2(n23_adj_4752), 
            .I3(n51154), .O(n51432));
    defparam i35798_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36175_4_lut (.I0(n24_adj_4749), .I1(n8_adj_4748), .I2(n45), 
            .I3(n51430), .O(n51810));   // verilog/motorControl.v(31[38:63])
    defparam i36175_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36172_3_lut (.I0(n51869), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4751), .I3(GND_net), .O(n51807));   // verilog/motorControl.v(31[38:63])
    defparam i36172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35800_4_lut (.I0(n43), .I1(n41_adj_4774), .I2(n39), .I3(n51912), 
            .O(n51434));
    defparam i35800_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36289_4_lut (.I0(n51807), .I1(n51810), .I2(n45), .I3(n51432), 
            .O(n51924));   // verilog/motorControl.v(31[38:63])
    defparam i36289_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35891_3_lut (.I0(n51942), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4774), .I3(GND_net), .O(n51526));   // verilog/motorControl.v(31[38:63])
    defparam i35891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36291_4_lut (.I0(n51526), .I1(n51924), .I2(n45), .I3(n51434), 
            .O(n51926));   // verilog/motorControl.v(31[38:63])
    defparam i36291_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4775));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i36237_3_lut (.I0(n4_adj_4775), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n51872));   // verilog/motorControl.v(31[10:34])
    defparam i36237_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36238_3_lut (.I0(n51872), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n51873));   // verilog/motorControl.v(31[10:34])
    defparam i36238_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35552_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n53164), 
            .I2(IntegralLimit[16]), .I3(n51489), .O(n51186));
    defparam i35552_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36316_4_lut (.I0(n30), .I1(n10_adj_4756), .I2(n53188), .I3(n51184), 
            .O(n51951));   // verilog/motorControl.v(31[10:34])
    defparam i36316_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36166_3_lut (.I0(n51873), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n51801));   // verilog/motorControl.v(31[10:34])
    defparam i36166_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36348_4_lut (.I0(n51801), .I1(n51951), .I2(n53188), .I3(n51186), 
            .O(n51983));   // verilog/motorControl.v(31[10:34])
    defparam i36348_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36349_3_lut (.I0(n51983), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n51984));   // verilog/motorControl.v(31[10:34])
    defparam i36349_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36329_3_lut (.I0(n51984), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n51964));   // verilog/motorControl.v(31[10:34])
    defparam i36329_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35540_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n53156), 
            .I2(IntegralLimit[21]), .I3(n51953), .O(n51174));
    defparam i35540_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_177_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n53154));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_177_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6621_8 (.CI(n40845), .I0(n18153[5]), .I1(n536), .CO(n40846));
    SB_LUT4 i36247_4_lut (.I0(n51799), .I1(n51804), .I2(n53154), .I3(n51172), 
            .O(n51882));   // verilog/motorControl.v(31[10:34])
    defparam i36247_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6621_7_lut (.I0(GND_net), .I1(n18153[4]), .I2(n463), .I3(n40844), 
            .O(n17673[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36321_3_lut (.I0(n51964), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[10:34])
    defparam i36321_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36292_3_lut (.I0(n51926), .I1(\PID_CONTROLLER.integral_23__N_3723 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3722 ));   // verilog/motorControl.v(31[38:63])
    defparam i36292_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36249_4_lut (.I0(n40), .I1(n51882), .I2(n53154), .I3(n51174), 
            .O(n51884));   // verilog/motorControl.v(31[10:34])
    defparam i36249_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_850_4_lut  (.I0(n51884), .I1(\PID_CONTROLLER.integral_23__N_3722 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3720 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_850_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 i35753_3_lut_4_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3772[2]), .O(n51387));   // verilog/motorControl.v(38[19:35])
    defparam i35753_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6621_7 (.CI(n40844), .I0(n18153[4]), .I1(n463), .CO(n40845));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n40654), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n40654), .I0(GND_net), .I1(n1[1]), 
            .CO(n40655));
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3723 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6621_6_lut (.I0(GND_net), .I1(n18153[3]), .I2(n390), .I3(n40843), 
            .O(n17673[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4783));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22139_2_lut (.I0(n34[23]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22139_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6621_6 (.CI(n40843), .I0(n18153[3]), .I1(n390), .CO(n40844));
    SB_LUT4 add_6782_9_lut (.I0(GND_net), .I1(n20057[6]), .I2(n630), .I3(n40745), 
            .O(n19913[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35794_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(PWMLimit[2]), .O(n51428));   // verilog/motorControl.v(36[10:25])
    defparam i35794_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_6782_8_lut (.I0(GND_net), .I1(n20057[5]), .I2(n557), .I3(n40744), 
            .O(n19913[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n40654));
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(GND_net), .O(n6_adj_4786));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n34[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22018_2_lut (.I0(n34[0]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22018_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22161_2_lut (.I0(n34[1]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6621_5_lut (.I0(GND_net), .I1(n18153[2]), .I2(n317), .I3(n40842), 
            .O(n17673[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4790));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n34[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4791));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4792));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4793));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4794));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6782_8 (.CI(n40744), .I0(n20057[5]), .I1(n557), .CO(n40745));
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4795));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26510_3_lut (.I0(\Kp[0] ), .I1(n137), .I2(n34[22]), .I3(GND_net), 
            .O(n20385[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26510_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 i2_4_lut_adj_1516 (.I0(n40268), .I1(\Kp[2] ), .I2(n20385[0]), 
            .I3(n34[20]), .O(n20368[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1516.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4796));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1517 (.I0(n4_adj_4797), .I1(\Kp[3] ), .I2(n20368[1]), 
            .I3(n34[19]), .O(n20337[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1517.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(n34[21]), .I2(GND_net), 
            .I3(GND_net), .O(n137));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4799));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26608_4_lut (.I0(n20385[0]), .I1(\Kp[2] ), .I2(n40268), .I3(n34[20]), 
            .O(n4_adj_4800));   // verilog/motorControl.v(34[16:22])
    defparam i26608_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n40653), .O(n34[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26639_4_lut (.I0(n20368[1]), .I1(\Kp[3] ), .I2(n4_adj_4797), 
            .I3(n34[19]), .O(n6_adj_4801));   // verilog/motorControl.v(34[16:22])
    defparam i26639_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i4_4_lut (.I0(n8_adj_4802), .I1(\Kp[0] ), .I2(n137), .I3(n34[22]), 
            .O(n14_adj_4803));   // verilog/motorControl.v(34[16:22])
    defparam i4_4_lut.LUT_INIT = 16'h6aaa;
    SB_LUT4 i2_4_lut_adj_1518 (.I0(\Kp[3] ), .I1(\Kp[0] ), .I2(n34[20]), 
            .I3(n34[23]), .O(n12_adj_4804));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1518.LUT_INIT = 16'h93a0;
    SB_CARRY add_6621_5 (.CI(n40842), .I0(n18153[2]), .I1(n317), .CO(n40843));
    SB_LUT4 i1_4_lut_adj_1519 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n34[19]), 
            .I3(n34[21]), .O(n11_adj_4805));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1519.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_6782_7_lut (.I0(GND_net), .I1(n20057[4]), .I2(n484), .I3(n40743), 
            .O(n19913[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut (.I0(n4_adj_4800), .I1(\Kp[1] ), .I2(n34[22]), .I3(GND_net), 
            .O(n15_adj_4806));   // verilog/motorControl.v(34[16:22])
    defparam i5_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 add_6621_4_lut (.I0(GND_net), .I1(n18153[1]), .I2(n244), .I3(n40841), 
            .O(n17673[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n40652), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_4_lut (.I0(\Kp[5] ), .I1(n14_adj_4803), .I2(n6_adj_4801), 
            .I3(n34[18]), .O(n17_adj_4807));   // verilog/motorControl.v(34[16:22])
    defparam i7_4_lut.LUT_INIT = 16'h963c;
    SB_CARRY add_6621_4 (.CI(n40841), .I0(n18153[1]), .I1(n244), .CO(n40842));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3648[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i9_4_lut_adj_1520 (.I0(n17_adj_4807), .I1(n15_adj_4806), .I2(n11_adj_4805), 
            .I3(n12_adj_4804), .O(n48333));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY sub_3_add_2_24 (.CI(n40652), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n40653));
    SB_LUT4 add_6621_3_lut (.I0(GND_net), .I1(n18153[0]), .I2(n171), .I3(n40840), 
            .O(n17673[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6782_7 (.CI(n40743), .I0(n20057[4]), .I1(n484), .CO(n40744));
    SB_CARRY add_6621_3 (.CI(n40840), .I0(n18153[0]), .I1(n171), .CO(n40841));
    SB_LUT4 i22160_2_lut (.I0(n34[2]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22159_2_lut (.I0(n34[3]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6621_2_lut (.I0(GND_net), .I1(n29_adj_4808), .I2(n98), 
            .I3(GND_net), .O(n17673[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6621_2 (.CI(GND_net), .I0(n29_adj_4808), .I1(n98), .CO(n40840));
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n40651), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_15_lut (.I0(GND_net), .I1(n18573[12]), .I2(n1050), 
            .I3(n40839), .O(n18153[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6782_6_lut (.I0(GND_net), .I1(n20057[3]), .I2(n411), .I3(n40742), 
            .O(n19913[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_14_lut (.I0(GND_net), .I1(n18573[11]), .I2(n977), 
            .I3(n40838), .O(n18153[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_14 (.CI(n40838), .I0(n18573[11]), .I1(n977), .CO(n40839));
    SB_LUT4 add_6650_13_lut (.I0(GND_net), .I1(n18573[10]), .I2(n904), 
            .I3(n40837), .O(n18153[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_13 (.CI(n40837), .I0(n18573[10]), .I1(n904), .CO(n40838));
    SB_CARRY sub_3_add_2_23 (.CI(n40651), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n40652));
    SB_LUT4 i22158_2_lut (.I0(n34[4]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6782_6 (.CI(n40742), .I0(n20057[3]), .I1(n411), .CO(n40743));
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6782_5_lut (.I0(GND_net), .I1(n20057[2]), .I2(n338), .I3(n40741), 
            .O(n19913[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6782_5 (.CI(n40741), .I0(n20057[2]), .I1(n338), .CO(n40742));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n34[23]), .I1(n11176[21]), .I2(GND_net), 
            .I3(n41502), .O(n10669[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n11176[20]), .I2(GND_net), 
            .I3(n41501), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n41501), .I0(n11176[20]), .I1(GND_net), 
            .CO(n41502));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n11176[19]), .I2(GND_net), 
            .I3(n41500), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n41500), .I0(n11176[19]), .I1(GND_net), 
            .CO(n41501));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n40650), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n11176[18]), .I2(GND_net), 
            .I3(n41499), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22157_2_lut (.I0(n34[5]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4812));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_21 (.CI(n41499), .I0(n11176[18]), .I1(GND_net), 
            .CO(n41500));
    SB_LUT4 add_6782_4_lut (.I0(GND_net), .I1(n20057[1]), .I2(n265), .I3(n40740), 
            .O(n19913[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n11176[17]), .I2(GND_net), 
            .I3(n41498), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6782_4 (.CI(n40740), .I0(n20057[1]), .I1(n265), .CO(n40741));
    SB_CARRY mult_10_add_1225_20 (.CI(n41498), .I0(n11176[17]), .I1(GND_net), 
            .CO(n41499));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n11176[16]), .I2(GND_net), 
            .I3(n41497), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_19 (.CI(n41497), .I0(n11176[16]), .I1(GND_net), 
            .CO(n41498));
    SB_LUT4 i22156_2_lut (.I0(n34[6]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22155_2_lut (.I0(n34[7]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n11176[15]), .I2(GND_net), 
            .I3(n41496), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4817));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_22 (.CI(n40650), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n40651));
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4818));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_18 (.CI(n41496), .I0(n11176[15]), .I1(GND_net), 
            .CO(n41497));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n11176[14]), .I2(GND_net), 
            .I3(n41495), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_12_lut (.I0(GND_net), .I1(n18573[9]), .I2(n831), 
            .I3(n40836), .O(n18153[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6650_12 (.CI(n40836), .I0(n18573[9]), .I1(n831), .CO(n40837));
    SB_CARRY mult_10_add_1225_17 (.CI(n41495), .I0(n11176[14]), .I1(GND_net), 
            .CO(n41496));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n11176[13]), .I2(n1096_adj_4820), 
            .I3(n41494), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n41494), .I0(n11176[13]), .I1(n1096_adj_4820), 
            .CO(n41495));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n11176[12]), .I2(n1023_adj_4821), 
            .I3(n41493), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_15 (.CI(n41493), .I0(n11176[12]), .I1(n1023_adj_4821), 
            .CO(n41494));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n11176[11]), .I2(n950_adj_4822), 
            .I3(n41492), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n41492), .I0(n11176[11]), .I1(n950_adj_4822), 
            .CO(n41493));
    SB_LUT4 add_6650_11_lut (.I0(GND_net), .I1(n18573[8]), .I2(n758), 
            .I3(n40835), .O(n18153[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n11176[10]), .I2(n877_adj_4819), 
            .I3(n41491), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n41491), .I0(n11176[10]), .I1(n877_adj_4819), 
            .CO(n41492));
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n11176[9]), .I2(n804_adj_4818), 
            .I3(n41490), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4821));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_12 (.CI(n41490), .I0(n11176[9]), .I1(n804_adj_4818), 
            .CO(n41491));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n11176[8]), .I2(n731_adj_4817), 
            .I3(n41489), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n41489), .I0(n11176[8]), .I1(n731_adj_4817), 
            .CO(n41490));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n11176[7]), .I2(n658_adj_4816), 
            .I3(n41488), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n41488), .I0(n11176[7]), .I1(n658_adj_4816), 
            .CO(n41489));
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4820));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n11176[6]), .I2(n585_adj_4812), 
            .I3(n41487), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n41487), .I0(n11176[6]), .I1(n585_adj_4812), 
            .CO(n41488));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n11176[5]), .I2(n512_adj_4810), 
            .I3(n41486), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_11 (.CI(n40835), .I0(n18573[8]), .I1(n758), .CO(n40836));
    SB_CARRY mult_10_add_1225_8 (.CI(n41486), .I0(n11176[5]), .I1(n512_adj_4810), 
            .CO(n41487));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n11176[4]), .I2(n439_adj_4796), 
            .I3(n41485), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6782_3_lut (.I0(GND_net), .I1(n20057[0]), .I2(n192), .I3(n40739), 
            .O(n19913[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n41485), .I0(n11176[4]), .I1(n439_adj_4796), 
            .CO(n41486));
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n11176[3]), .I2(n366_adj_4795), 
            .I3(n41484), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_10_lut (.I0(GND_net), .I1(n18573[7]), .I2(n685), 
            .I3(n40834), .O(n18153[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n41484), .I0(n11176[3]), .I1(n366_adj_4795), 
            .CO(n41485));
    SB_CARRY add_6782_3 (.CI(n40739), .I0(n20057[0]), .I1(n192), .CO(n40740));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n11176[2]), .I2(n293_adj_4794), 
            .I3(n41483), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n41483), .I0(n11176[2]), .I1(n293_adj_4794), 
            .CO(n41484));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n11176[1]), .I2(n220_adj_4793), 
            .I3(n41482), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_10 (.CI(n40834), .I0(n18573[7]), .I1(n685), .CO(n40835));
    SB_CARRY mult_10_add_1225_4 (.CI(n41482), .I0(n11176[1]), .I1(n220_adj_4793), 
            .CO(n41483));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n11176[0]), .I2(n147_adj_4792), 
            .I3(n41481), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6782_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n19913[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6782_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6782_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n40739));
    SB_CARRY mult_10_add_1225_3 (.CI(n41481), .I0(n11176[0]), .I1(n147_adj_4792), 
            .CO(n41482));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4791), .I2(n74_adj_4790), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n40649), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4791), .I1(n74_adj_4790), 
            .CO(n41481));
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4809_23_lut (.I0(GND_net), .I1(n13140[20]), .I2(GND_net), 
            .I3(n41480), .O(n11176[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4809_22_lut (.I0(GND_net), .I1(n13140[19]), .I2(GND_net), 
            .I3(n41479), .O(n11176[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n40649), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n40650));
    SB_LUT4 add_957_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4230[23]), .I3(n40578), .O(\PID_CONTROLLER.integral_23__N_3672 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_22 (.CI(n41479), .I0(n13140[19]), .I1(GND_net), 
            .CO(n41480));
    SB_LUT4 add_4809_21_lut (.I0(GND_net), .I1(n13140[18]), .I2(GND_net), 
            .I3(n41478), .O(n11176[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n40648), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_21 (.CI(n41478), .I0(n13140[18]), .I1(GND_net), 
            .CO(n41479));
    SB_LUT4 add_4809_20_lut (.I0(GND_net), .I1(n13140[17]), .I2(GND_net), 
            .I3(n41477), .O(n11176[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22154_2_lut (.I0(n34[8]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22154_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4809_20 (.CI(n41477), .I0(n13140[17]), .I1(GND_net), 
            .CO(n41478));
    SB_LUT4 i22153_2_lut (.I0(n34[9]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4809_19_lut (.I0(GND_net), .I1(n13140[16]), .I2(GND_net), 
            .I3(n41476), .O(n11176[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_19 (.CI(n41476), .I0(n13140[16]), .I1(GND_net), 
            .CO(n41477));
    SB_LUT4 add_4809_18_lut (.I0(GND_net), .I1(n13140[15]), .I2(GND_net), 
            .I3(n41475), .O(n11176[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_18 (.CI(n41475), .I0(n13140[15]), .I1(GND_net), 
            .CO(n41476));
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4809_17_lut (.I0(GND_net), .I1(n13140[14]), .I2(GND_net), 
            .I3(n41474), .O(n11176[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6797_8_lut (.I0(GND_net), .I1(n20169[5]), .I2(n560_adj_4741), 
            .I3(n40738), .O(n20057[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n40648), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n40649));
    SB_CARRY add_4809_17 (.CI(n41474), .I0(n13140[14]), .I1(GND_net), 
            .CO(n41475));
    SB_LUT4 add_4809_16_lut (.I0(GND_net), .I1(n13140[13]), .I2(n1099), 
            .I3(n41473), .O(n11176[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_957_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4230[22]), .I3(n40577), .O(\PID_CONTROLLER.integral_23__N_3672 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_9_lut (.I0(GND_net), .I1(n18573[6]), .I2(n612), .I3(n40833), 
            .O(n18153[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_16 (.CI(n41473), .I0(n13140[13]), .I1(n1099), .CO(n41474));
    SB_LUT4 add_4809_15_lut (.I0(GND_net), .I1(n13140[12]), .I2(n1026), 
            .I3(n41472), .O(n11176[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22152_2_lut (.I0(n34[10]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22152_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4809_15 (.CI(n41472), .I0(n13140[12]), .I1(n1026), .CO(n41473));
    SB_LUT4 add_4809_14_lut (.I0(GND_net), .I1(n13140[11]), .I2(n953), 
            .I3(n41471), .O(n11176[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_9 (.CI(n40833), .I0(n18573[6]), .I1(n612), .CO(n40834));
    SB_CARRY add_4809_14 (.CI(n41471), .I0(n13140[11]), .I1(n953), .CO(n41472));
    SB_LUT4 add_4809_13_lut (.I0(GND_net), .I1(n13140[10]), .I2(n880), 
            .I3(n41470), .O(n11176[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_13 (.CI(n41470), .I0(n13140[10]), .I1(n880), .CO(n41471));
    SB_LUT4 add_4809_12_lut (.I0(GND_net), .I1(n13140[9]), .I2(n807), 
            .I3(n41469), .O(n11176[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6797_7_lut (.I0(GND_net), .I1(n20169[4]), .I2(n487_adj_4739), 
            .I3(n40737), .O(n20057[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_12 (.CI(n41469), .I0(n13140[9]), .I1(n807), .CO(n41470));
    SB_LUT4 add_4809_11_lut (.I0(GND_net), .I1(n13140[8]), .I2(n734), 
            .I3(n41468), .O(n11176[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_11 (.CI(n41468), .I0(n13140[8]), .I1(n734), .CO(n41469));
    SB_LUT4 add_4809_10_lut (.I0(GND_net), .I1(n13140[7]), .I2(n661), 
            .I3(n41467), .O(n11176[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_10 (.CI(n41467), .I0(n13140[7]), .I1(n661), .CO(n41468));
    SB_LUT4 add_4809_9_lut (.I0(GND_net), .I1(n13140[6]), .I2(n588), .I3(n41466), 
            .O(n11176[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n40647), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6797_7 (.CI(n40737), .I0(n20169[4]), .I1(n487_adj_4739), 
            .CO(n40738));
    SB_CARRY add_4809_9 (.CI(n41466), .I0(n13140[6]), .I1(n588), .CO(n41467));
    SB_LUT4 add_4809_8_lut (.I0(GND_net), .I1(n13140[5]), .I2(n515), .I3(n41465), 
            .O(n11176[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_8 (.CI(n41465), .I0(n13140[5]), .I1(n515), .CO(n41466));
    SB_LUT4 add_6650_8_lut (.I0(GND_net), .I1(n18573[5]), .I2(n539), .I3(n40832), 
            .O(n18153[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4809_7_lut (.I0(GND_net), .I1(n13140[4]), .I2(n442), .I3(n41464), 
            .O(n11176[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_7 (.CI(n41464), .I0(n13140[4]), .I1(n442), .CO(n41465));
    SB_LUT4 add_4809_6_lut (.I0(GND_net), .I1(n13140[3]), .I2(n369), .I3(n41463), 
            .O(n11176[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4830));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4832));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4833));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4835));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4836));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22151_2_lut (.I0(n34[11]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4809_6 (.CI(n41463), .I0(n13140[3]), .I1(n369), .CO(n41464));
    SB_CARRY sub_3_add_2_19 (.CI(n40647), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n40648));
    SB_LUT4 add_4809_5_lut (.I0(GND_net), .I1(n13140[2]), .I2(n296), .I3(n41462), 
            .O(n11176[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_5 (.CI(n41462), .I0(n13140[2]), .I1(n296), .CO(n41463));
    SB_LUT4 add_4809_4_lut (.I0(GND_net), .I1(n13140[1]), .I2(n223), .I3(n41461), 
            .O(n11176[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_4 (.CI(n41461), .I0(n13140[1]), .I1(n223), .CO(n41462));
    SB_LUT4 add_4809_3_lut (.I0(GND_net), .I1(n13140[0]), .I2(n150), .I3(n41460), 
            .O(n11176[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_3 (.CI(n41460), .I0(n13140[0]), .I1(n150), .CO(n41461));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n40646), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4809_2_lut (.I0(GND_net), .I1(n8_adj_4738), .I2(n77), 
            .I3(GND_net), .O(n11176[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4809_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4809_2 (.CI(GND_net), .I0(n8_adj_4738), .I1(n77), .CO(n41460));
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4838));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4839));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6650_8 (.CI(n40832), .I0(n18573[5]), .I1(n539), .CO(n40833));
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_957_24 (.CI(n40577), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4230[22]), .CO(n40578));
    SB_CARRY sub_3_add_2_18 (.CI(n40646), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n40647));
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n40645), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6650_7_lut (.I0(GND_net), .I1(n18573[4]), .I2(n466), .I3(n40831), 
            .O(n18153[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_7 (.CI(n40831), .I0(n18573[4]), .I1(n466), .CO(n40832));
    SB_LUT4 add_6650_6_lut (.I0(GND_net), .I1(n18573[3]), .I2(n393), .I3(n40830), 
            .O(n18153[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6797_6_lut (.I0(GND_net), .I1(n20169[3]), .I2(n414_adj_4737), 
            .I3(n40736), .O(n20057[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6797_6 (.CI(n40736), .I0(n20169[3]), .I1(n414_adj_4737), 
            .CO(n40737));
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4842));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6650_6 (.CI(n40830), .I0(n18573[3]), .I1(n393), .CO(n40831));
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4843));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4844));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6650_5_lut (.I0(GND_net), .I1(n18573[2]), .I2(n320), .I3(n40829), 
            .O(n18153[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6797_5_lut (.I0(GND_net), .I1(n20169[2]), .I2(n341), .I3(n40735), 
            .O(n20057[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n40645), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n40646));
    SB_CARRY add_6797_5 (.CI(n40735), .I0(n20169[2]), .I1(n341), .CO(n40736));
    SB_LUT4 add_957_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4230[21]), .I3(n40576), .O(\PID_CONTROLLER.integral_23__N_3672 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_5 (.CI(n40829), .I0(n18573[2]), .I1(n320), .CO(n40830));
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6650_4_lut (.I0(GND_net), .I1(n18573[1]), .I2(n247), .I3(n40828), 
            .O(n18153[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_4 (.CI(n40828), .I0(n18573[1]), .I1(n247), .CO(n40829));
    SB_LUT4 add_6650_3_lut (.I0(GND_net), .I1(n18573[0]), .I2(n174), .I3(n40827), 
            .O(n18153[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6650_3 (.CI(n40827), .I0(n18573[0]), .I1(n174), .CO(n40828));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n40644), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6797_4_lut (.I0(GND_net), .I1(n20169[1]), .I2(n268), .I3(n40734), 
            .O(n20057[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_23 (.CI(n40576), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4230[21]), .CO(n40577));
    SB_CARRY sub_3_add_2_16 (.CI(n40644), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n40645));
    SB_LUT4 add_6650_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18153[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6650_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6650_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n40827));
    SB_CARRY add_6797_4 (.CI(n40734), .I0(n20169[1]), .I1(n268), .CO(n40735));
    SB_LUT4 add_6797_3_lut (.I0(GND_net), .I1(n20169[0]), .I2(n195), .I3(n40733), 
            .O(n20057[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n40643), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6804_8_lut (.I0(GND_net), .I1(n20217[5]), .I2(n560), .I3(n40826), 
            .O(n20120[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n40643), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n40644));
    SB_LUT4 add_957_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4230[20]), .I3(n40575), .O(\PID_CONTROLLER.integral_23__N_3672 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4808));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6804_7_lut (.I0(GND_net), .I1(n20217[4]), .I2(n487), .I3(n40825), 
            .O(n20120[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5774_22_lut (.I0(GND_net), .I1(n14671[19]), .I2(GND_net), 
            .I3(n41436), .O(n13140[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5774_21_lut (.I0(GND_net), .I1(n14671[18]), .I2(GND_net), 
            .I3(n41435), .O(n13140[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6804_7 (.CI(n40825), .I0(n20217[4]), .I1(n487), .CO(n40826));
    SB_CARRY add_5774_21 (.CI(n41435), .I0(n14671[18]), .I1(GND_net), 
            .CO(n41436));
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5774_20_lut (.I0(GND_net), .I1(n14671[17]), .I2(GND_net), 
            .I3(n41434), .O(n13140[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_20 (.CI(n41434), .I0(n14671[17]), .I1(GND_net), 
            .CO(n41435));
    SB_LUT4 add_5774_19_lut (.I0(GND_net), .I1(n14671[16]), .I2(GND_net), 
            .I3(n41433), .O(n13140[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_19 (.CI(n41433), .I0(n14671[16]), .I1(GND_net), 
            .CO(n41434));
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5774_18_lut (.I0(GND_net), .I1(n14671[15]), .I2(GND_net), 
            .I3(n41432), .O(n13140[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_18 (.CI(n41432), .I0(n14671[15]), .I1(GND_net), 
            .CO(n41433));
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5774_17_lut (.I0(GND_net), .I1(n14671[14]), .I2(GND_net), 
            .I3(n41431), .O(n13140[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6797_3 (.CI(n40733), .I0(n20169[0]), .I1(n195), .CO(n40734));
    SB_CARRY add_5774_17 (.CI(n41431), .I0(n14671[14]), .I1(GND_net), 
            .CO(n41432));
    SB_LUT4 add_5774_16_lut (.I0(GND_net), .I1(n14671[13]), .I2(n1102), 
            .I3(n41430), .O(n13140[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_16 (.CI(n41430), .I0(n14671[13]), .I1(n1102), .CO(n41431));
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5774_15_lut (.I0(GND_net), .I1(n14671[12]), .I2(n1029), 
            .I3(n41429), .O(n13140[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_15 (.CI(n41429), .I0(n14671[12]), .I1(n1029), .CO(n41430));
    SB_LUT4 add_5774_14_lut (.I0(GND_net), .I1(n14671[11]), .I2(n956), 
            .I3(n41428), .O(n13140[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_14 (.CI(n41428), .I0(n14671[11]), .I1(n956), .CO(n41429));
    SB_LUT4 add_5774_13_lut (.I0(GND_net), .I1(n14671[10]), .I2(n883), 
            .I3(n41427), .O(n13140[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_13 (.CI(n41427), .I0(n14671[10]), .I1(n883), .CO(n41428));
    SB_LUT4 add_5774_12_lut (.I0(GND_net), .I1(n14671[9]), .I2(n810), 
            .I3(n41426), .O(n13140[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_12 (.CI(n41426), .I0(n14671[9]), .I1(n810), .CO(n41427));
    SB_LUT4 add_5774_11_lut (.I0(GND_net), .I1(n14671[8]), .I2(n737), 
            .I3(n41425), .O(n13140[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_11 (.CI(n41425), .I0(n14671[8]), .I1(n737), .CO(n41426));
    SB_LUT4 add_5774_10_lut (.I0(GND_net), .I1(n14671[7]), .I2(n664), 
            .I3(n41424), .O(n13140[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_10 (.CI(n41424), .I0(n14671[7]), .I1(n664), .CO(n41425));
    SB_LUT4 add_5774_9_lut (.I0(GND_net), .I1(n14671[6]), .I2(n591), .I3(n41423), 
            .O(n13140[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_9 (.CI(n41423), .I0(n14671[6]), .I1(n591), .CO(n41424));
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5774_8_lut (.I0(GND_net), .I1(n14671[5]), .I2(n518), .I3(n41422), 
            .O(n13140[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_8 (.CI(n41422), .I0(n14671[5]), .I1(n518), .CO(n41423));
    SB_LUT4 add_5774_7_lut (.I0(GND_net), .I1(n14671[4]), .I2(n445), .I3(n41421), 
            .O(n13140[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6797_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20057[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6797_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_7 (.CI(n41421), .I0(n14671[4]), .I1(n445), .CO(n41422));
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5774_6_lut (.I0(GND_net), .I1(n14671[3]), .I2(n372), .I3(n41420), 
            .O(n13140[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5774_6 (.CI(n41420), .I0(n14671[3]), .I1(n372), .CO(n41421));
    SB_LUT4 add_5774_5_lut (.I0(GND_net), .I1(n14671[2]), .I2(n299), .I3(n41419), 
            .O(n13140[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4848));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4849));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5774_5 (.CI(n41419), .I0(n14671[2]), .I1(n299), .CO(n41420));
    SB_LUT4 add_5774_4_lut (.I0(GND_net), .I1(n14671[1]), .I2(n226), .I3(n41418), 
            .O(n13140[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_4 (.CI(n41418), .I0(n14671[1]), .I1(n226), .CO(n41419));
    SB_LUT4 add_5774_3_lut (.I0(GND_net), .I1(n14671[0]), .I2(n153), .I3(n41417), 
            .O(n13140[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5774_3 (.CI(n41417), .I0(n14671[0]), .I1(n153), .CO(n41418));
    SB_LUT4 add_5774_2_lut (.I0(GND_net), .I1(n11_adj_4733), .I2(n80), 
            .I3(GND_net), .O(n13140[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5774_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5774_2 (.CI(GND_net), .I0(n11_adj_4733), .I1(n80), .CO(n41417));
    SB_CARRY add_6797_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n40733));
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n40642), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6464_21_lut (.I0(GND_net), .I1(n15472[18]), .I2(GND_net), 
            .I3(n41416), .O(n14671[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_22 (.CI(n40575), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4230[20]), .CO(n40576));
    SB_LUT4 add_6464_20_lut (.I0(GND_net), .I1(n15472[17]), .I2(GND_net), 
            .I3(n41415), .O(n14671[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_20 (.CI(n41415), .I0(n15472[17]), .I1(GND_net), 
            .CO(n41416));
    SB_LUT4 add_6464_19_lut (.I0(GND_net), .I1(n15472[16]), .I2(GND_net), 
            .I3(n41414), .O(n14671[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6804_6_lut (.I0(GND_net), .I1(n20217[3]), .I2(n414), .I3(n40824), 
            .O(n20120[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_19 (.CI(n41414), .I0(n15472[16]), .I1(GND_net), 
            .CO(n41415));
    SB_LUT4 add_6464_18_lut (.I0(GND_net), .I1(n15472[15]), .I2(GND_net), 
            .I3(n41413), .O(n14671[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_18 (.CI(n41413), .I0(n15472[15]), .I1(GND_net), 
            .CO(n41414));
    SB_LUT4 add_6464_17_lut (.I0(GND_net), .I1(n15472[14]), .I2(GND_net), 
            .I3(n41412), .O(n14671[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6804_6 (.CI(n40824), .I0(n20217[3]), .I1(n414), .CO(n40825));
    SB_CARRY add_6464_17 (.CI(n41412), .I0(n15472[14]), .I1(GND_net), 
            .CO(n41413));
    SB_LUT4 add_6810_7_lut (.I0(GND_net), .I1(n47913), .I2(n490), .I3(n40732), 
            .O(n20169[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n40642), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n40643));
    SB_LUT4 add_6464_16_lut (.I0(GND_net), .I1(n15472[13]), .I2(n1105), 
            .I3(n41411), .O(n14671[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6810_6_lut (.I0(GND_net), .I1(n20253[3]), .I2(n417_adj_4852), 
            .I3(n40731), .O(n20169[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_16 (.CI(n41411), .I0(n15472[13]), .I1(n1105), .CO(n41412));
    SB_LUT4 add_6804_5_lut (.I0(GND_net), .I1(n20217[2]), .I2(n341_adj_4853), 
            .I3(n40823), .O(n20120[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6464_15_lut (.I0(GND_net), .I1(n15472[12]), .I2(n1032), 
            .I3(n41410), .O(n14671[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4854));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6464_15 (.CI(n41410), .I0(n15472[12]), .I1(n1032), .CO(n41411));
    SB_CARRY add_6804_5 (.CI(n40823), .I0(n20217[2]), .I1(n341_adj_4853), 
            .CO(n40824));
    SB_LUT4 add_6804_4_lut (.I0(GND_net), .I1(n20217[1]), .I2(n268_adj_4855), 
            .I3(n40822), .O(n20120[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6464_14_lut (.I0(GND_net), .I1(n15472[11]), .I2(n959), 
            .I3(n41409), .O(n14671[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_14 (.CI(n41409), .I0(n15472[11]), .I1(n959), .CO(n41410));
    SB_LUT4 add_957_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4230[19]), .I3(n40574), .O(\PID_CONTROLLER.integral_23__N_3672 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6464_13_lut (.I0(GND_net), .I1(n15472[10]), .I2(n886), 
            .I3(n41408), .O(n14671[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_13 (.CI(n41408), .I0(n15472[10]), .I1(n886), .CO(n41409));
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4856));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4858));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4859));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4860));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4862));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_12_lut (.I0(GND_net), .I1(n15472[9]), .I2(n813), 
            .I3(n41407), .O(n14671[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_21 (.CI(n40574), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4230[19]), .CO(n40575));
    SB_CARRY add_6464_12 (.CI(n41407), .I0(n15472[9]), .I1(n813), .CO(n41408));
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4863));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_11_lut (.I0(GND_net), .I1(n15472[8]), .I2(n740), 
            .I3(n41406), .O(n14671[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_11 (.CI(n41406), .I0(n15472[8]), .I1(n740), .CO(n41407));
    SB_LUT4 add_6464_10_lut (.I0(GND_net), .I1(n15472[7]), .I2(n667), 
            .I3(n41405), .O(n14671[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_10 (.CI(n41405), .I0(n15472[7]), .I1(n667), .CO(n41406));
    SB_CARRY add_6810_6 (.CI(n40731), .I0(n20253[3]), .I1(n417_adj_4852), 
            .CO(n40732));
    SB_LUT4 add_6810_5_lut (.I0(GND_net), .I1(n20253[2]), .I2(n344_adj_4864), 
            .I3(n40730), .O(n20169[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_9_lut (.I0(GND_net), .I1(n15472[6]), .I2(n594), .I3(n41404), 
            .O(n14671[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_9 (.CI(n41404), .I0(n15472[6]), .I1(n594), .CO(n41405));
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4865));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_8_lut (.I0(GND_net), .I1(n15472[5]), .I2(n521), .I3(n41403), 
            .O(n14671[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6464_8 (.CI(n41403), .I0(n15472[5]), .I1(n521), .CO(n41404));
    SB_LUT4 add_6464_7_lut (.I0(GND_net), .I1(n15472[4]), .I2(n448), .I3(n41402), 
            .O(n14671[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_7 (.CI(n41402), .I0(n15472[4]), .I1(n448), .CO(n41403));
    SB_LUT4 add_6464_6_lut (.I0(GND_net), .I1(n15472[3]), .I2(n375), .I3(n41401), 
            .O(n14671[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_6 (.CI(n41401), .I0(n15472[3]), .I1(n375), .CO(n41402));
    SB_LUT4 add_6464_5_lut (.I0(GND_net), .I1(n15472[2]), .I2(n302), .I3(n41400), 
            .O(n14671[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6810_5 (.CI(n40730), .I0(n20253[2]), .I1(n344_adj_4864), 
            .CO(n40731));
    SB_LUT4 add_957_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4230[18]), .I3(n40573), .O(\PID_CONTROLLER.integral_23__N_3672 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_5 (.CI(n41400), .I0(n15472[2]), .I1(n302), .CO(n41401));
    SB_LUT4 add_6464_4_lut (.I0(GND_net), .I1(n15472[1]), .I2(n229), .I3(n41399), 
            .O(n14671[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6810_4_lut (.I0(GND_net), .I1(n20253[1]), .I2(n271_adj_4866), 
            .I3(n40729), .O(n20169[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_4 (.CI(n41399), .I0(n15472[1]), .I1(n229), .CO(n41400));
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_3_lut (.I0(GND_net), .I1(n15472[0]), .I2(n156), .I3(n41398), 
            .O(n14671[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6464_3 (.CI(n41398), .I0(n15472[0]), .I1(n156), .CO(n41399));
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6464_2_lut (.I0(GND_net), .I1(n14_adj_4867), .I2(n83), 
            .I3(GND_net), .O(n14671[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6464_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6464_2 (.CI(GND_net), .I0(n14_adj_4867), .I1(n83), .CO(n41398));
    SB_LUT4 add_6504_20_lut (.I0(GND_net), .I1(n16193[17]), .I2(GND_net), 
            .I3(n41397), .O(n15472[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6504_19_lut (.I0(GND_net), .I1(n16193[16]), .I2(GND_net), 
            .I3(n41396), .O(n15472[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n40641), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_19 (.CI(n41396), .I0(n16193[16]), .I1(GND_net), 
            .CO(n41397));
    SB_LUT4 add_6504_18_lut (.I0(GND_net), .I1(n16193[15]), .I2(GND_net), 
            .I3(n41395), .O(n15472[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_18 (.CI(n41395), .I0(n16193[15]), .I1(GND_net), 
            .CO(n41396));
    SB_CARRY add_957_20 (.CI(n40573), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4230[18]), .CO(n40574));
    SB_LUT4 add_6504_17_lut (.I0(GND_net), .I1(n16193[14]), .I2(GND_net), 
            .I3(n41394), .O(n15472[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_17 (.CI(n41394), .I0(n16193[14]), .I1(GND_net), 
            .CO(n41395));
    SB_LUT4 add_6504_16_lut (.I0(GND_net), .I1(n16193[13]), .I2(n1108), 
            .I3(n41393), .O(n15472[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n40641), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n40642));
    SB_LUT4 add_957_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4230[17]), .I3(n40572), .O(\PID_CONTROLLER.integral_23__N_3672 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_16 (.CI(n41393), .I0(n16193[13]), .I1(n1108), .CO(n41394));
    SB_CARRY add_6804_4 (.CI(n40822), .I0(n20217[1]), .I1(n268_adj_4855), 
            .CO(n40823));
    SB_LUT4 add_6504_15_lut (.I0(GND_net), .I1(n16193[12]), .I2(n1035), 
            .I3(n41392), .O(n15472[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_15 (.CI(n41392), .I0(n16193[12]), .I1(n1035), .CO(n41393));
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n40640), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6504_14_lut (.I0(GND_net), .I1(n16193[11]), .I2(n962), 
            .I3(n41391), .O(n15472[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_14 (.CI(n41391), .I0(n16193[11]), .I1(n962), .CO(n41392));
    SB_CARRY add_6810_4 (.CI(n40729), .I0(n20253[1]), .I1(n271_adj_4866), 
            .CO(n40730));
    SB_LUT4 add_6504_13_lut (.I0(GND_net), .I1(n16193[10]), .I2(n889), 
            .I3(n41390), .O(n15472[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_19 (.CI(n40572), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4230[17]), .CO(n40573));
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_13 (.CI(n41390), .I0(n16193[10]), .I1(n889), .CO(n41391));
    SB_LUT4 add_6504_12_lut (.I0(GND_net), .I1(n16193[9]), .I2(n816), 
            .I3(n41389), .O(n15472[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_12 (.CI(n41389), .I0(n16193[9]), .I1(n816), .CO(n41390));
    SB_LUT4 add_6504_11_lut (.I0(GND_net), .I1(n16193[8]), .I2(n743), 
            .I3(n41388), .O(n15472[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_11 (.CI(n41388), .I0(n16193[8]), .I1(n743), .CO(n41389));
    SB_LUT4 add_6504_10_lut (.I0(GND_net), .I1(n16193[7]), .I2(n670), 
            .I3(n41387), .O(n15472[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_10 (.CI(n41387), .I0(n16193[7]), .I1(n670), .CO(n41388));
    SB_LUT4 add_6504_9_lut (.I0(GND_net), .I1(n16193[6]), .I2(n597), .I3(n41386), 
            .O(n15472[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_9 (.CI(n41386), .I0(n16193[6]), .I1(n597), .CO(n41387));
    SB_LUT4 add_6504_8_lut (.I0(GND_net), .I1(n16193[5]), .I2(n524), .I3(n41385), 
            .O(n15472[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_8 (.CI(n41385), .I0(n16193[5]), .I1(n524), .CO(n41386));
    SB_LUT4 add_6504_7_lut (.I0(GND_net), .I1(n16193[4]), .I2(n451), .I3(n41384), 
            .O(n15472[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_7 (.CI(n41384), .I0(n16193[4]), .I1(n451), .CO(n41385));
    SB_LUT4 add_6504_6_lut (.I0(GND_net), .I1(n16193[3]), .I2(n378), .I3(n41383), 
            .O(n15472[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_6 (.CI(n41383), .I0(n16193[3]), .I1(n378), .CO(n41384));
    SB_LUT4 add_6504_5_lut (.I0(GND_net), .I1(n16193[2]), .I2(n305), .I3(n41382), 
            .O(n15472[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_5 (.CI(n41382), .I0(n16193[2]), .I1(n305), .CO(n41383));
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4869));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6504_4_lut (.I0(GND_net), .I1(n16193[1]), .I2(n232), .I3(n41381), 
            .O(n15472[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_4 (.CI(n41381), .I0(n16193[1]), .I1(n232), .CO(n41382));
    SB_LUT4 add_6504_3_lut (.I0(GND_net), .I1(n16193[0]), .I2(n159), .I3(n41380), 
            .O(n15472[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6804_3_lut (.I0(GND_net), .I1(n20217[0]), .I2(n195_adj_4871), 
            .I3(n40821), .O(n20120[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6504_3 (.CI(n41380), .I0(n16193[0]), .I1(n159), .CO(n41381));
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6504_2_lut (.I0(GND_net), .I1(n17_adj_4872), .I2(n86), 
            .I3(GND_net), .O(n15472[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6504_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6504_2 (.CI(GND_net), .I0(n17_adj_4872), .I1(n86), .CO(n41380));
    SB_LUT4 add_6540_19_lut (.I0(GND_net), .I1(n16840[16]), .I2(GND_net), 
            .I3(n41379), .O(n16193[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6810_3_lut (.I0(GND_net), .I1(n20253[0]), .I2(n198_adj_4873), 
            .I3(n40728), .O(n20169[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_6540_18_lut (.I0(GND_net), .I1(n16840[15]), .I2(GND_net), 
            .I3(n41378), .O(n16193[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_957_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4230[16]), .I3(n40571), .O(\PID_CONTROLLER.integral_23__N_3672 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_18 (.CI(n41378), .I0(n16840[15]), .I1(GND_net), 
            .CO(n41379));
    SB_LUT4 add_6540_17_lut (.I0(GND_net), .I1(n16840[14]), .I2(GND_net), 
            .I3(n41377), .O(n16193[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6810_3 (.CI(n40728), .I0(n20253[0]), .I1(n198_adj_4873), 
            .CO(n40729));
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6540_17 (.CI(n41377), .I0(n16840[14]), .I1(GND_net), 
            .CO(n41378));
    SB_CARRY sub_3_add_2_12 (.CI(n40640), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n40641));
    SB_CARRY add_6804_3 (.CI(n40821), .I0(n20217[0]), .I1(n195_adj_4871), 
            .CO(n40822));
    SB_LUT4 add_6540_16_lut (.I0(GND_net), .I1(n16840[13]), .I2(n1111), 
            .I3(n41376), .O(n16193[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_16 (.CI(n41376), .I0(n16840[13]), .I1(n1111), .CO(n41377));
    SB_LUT4 add_6540_15_lut (.I0(GND_net), .I1(n16840[12]), .I2(n1038), 
            .I3(n41375), .O(n16193[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_6540_15 (.CI(n41375), .I0(n16840[12]), .I1(n1038), .CO(n41376));
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_6540_14_lut (.I0(GND_net), .I1(n16840[11]), .I2(n965), 
            .I3(n41374), .O(n16193[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_6540_14 (.CI(n41374), .I0(n16840[11]), .I1(n965), .CO(n41375));
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_6540_13_lut (.I0(GND_net), .I1(n16840[10]), .I2(n892), 
            .I3(n41373), .O(n16193[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_6540_13 (.CI(n41373), .I0(n16840[10]), .I1(n892), .CO(n41374));
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3648[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3648[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3648[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3648[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3648[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3648[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3648[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3648[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3648[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3648[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3648[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_6540_12_lut (.I0(GND_net), .I1(n16840[9]), .I2(n819), 
            .I3(n41372), .O(n16193[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3648[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3648[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3648[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6540_12 (.CI(n41372), .I0(n16840[9]), .I1(n819), .CO(n41373));
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_11_lut (.I0(GND_net), .I1(n16840[8]), .I2(n746), 
            .I3(n41371), .O(n16193[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3648[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_6540_11 (.CI(n41371), .I0(n16840[8]), .I1(n746), .CO(n41372));
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3648[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3648[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3648[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3648[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3648[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3648[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3648[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3648[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4876));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_10_lut (.I0(GND_net), .I1(n16840[7]), .I2(n673), 
            .I3(n41370), .O(n16193[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_10 (.CI(n41370), .I0(n16840[7]), .I1(n673), .CO(n41371));
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_9_lut (.I0(GND_net), .I1(n16840[6]), .I2(n600), .I3(n41369), 
            .O(n16193[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4878));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6540_9 (.CI(n41369), .I0(n16840[6]), .I1(n600), .CO(n41370));
    SB_LUT4 add_6540_8_lut (.I0(GND_net), .I1(n16840[5]), .I2(n527), .I3(n41368), 
            .O(n16193[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6540_8 (.CI(n41368), .I0(n16840[5]), .I1(n527), .CO(n41369));
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4881));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_7_lut (.I0(GND_net), .I1(n16840[4]), .I2(n454), .I3(n41367), 
            .O(n16193[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_7 (.CI(n41367), .I0(n16840[4]), .I1(n454), .CO(n41368));
    SB_LUT4 add_6540_6_lut (.I0(GND_net), .I1(n16840[3]), .I2(n381), .I3(n41366), 
            .O(n16193[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_6 (.CI(n41366), .I0(n16840[3]), .I1(n381), .CO(n41367));
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4882));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_5_lut (.I0(GND_net), .I1(n16840[2]), .I2(n308), .I3(n41365), 
            .O(n16193[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n40639), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_5 (.CI(n41365), .I0(n16840[2]), .I1(n308), .CO(n41366));
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_4_lut (.I0(GND_net), .I1(n16840[1]), .I2(n235), .I3(n41364), 
            .O(n16193[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6540_4 (.CI(n41364), .I0(n16840[1]), .I1(n235), .CO(n41365));
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4884));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6540_3_lut (.I0(GND_net), .I1(n16840[0]), .I2(n162), .I3(n41363), 
            .O(n16193[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4885));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6810_2_lut (.I0(GND_net), .I1(n56_adj_4886), .I2(n125_adj_4887), 
            .I3(GND_net), .O(n20169[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6810_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6810_2 (.CI(GND_net), .I0(n56_adj_4886), .I1(n125_adj_4887), 
            .CO(n40728));
    SB_LUT4 add_6804_2_lut (.I0(GND_net), .I1(n53_adj_4888), .I2(n122_adj_4889), 
            .I3(GND_net), .O(n20120[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6804_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4890));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6540_3 (.CI(n41363), .I0(n16840[0]), .I1(n162), .CO(n41364));
    SB_CARRY add_6804_2 (.CI(GND_net), .I0(n53_adj_4888), .I1(n122_adj_4889), 
            .CO(n40821));
    SB_LUT4 add_6540_2_lut (.I0(GND_net), .I1(n20_adj_4891), .I2(n89), 
            .I3(GND_net), .O(n16193[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6540_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6540_2 (.CI(GND_net), .I0(n20_adj_4891), .I1(n89), .CO(n41363));
    SB_LUT4 add_6574_18_lut (.I0(GND_net), .I1(n17417[15]), .I2(GND_net), 
            .I3(n41362), .O(n16840[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n40639), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n40640));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n40638), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6574_17_lut (.I0(GND_net), .I1(n17417[14]), .I2(GND_net), 
            .I3(n41361), .O(n16840[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_17 (.CI(n41361), .I0(n17417[14]), .I1(GND_net), 
            .CO(n41362));
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4893));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4894));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6574_16_lut (.I0(GND_net), .I1(n17417[13]), .I2(n1114_adj_4895), 
            .I3(n41360), .O(n16840[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_16 (.CI(n41360), .I0(n17417[13]), .I1(n1114_adj_4895), 
            .CO(n41361));
    SB_LUT4 add_6574_15_lut (.I0(GND_net), .I1(n17417[12]), .I2(n1041_adj_4896), 
            .I3(n41359), .O(n16840[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_15 (.CI(n41359), .I0(n17417[12]), .I1(n1041_adj_4896), 
            .CO(n41360));
    SB_LUT4 add_6574_14_lut (.I0(GND_net), .I1(n17417[11]), .I2(n968_adj_4897), 
            .I3(n41358), .O(n16840[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_14 (.CI(n41358), .I0(n17417[11]), .I1(n968_adj_4897), 
            .CO(n41359));
    SB_LUT4 add_6574_13_lut (.I0(GND_net), .I1(n17417[10]), .I2(n895_adj_4898), 
            .I3(n41357), .O(n16840[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_13 (.CI(n41357), .I0(n17417[10]), .I1(n895_adj_4898), 
            .CO(n41358));
    SB_LUT4 add_6574_12_lut (.I0(GND_net), .I1(n17417[9]), .I2(n822_adj_4899), 
            .I3(n41356), .O(n16840[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4900));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6574_12 (.CI(n41356), .I0(n17417[9]), .I1(n822_adj_4899), 
            .CO(n41357));
    SB_LUT4 add_6574_11_lut (.I0(GND_net), .I1(n17417[8]), .I2(n749_adj_4901), 
            .I3(n41355), .O(n16840[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_11 (.CI(n41355), .I0(n17417[8]), .I1(n749_adj_4901), 
            .CO(n41356));
    SB_LUT4 add_6574_10_lut (.I0(GND_net), .I1(n17417[7]), .I2(n676_adj_4902), 
            .I3(n41354), .O(n16840[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_10 (.CI(n41354), .I0(n17417[7]), .I1(n676_adj_4902), 
            .CO(n41355));
    SB_LUT4 add_6574_9_lut (.I0(GND_net), .I1(n17417[6]), .I2(n603_adj_4903), 
            .I3(n41353), .O(n16840[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_9 (.CI(n41353), .I0(n17417[6]), .I1(n603_adj_4903), 
            .CO(n41354));
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6574_8_lut (.I0(GND_net), .I1(n17417[5]), .I2(n530_adj_4905), 
            .I3(n41352), .O(n16840[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_8 (.CI(n41352), .I0(n17417[5]), .I1(n530_adj_4905), 
            .CO(n41353));
    SB_LUT4 add_6574_7_lut (.I0(GND_net), .I1(n17417[4]), .I2(n457_adj_4906), 
            .I3(n41351), .O(n16840[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4908));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6574_7 (.CI(n41351), .I0(n17417[4]), .I1(n457_adj_4906), 
            .CO(n41352));
    SB_LUT4 add_6574_6_lut (.I0(GND_net), .I1(n17417[3]), .I2(n384_adj_4909), 
            .I3(n41350), .O(n16840[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_6 (.CI(n41350), .I0(n17417[3]), .I1(n384_adj_4909), 
            .CO(n41351));
    SB_LUT4 add_6574_5_lut (.I0(GND_net), .I1(n17417[2]), .I2(n311_adj_4910), 
            .I3(n41349), .O(n16840[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n40638), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n40639));
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_957_18 (.CI(n40571), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4230[16]), .CO(n40572));
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4912));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4913));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6574_5 (.CI(n41349), .I0(n17417[2]), .I1(n311_adj_4910), 
            .CO(n41350));
    SB_LUT4 add_6574_4_lut (.I0(GND_net), .I1(n17417[1]), .I2(n238_adj_4914), 
            .I3(n41348), .O(n16840[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_4 (.CI(n41348), .I0(n17417[1]), .I1(n238_adj_4914), 
            .CO(n41349));
    SB_LUT4 add_6574_3_lut (.I0(GND_net), .I1(n17417[0]), .I2(n165_adj_4915), 
            .I3(n41347), .O(n16840[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6574_3 (.CI(n41347), .I0(n17417[0]), .I1(n165_adj_4915), 
            .CO(n41348));
    SB_LUT4 add_6574_2_lut (.I0(GND_net), .I1(n23_adj_4916), .I2(n92_adj_4917), 
            .I3(GND_net), .O(n16840[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6574_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n40637), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6574_2 (.CI(GND_net), .I0(n23_adj_4916), .I1(n92_adj_4917), 
            .CO(n41347));
    SB_CARRY sub_3_add_2_9 (.CI(n40637), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n40638));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n40636), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6606_17_lut (.I0(GND_net), .I1(n17928[14]), .I2(GND_net), 
            .I3(n41346), .O(n17417[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_957_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4230[15]), .I3(n40570), .O(\PID_CONTROLLER.integral_23__N_3672 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n40636), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n40637));
    SB_LUT4 add_6606_16_lut (.I0(GND_net), .I1(n17928[13]), .I2(n1117_adj_4918), 
            .I3(n41345), .O(n17417[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n40635), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n40635), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n40636));
    SB_CARRY add_6606_16 (.CI(n41345), .I0(n17928[13]), .I1(n1117_adj_4918), 
            .CO(n41346));
    SB_LUT4 add_6606_15_lut (.I0(GND_net), .I1(n17928[12]), .I2(n1044_adj_4919), 
            .I3(n41344), .O(n17417[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_15 (.CI(n41344), .I0(n17928[12]), .I1(n1044_adj_4919), 
            .CO(n41345));
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4920));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4921));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6606_14_lut (.I0(GND_net), .I1(n17928[11]), .I2(n971_adj_4922), 
            .I3(n41343), .O(n17417[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_14 (.CI(n41343), .I0(n17928[11]), .I1(n971_adj_4922), 
            .CO(n41344));
    SB_LUT4 add_6606_13_lut (.I0(GND_net), .I1(n17928[10]), .I2(n898_adj_4923), 
            .I3(n41342), .O(n17417[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_13 (.CI(n41342), .I0(n17928[10]), .I1(n898_adj_4923), 
            .CO(n41343));
    SB_LUT4 add_6606_12_lut (.I0(GND_net), .I1(n17928[9]), .I2(n825_adj_4924), 
            .I3(n41341), .O(n17417[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n40634), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4925));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4926));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6606_12 (.CI(n41341), .I0(n17928[9]), .I1(n825_adj_4924), 
            .CO(n41342));
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4929));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4930));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4931));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4932));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4933));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4934));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4936));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3772[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4937));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3772[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4938));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4939));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3772[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4940));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4941));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_957_17 (.CI(n40570), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4230[15]), .CO(n40571));
    SB_LUT4 duty_23__I_851_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3772[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4942));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3772[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4943));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3772[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4944));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6606_11_lut (.I0(GND_net), .I1(n17928[8]), .I2(n752_adj_4945), 
            .I3(n41340), .O(n17417[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4946));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3772[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4947));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3772[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4948));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3772[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4949));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6606_11 (.CI(n41340), .I0(n17928[8]), .I1(n752_adj_4945), 
            .CO(n41341));
    SB_LUT4 add_6606_10_lut (.I0(GND_net), .I1(n17928[7]), .I2(n679_adj_4950), 
            .I3(n41339), .O(n17417[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4951));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_6 (.CI(n40634), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n40635));
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4952));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6606_10 (.CI(n41339), .I0(n17928[7]), .I1(n679_adj_4950), 
            .CO(n41340));
    SB_LUT4 duty_23__I_851_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3772[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4953));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3772[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4954));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3772[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4955));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3772[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4956));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4958));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4960));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6606_9_lut (.I0(GND_net), .I1(n17928[6]), .I2(n606_adj_4961), 
            .I3(n41338), .O(n17417[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4963));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3772[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4964));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3772[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4965));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6606_9 (.CI(n41338), .I0(n17928[6]), .I1(n606_adj_4961), 
            .CO(n41339));
    SB_LUT4 duty_23__I_851_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3772[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4966));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6606_8_lut (.I0(GND_net), .I1(n17928[5]), .I2(n533_adj_4967), 
            .I3(n41337), .O(n17417[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_8 (.CI(n41337), .I0(n17928[5]), .I1(n533_adj_4967), 
            .CO(n41338));
    SB_LUT4 add_6606_7_lut (.I0(GND_net), .I1(n17928[4]), .I2(n460_adj_4968), 
            .I3(n41336), .O(n17417[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3772[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4969));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35784_4_lut (.I0(n21_adj_4969), .I1(n19_adj_4966), .I2(n17_adj_4965), 
            .I3(n9_adj_4964), .O(n51418));
    defparam i35784_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4970));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6606_7 (.CI(n41336), .I0(n17928[4]), .I1(n460_adj_4968), 
            .CO(n41337));
    SB_LUT4 add_6606_6_lut (.I0(GND_net), .I1(n17928[3]), .I2(n387_adj_4971), 
            .I3(n41335), .O(n17417[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n40633), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35777_4_lut (.I0(n27_adj_4956), .I1(n15_adj_4955), .I2(n13_adj_4954), 
            .I3(n11_adj_4953), .O(n51411));
    defparam i35777_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6606_6 (.CI(n41335), .I0(n17928[3]), .I1(n387_adj_4971), 
            .CO(n41336));
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4972));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i12_3_lut (.I0(duty_23__N_3772[7]), .I1(duty_23__N_3772[16]), 
            .I2(n33_adj_4963), .I3(GND_net), .O(n12_adj_4973));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6606_5_lut (.I0(GND_net), .I1(n17928[2]), .I2(n314_adj_4974), 
            .I3(n41334), .O(n17417[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i10_3_lut (.I0(duty_23__N_3772[5]), .I1(duty_23__N_3772[6]), 
            .I2(n13_adj_4954), .I3(GND_net), .O(n10_adj_4975));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6606_5 (.CI(n41334), .I0(n17928[2]), .I1(n314_adj_4974), 
            .CO(n41335));
    SB_LUT4 duty_23__I_851_i30_3_lut (.I0(n12_adj_4973), .I1(duty_23__N_3772[17]), 
            .I2(n35_adj_4949), .I3(GND_net), .O(n30_adj_4976));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6606_4_lut (.I0(GND_net), .I1(n17928[1]), .I2(n241_adj_4977), 
            .I3(n41333), .O(n17417[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_4 (.CI(n41333), .I0(n17928[1]), .I1(n241_adj_4977), 
            .CO(n41334));
    SB_LUT4 i36017_4_lut (.I0(n13_adj_4954), .I1(n11_adj_4953), .I2(n9_adj_4964), 
            .I3(n51428), .O(n51652));
    defparam i36017_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36013_4_lut (.I0(n19_adj_4966), .I1(n17_adj_4965), .I2(n15_adj_4955), 
            .I3(n51652), .O(n51648));
    defparam i36013_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36275_4_lut (.I0(n25_adj_4943), .I1(n23_adj_4942), .I2(n21_adj_4969), 
            .I3(n51648), .O(n51910));
    defparam i36275_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36129_4_lut (.I0(n31_adj_4948), .I1(n29_adj_4947), .I2(n27_adj_4956), 
            .I3(n51910), .O(n51764));
    defparam i36129_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36312_4_lut (.I0(n37_adj_4944), .I1(n35_adj_4949), .I2(n33_adj_4963), 
            .I3(n51764), .O(n51947));
    defparam i36312_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4978));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4979));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6606_3_lut (.I0(GND_net), .I1(n17928[0]), .I2(n168_adj_4980), 
            .I3(n41332), .O(n17417[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6606_3 (.CI(n41332), .I0(n17928[0]), .I1(n168_adj_4980), 
            .CO(n41333));
    SB_LUT4 add_6606_2_lut (.I0(GND_net), .I1(n26_adj_4981), .I2(n95_adj_4982), 
            .I3(GND_net), .O(n17417[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6606_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i16_3_lut (.I0(duty_23__N_3772[9]), .I1(duty_23__N_3772[21]), 
            .I2(n43_adj_4941), .I3(GND_net), .O(n16_adj_4983));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36199_3_lut (.I0(n6_adj_4786), .I1(duty_23__N_3772[10]), .I2(n21_adj_4969), 
            .I3(GND_net), .O(n51834));   // verilog/motorControl.v(36[10:25])
    defparam i36199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36200_3_lut (.I0(n51834), .I1(duty_23__N_3772[11]), .I2(n23_adj_4942), 
            .I3(GND_net), .O(n51835));   // verilog/motorControl.v(36[10:25])
    defparam i36200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i8_3_lut (.I0(duty_23__N_3772[4]), .I1(duty_23__N_3772[8]), 
            .I2(n17_adj_4965), .I3(GND_net), .O(n8_adj_4984));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i24_3_lut (.I0(n16_adj_4983), .I1(duty_23__N_3772[22]), 
            .I2(n45_adj_4940), .I3(GND_net), .O(n24_adj_4985));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35758_4_lut (.I0(n43_adj_4941), .I1(n25_adj_4943), .I2(n23_adj_4942), 
            .I3(n51418), .O(n51392));
    defparam i35758_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36177_4_lut (.I0(n24_adj_4985), .I1(n8_adj_4984), .I2(n45_adj_4940), 
            .I3(n51389), .O(n51812));   // verilog/motorControl.v(36[10:25])
    defparam i36177_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35893_3_lut (.I0(n51835), .I1(duty_23__N_3772[12]), .I2(n25_adj_4943), 
            .I3(GND_net), .O(n51528));   // verilog/motorControl.v(36[10:25])
    defparam i35893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4986));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4987));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4988));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(duty_23__N_3772[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4989));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i36197_3_lut (.I0(n4_adj_4989), .I1(duty_23__N_3772[13]), .I2(n27_adj_4956), 
            .I3(GND_net), .O(n51832));   // verilog/motorControl.v(36[10:25])
    defparam i36197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36198_3_lut (.I0(n51832), .I1(duty_23__N_3772[14]), .I2(n29_adj_4947), 
            .I3(GND_net), .O(n51833));   // verilog/motorControl.v(36[10:25])
    defparam i36198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35771_4_lut (.I0(n33_adj_4963), .I1(n31_adj_4948), .I2(n29_adj_4947), 
            .I3(n51411), .O(n51405));
    defparam i35771_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4990));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36279_4_lut (.I0(n30_adj_4976), .I1(n10_adj_4975), .I2(n35_adj_4949), 
            .I3(n51402), .O(n51914));   // verilog/motorControl.v(36[10:25])
    defparam i36279_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35895_3_lut (.I0(n51833), .I1(duty_23__N_3772[15]), .I2(n31_adj_4948), 
            .I3(GND_net), .O(n51530));   // verilog/motorControl.v(36[10:25])
    defparam i35895_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_5 (.CI(n40633), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n40634));
    SB_CARRY add_6606_2 (.CI(GND_net), .I0(n26_adj_4981), .I1(n95_adj_4982), 
            .CO(n41332));
    SB_LUT4 i36346_4_lut (.I0(n51530), .I1(n51914), .I2(n35_adj_4949), 
            .I3(n51405), .O(n51981));   // verilog/motorControl.v(36[10:25])
    defparam i36346_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36347_3_lut (.I0(n51981), .I1(duty_23__N_3772[18]), .I2(n37_adj_4944), 
            .I3(GND_net), .O(n51982));   // verilog/motorControl.v(36[10:25])
    defparam i36347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4991));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4992));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36335_3_lut (.I0(n51982), .I1(duty_23__N_3772[19]), .I2(n39_adj_4938), 
            .I3(GND_net), .O(n51970));   // verilog/motorControl.v(36[10:25])
    defparam i36335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35760_4_lut (.I0(n43_adj_4941), .I1(n41_adj_4937), .I2(n39_adj_4938), 
            .I3(n51947), .O(n51394));
    defparam i35760_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36293_4_lut (.I0(n51528), .I1(n51812), .I2(n45_adj_4940), 
            .I3(n51392), .O(n51928));   // verilog/motorControl.v(36[10:25])
    defparam i36293_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35901_3_lut (.I0(n51970), .I1(duty_23__N_3772[20]), .I2(n41_adj_4937), 
            .I3(GND_net), .O(n51536));   // verilog/motorControl.v(36[10:25])
    defparam i35901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36295_4_lut (.I0(n51536), .I1(n51928), .I2(n45_adj_4940), 
            .I3(n51394), .O(n51930));   // verilog/motorControl.v(36[10:25])
    defparam i36295_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36296_3_lut (.I0(n51930), .I1(PWMLimit[23]), .I2(duty_23__N_3772[23]), 
            .I3(GND_net), .O(duty_23__N_3771));   // verilog/motorControl.v(36[10:25])
    defparam i36296_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4994));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4995));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4996));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4997));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4999));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5001));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5002));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_5004));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_5005));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_5007));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5008));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n40632), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5009));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5010));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5011));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5012));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5013));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5015));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5016));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5017));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5018));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_5019));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5020));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5022));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5023));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5024));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5025));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5027));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_5028));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_957_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4230[14]), .I3(n40569), .O(\PID_CONTROLLER.integral_23__N_3672 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35743_4_lut (.I0(n21_adj_5027), .I1(n19_adj_5025), .I2(n17_adj_5024), 
            .I3(n9_adj_5023), .O(n51377));
    defparam i35743_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35737_4_lut (.I0(n27_adj_5022), .I1(n15_adj_5020), .I2(n13_adj_5018), 
            .I3(n11_adj_5017), .O(n51371));
    defparam i35737_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_5015), 
            .I3(GND_net), .O(n12_adj_5030));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_5031));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_5033));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_5018), 
            .I3(GND_net), .O(n10_adj_5034));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_5030), .I1(n257[17]), .I2(n35_adj_5013), 
            .I3(GND_net), .O(n30_adj_5035));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35985_4_lut (.I0(n13_adj_5018), .I1(n11_adj_5017), .I2(n9_adj_5023), 
            .I3(n51387), .O(n51620));
    defparam i35985_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35981_4_lut (.I0(n19_adj_5025), .I1(n17_adj_5024), .I2(n15_adj_5020), 
            .I3(n51620), .O(n51616));
    defparam i35981_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36269_4_lut (.I0(n25_adj_5009), .I1(n23_adj_5008), .I2(n21_adj_5027), 
            .I3(n51616), .O(n51904));
    defparam i36269_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36111_4_lut (.I0(n31_adj_5012), .I1(n29_adj_5011), .I2(n27_adj_5022), 
            .I3(n51904), .O(n51746));
    defparam i36111_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36310_4_lut (.I0(n37_adj_5010), .I1(n35_adj_5013), .I2(n33_adj_5015), 
            .I3(n51746), .O(n51945));
    defparam i36310_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_5002), 
            .I3(GND_net), .O(n16_adj_5036));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5037));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36193_3_lut (.I0(n6_adj_4783), .I1(n257[10]), .I2(n21_adj_5027), 
            .I3(GND_net), .O(n51828));   // verilog/motorControl.v(38[19:35])
    defparam i36193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36194_3_lut (.I0(n51828), .I1(n257[11]), .I2(n23_adj_5008), 
            .I3(GND_net), .O(n51829));   // verilog/motorControl.v(38[19:35])
    defparam i36194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_5024), 
            .I3(GND_net), .O(n8_adj_5039));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_5036), .I1(n257[22]), .I2(n45_adj_5001), 
            .I3(GND_net), .O(n24_adj_5040));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35720_4_lut (.I0(n43_adj_5002), .I1(n25_adj_5009), .I2(n23_adj_5008), 
            .I3(n51377), .O(n51354));
    defparam i35720_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36179_4_lut (.I0(n24_adj_5040), .I1(n8_adj_5039), .I2(n45_adj_5001), 
            .I3(n51352), .O(n51814));   // verilog/motorControl.v(38[19:35])
    defparam i36179_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35903_3_lut (.I0(n51829), .I1(n257[12]), .I2(n25_adj_5009), 
            .I3(GND_net), .O(n51538));   // verilog/motorControl.v(38[19:35])
    defparam i35903_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_957_16 (.CI(n40569), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4230[14]), .CO(n40570));
    SB_CARRY sub_3_add_2_4 (.CI(n40632), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n40633));
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(n257[1]), 
            .I2(duty_23__N_3772[1]), .I3(n257[0]), .O(n4_adj_5041));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n40631), .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5042));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36191_3_lut (.I0(n4_adj_5041), .I1(n257[13]), .I2(n27_adj_5022), 
            .I3(GND_net), .O(n51826));   // verilog/motorControl.v(38[19:35])
    defparam i36191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36192_3_lut (.I0(n51826), .I1(n257[14]), .I2(n29_adj_5011), 
            .I3(GND_net), .O(n51827));   // verilog/motorControl.v(38[19:35])
    defparam i36192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35733_4_lut (.I0(n33_adj_5015), .I1(n31_adj_5012), .I2(n29_adj_5011), 
            .I3(n51371), .O(n51367));
    defparam i35733_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36281_4_lut (.I0(n30_adj_5035), .I1(n10_adj_5034), .I2(n35_adj_5013), 
            .I3(n51365), .O(n51916));   // verilog/motorControl.v(38[19:35])
    defparam i36281_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35905_3_lut (.I0(n51827), .I1(n257[15]), .I2(n31_adj_5012), 
            .I3(GND_net), .O(n51540));   // verilog/motorControl.v(38[19:35])
    defparam i35905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36326_4_lut (.I0(n51540), .I1(n51916), .I2(n35_adj_5013), 
            .I3(n51367), .O(n51961));   // verilog/motorControl.v(38[19:35])
    defparam i36326_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36327_3_lut (.I0(n51961), .I1(n257[18]), .I2(n37_adj_5010), 
            .I3(GND_net), .O(n51962));   // verilog/motorControl.v(38[19:35])
    defparam i36327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36325_3_lut (.I0(n51962), .I1(n257[19]), .I2(n39_adj_4994), 
            .I3(GND_net), .O(n51960));   // verilog/motorControl.v(38[19:35])
    defparam i36325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35723_4_lut (.I0(n43_adj_5002), .I1(n41_adj_4995), .I2(n39_adj_4994), 
            .I3(n51945), .O(n51357));
    defparam i35723_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36297_4_lut (.I0(n51538), .I1(n51814), .I2(n45_adj_5001), 
            .I3(n51354), .O(n51932));   // verilog/motorControl.v(38[19:35])
    defparam i36297_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35911_3_lut (.I0(n51960), .I1(n257[20]), .I2(n41_adj_4995), 
            .I3(GND_net), .O(n51546));   // verilog/motorControl.v(38[19:35])
    defparam i35911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36299_4_lut (.I0(n51546), .I1(n51932), .I2(n45_adj_5001), 
            .I3(n51357), .O(n51934));   // verilog/motorControl.v(38[19:35])
    defparam i36299_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36300_3_lut (.I0(n51934), .I1(duty_23__N_3772[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_5043));   // verilog/motorControl.v(38[19:35])
    defparam i36300_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3772[0]), .I1(n257[0]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3747[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_3 (.CI(n40631), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n40632));
    SB_LUT4 add_957_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4230[13]), .I3(n40568), .O(\PID_CONTROLLER.integral_23__N_3672 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n34[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_957_15 (.CI(n40568), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4230[13]), .CO(n40569));
    SB_LUT4 add_6677_14_lut (.I0(GND_net), .I1(n18937[11]), .I2(n980), 
            .I3(n40813), .O(n18573[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6636_16_lut (.I0(GND_net), .I1(n18377[13]), .I2(n1120_adj_5044), 
            .I3(n41309), .O(n17928[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6677_13_lut (.I0(GND_net), .I1(n18937[10]), .I2(n907), 
            .I3(n40812), .O(n18573[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6636_15_lut (.I0(GND_net), .I1(n18377[12]), .I2(n1047_adj_5045), 
            .I3(n41308), .O(n17928[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_15 (.CI(n41308), .I0(n18377[12]), .I1(n1047_adj_5045), 
            .CO(n41309));
    SB_LUT4 add_6636_14_lut (.I0(GND_net), .I1(n18377[11]), .I2(n974_adj_5046), 
            .I3(n41307), .O(n17928[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_14 (.CI(n41307), .I0(n18377[11]), .I1(n974_adj_5046), 
            .CO(n41308));
    SB_CARRY add_6677_13 (.CI(n40812), .I0(n18937[10]), .I1(n907), .CO(n40813));
    SB_LUT4 add_6636_13_lut (.I0(GND_net), .I1(n18377[10]), .I2(n901_adj_5047), 
            .I3(n41306), .O(n17928[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_13 (.CI(n41306), .I0(n18377[10]), .I1(n901_adj_5047), 
            .CO(n41307));
    SB_LUT4 add_6677_12_lut (.I0(GND_net), .I1(n18937[9]), .I2(n834), 
            .I3(n40811), .O(n18573[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_12 (.CI(n40811), .I0(n18937[9]), .I1(n834), .CO(n40812));
    SB_LUT4 add_6636_12_lut (.I0(GND_net), .I1(n18377[9]), .I2(n828_adj_5048), 
            .I3(n41305), .O(n17928[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_12 (.CI(n41305), .I0(n18377[9]), .I1(n828_adj_5048), 
            .CO(n41306));
    SB_LUT4 add_6636_11_lut (.I0(GND_net), .I1(n18377[8]), .I2(n755_adj_5049), 
            .I3(n41304), .O(n17928[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_11 (.CI(n41304), .I0(n18377[8]), .I1(n755_adj_5049), 
            .CO(n41305));
    SB_LUT4 add_6636_10_lut (.I0(GND_net), .I1(n18377[7]), .I2(n682_adj_5050), 
            .I3(n41303), .O(n17928[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_10 (.CI(n41303), .I0(n18377[7]), .I1(n682_adj_5050), 
            .CO(n41304));
    SB_LUT4 add_6636_9_lut (.I0(GND_net), .I1(n18377[6]), .I2(n609_adj_5051), 
            .I3(n41302), .O(n17928[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_9 (.CI(n41302), .I0(n18377[6]), .I1(n609_adj_5051), 
            .CO(n41303));
    SB_LUT4 add_6636_8_lut (.I0(GND_net), .I1(n18377[5]), .I2(n536_adj_5052), 
            .I3(n41301), .O(n17928[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_8 (.CI(n41301), .I0(n18377[5]), .I1(n536_adj_5052), 
            .CO(n41302));
    SB_LUT4 add_6636_7_lut (.I0(GND_net), .I1(n18377[4]), .I2(n463_adj_5053), 
            .I3(n41300), .O(n17928[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_7 (.CI(n41300), .I0(n18377[4]), .I1(n463_adj_5053), 
            .CO(n41301));
    SB_LUT4 add_6636_6_lut (.I0(GND_net), .I1(n18377[3]), .I2(n390_adj_5054), 
            .I3(n41299), .O(n17928[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_6 (.CI(n41299), .I0(n18377[3]), .I1(n390_adj_5054), 
            .CO(n41300));
    SB_LUT4 add_6636_5_lut (.I0(GND_net), .I1(n18377[2]), .I2(n317_adj_5055), 
            .I3(n41298), .O(n17928[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_5 (.CI(n41298), .I0(n18377[2]), .I1(n317_adj_5055), 
            .CO(n41299));
    SB_LUT4 add_6636_4_lut (.I0(GND_net), .I1(n18377[1]), .I2(n244_adj_5056), 
            .I3(n41297), .O(n17928[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_4 (.CI(n41297), .I0(n18377[1]), .I1(n244_adj_5056), 
            .CO(n41298));
    SB_LUT4 add_6636_3_lut (.I0(GND_net), .I1(n18377[0]), .I2(n171_adj_5057), 
            .I3(n41296), .O(n17928[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6636_3 (.CI(n41296), .I0(n18377[0]), .I1(n171_adj_5057), 
            .CO(n41297));
    SB_LUT4 add_6677_11_lut (.I0(GND_net), .I1(n18937[8]), .I2(n761), 
            .I3(n40810), .O(n18573[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_11 (.CI(n40810), .I0(n18937[8]), .I1(n761), .CO(n40811));
    SB_LUT4 add_6636_2_lut (.I0(GND_net), .I1(n29_adj_5058), .I2(n98_adj_5059), 
            .I3(GND_net), .O(n17928[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6636_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6677_10_lut (.I0(GND_net), .I1(n18937[7]), .I2(n688), 
            .I3(n40809), .O(n18573[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n40631));
    SB_CARRY add_6636_2 (.CI(GND_net), .I0(n29_adj_5058), .I1(n98_adj_5059), 
            .CO(n41296));
    SB_LUT4 add_6664_15_lut (.I0(GND_net), .I1(n18768[12]), .I2(n1050_adj_5060), 
            .I3(n41295), .O(n18377[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6664_14_lut (.I0(GND_net), .I1(n18768[11]), .I2(n977_adj_5061), 
            .I3(n41294), .O(n18377[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_14 (.CI(n41294), .I0(n18768[11]), .I1(n977_adj_5061), 
            .CO(n41295));
    SB_LUT4 add_6664_13_lut (.I0(GND_net), .I1(n18768[10]), .I2(n904_adj_5062), 
            .I3(n41293), .O(n18377[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_13 (.CI(n41293), .I0(n18768[10]), .I1(n904_adj_5062), 
            .CO(n41294));
    SB_LUT4 add_6664_12_lut (.I0(GND_net), .I1(n18768[9]), .I2(n831_adj_5063), 
            .I3(n41292), .O(n18377[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_12 (.CI(n41292), .I0(n18768[9]), .I1(n831_adj_5063), 
            .CO(n41293));
    SB_LUT4 add_6664_11_lut (.I0(GND_net), .I1(n18768[8]), .I2(n758_adj_5064), 
            .I3(n41291), .O(n18377[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_11 (.CI(n41291), .I0(n18768[8]), .I1(n758_adj_5064), 
            .CO(n41292));
    SB_LUT4 add_6664_10_lut (.I0(GND_net), .I1(n18768[7]), .I2(n685_adj_5065), 
            .I3(n41290), .O(n18377[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_10 (.CI(n41290), .I0(n18768[7]), .I1(n685_adj_5065), 
            .CO(n41291));
    SB_CARRY add_6677_10 (.CI(n40809), .I0(n18937[7]), .I1(n688), .CO(n40810));
    SB_LUT4 add_6664_9_lut (.I0(GND_net), .I1(n18768[6]), .I2(n612_adj_5066), 
            .I3(n41289), .O(n18377[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_9 (.CI(n41289), .I0(n18768[6]), .I1(n612_adj_5066), 
            .CO(n41290));
    SB_LUT4 add_6664_8_lut (.I0(GND_net), .I1(n18768[5]), .I2(n539_adj_5067), 
            .I3(n41288), .O(n18377[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_8 (.CI(n41288), .I0(n18768[5]), .I1(n539_adj_5067), 
            .CO(n41289));
    SB_LUT4 add_6677_9_lut (.I0(GND_net), .I1(n18937[6]), .I2(n615), .I3(n40808), 
            .O(n18573[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6664_7_lut (.I0(GND_net), .I1(n18768[4]), .I2(n466_adj_5068), 
            .I3(n41287), .O(n18377[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_7 (.CI(n41287), .I0(n18768[4]), .I1(n466_adj_5068), 
            .CO(n41288));
    SB_LUT4 add_6664_6_lut (.I0(GND_net), .I1(n18768[3]), .I2(n393_adj_5069), 
            .I3(n41286), .O(n18377[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_6 (.CI(n41286), .I0(n18768[3]), .I1(n393_adj_5069), 
            .CO(n41287));
    SB_CARRY add_6677_9 (.CI(n40808), .I0(n18937[6]), .I1(n615), .CO(n40809));
    SB_LUT4 add_957_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4230[12]), .I3(n40567), .O(\PID_CONTROLLER.integral_23__N_3672 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6664_5_lut (.I0(GND_net), .I1(n18768[2]), .I2(n320_adj_5070), 
            .I3(n41285), .O(n18377[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_5 (.CI(n41285), .I0(n18768[2]), .I1(n320_adj_5070), 
            .CO(n41286));
    SB_LUT4 add_6664_4_lut (.I0(GND_net), .I1(n18768[1]), .I2(n247_adj_5071), 
            .I3(n41284), .O(n18377[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_4 (.CI(n41284), .I0(n18768[1]), .I1(n247_adj_5071), 
            .CO(n41285));
    SB_LUT4 add_6677_8_lut (.I0(GND_net), .I1(n18937[5]), .I2(n542), .I3(n40807), 
            .O(n18573[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6664_3_lut (.I0(GND_net), .I1(n18768[0]), .I2(n174_adj_5072), 
            .I3(n41283), .O(n18377[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_3 (.CI(n41283), .I0(n18768[0]), .I1(n174_adj_5072), 
            .CO(n41284));
    SB_LUT4 add_6664_2_lut (.I0(GND_net), .I1(n32_adj_5073), .I2(n101_adj_5074), 
            .I3(GND_net), .O(n18377[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6664_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6664_2 (.CI(GND_net), .I0(n32_adj_5073), .I1(n101_adj_5074), 
            .CO(n41283));
    SB_LUT4 add_6690_14_lut (.I0(GND_net), .I1(n19105[11]), .I2(n980_adj_5075), 
            .I3(n41282), .O(n18768[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6690_13_lut (.I0(GND_net), .I1(n19105[10]), .I2(n907_adj_5076), 
            .I3(n41281), .O(n18768[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_8 (.CI(n40807), .I0(n18937[5]), .I1(n542), .CO(n40808));
    SB_LUT4 add_6677_7_lut (.I0(GND_net), .I1(n18937[4]), .I2(n469), .I3(n40806), 
            .O(n18573[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_13 (.CI(n41281), .I0(n19105[10]), .I1(n907_adj_5076), 
            .CO(n41282));
    SB_LUT4 add_6690_12_lut (.I0(GND_net), .I1(n19105[9]), .I2(n834_adj_5077), 
            .I3(n41280), .O(n18768[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_12 (.CI(n41280), .I0(n19105[9]), .I1(n834_adj_5077), 
            .CO(n41281));
    SB_LUT4 add_6690_11_lut (.I0(GND_net), .I1(n19105[8]), .I2(n761_adj_5078), 
            .I3(n41279), .O(n18768[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_7 (.CI(n40806), .I0(n18937[4]), .I1(n469), .CO(n40807));
    SB_CARRY add_6690_11 (.CI(n41279), .I0(n19105[8]), .I1(n761_adj_5078), 
            .CO(n41280));
    SB_LUT4 add_6690_10_lut (.I0(GND_net), .I1(n19105[7]), .I2(n688_adj_5079), 
            .I3(n41278), .O(n18768[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_10 (.CI(n41278), .I0(n19105[7]), .I1(n688_adj_5079), 
            .CO(n41279));
    SB_LUT4 add_6690_9_lut (.I0(GND_net), .I1(n19105[6]), .I2(n615_adj_5080), 
            .I3(n41277), .O(n18768[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_9 (.CI(n41277), .I0(n19105[6]), .I1(n615_adj_5080), 
            .CO(n41278));
    SB_LUT4 add_6690_8_lut (.I0(GND_net), .I1(n19105[5]), .I2(n542_adj_5081), 
            .I3(n41276), .O(n18768[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_8 (.CI(n41276), .I0(n19105[5]), .I1(n542_adj_5081), 
            .CO(n41277));
    SB_LUT4 add_6690_7_lut (.I0(GND_net), .I1(n19105[4]), .I2(n469_adj_5082), 
            .I3(n41275), .O(n18768[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_7 (.CI(n41275), .I0(n19105[4]), .I1(n469_adj_5082), 
            .CO(n41276));
    SB_LUT4 add_6690_6_lut (.I0(GND_net), .I1(n19105[3]), .I2(n396), .I3(n41274), 
            .O(n18768[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_6 (.CI(n41274), .I0(n19105[3]), .I1(n396), .CO(n41275));
    SB_LUT4 add_6690_5_lut (.I0(GND_net), .I1(n19105[2]), .I2(n323), .I3(n41273), 
            .O(n18768[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_5 (.CI(n41273), .I0(n19105[2]), .I1(n323), .CO(n41274));
    SB_LUT4 add_6690_4_lut (.I0(GND_net), .I1(n19105[1]), .I2(n250), .I3(n41272), 
            .O(n18768[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_4 (.CI(n41272), .I0(n19105[1]), .I1(n250), .CO(n41273));
    SB_LUT4 add_6690_3_lut (.I0(GND_net), .I1(n19105[0]), .I2(n177), .I3(n41271), 
            .O(n18768[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_3 (.CI(n41271), .I0(n19105[0]), .I1(n177), .CO(n41272));
    SB_LUT4 add_6690_2_lut (.I0(GND_net), .I1(n35_adj_5083), .I2(n104_adj_5084), 
            .I3(GND_net), .O(n18768[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6690_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6690_2 (.CI(GND_net), .I0(n35_adj_5083), .I1(n104_adj_5084), 
            .CO(n41271));
    SB_LUT4 add_6714_13_lut (.I0(GND_net), .I1(n19392[10]), .I2(n910_adj_5085), 
            .I3(n41270), .O(n19105[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6677_6_lut (.I0(GND_net), .I1(n18937[3]), .I2(n396_adj_5086), 
            .I3(n40805), .O(n18573[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6714_12_lut (.I0(GND_net), .I1(n19392[9]), .I2(n837_adj_5087), 
            .I3(n41269), .O(n19105[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_6 (.CI(n40805), .I0(n18937[3]), .I1(n396_adj_5086), 
            .CO(n40806));
    SB_CARRY add_6714_12 (.CI(n41269), .I0(n19392[9]), .I1(n837_adj_5087), 
            .CO(n41270));
    SB_LUT4 add_6714_11_lut (.I0(GND_net), .I1(n19392[8]), .I2(n764_adj_5088), 
            .I3(n41268), .O(n19105[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_11 (.CI(n41268), .I0(n19392[8]), .I1(n764_adj_5088), 
            .CO(n41269));
    SB_LUT4 add_6714_10_lut (.I0(GND_net), .I1(n19392[7]), .I2(n691_adj_5089), 
            .I3(n41267), .O(n19105[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_10 (.CI(n41267), .I0(n19392[7]), .I1(n691_adj_5089), 
            .CO(n41268));
    SB_LUT4 add_6714_9_lut (.I0(GND_net), .I1(n19392[6]), .I2(n618_adj_5090), 
            .I3(n41266), .O(n19105[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_9 (.CI(n41266), .I0(n19392[6]), .I1(n618_adj_5090), 
            .CO(n41267));
    SB_LUT4 add_6714_8_lut (.I0(GND_net), .I1(n19392[5]), .I2(n545_adj_5091), 
            .I3(n41265), .O(n19105[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_8 (.CI(n41265), .I0(n19392[5]), .I1(n545_adj_5091), 
            .CO(n41266));
    SB_LUT4 add_6714_7_lut (.I0(GND_net), .I1(n19392[4]), .I2(n472_adj_5092), 
            .I3(n41264), .O(n19105[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_7 (.CI(n41264), .I0(n19392[4]), .I1(n472_adj_5092), 
            .CO(n41265));
    SB_LUT4 add_6677_5_lut (.I0(GND_net), .I1(n18937[2]), .I2(n323_adj_5093), 
            .I3(n40804), .O(n18573[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6714_6_lut (.I0(GND_net), .I1(n19392[3]), .I2(n399_adj_5094), 
            .I3(n41263), .O(n19105[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_6 (.CI(n41263), .I0(n19392[3]), .I1(n399_adj_5094), 
            .CO(n41264));
    SB_CARRY add_6677_5 (.CI(n40804), .I0(n18937[2]), .I1(n323_adj_5093), 
            .CO(n40805));
    SB_LUT4 add_6714_5_lut (.I0(GND_net), .I1(n19392[2]), .I2(n326_adj_5095), 
            .I3(n41262), .O(n19105[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6677_4_lut (.I0(GND_net), .I1(n18937[1]), .I2(n250_adj_5096), 
            .I3(n40803), .O(n18573[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_4 (.CI(n40803), .I0(n18937[1]), .I1(n250_adj_5096), 
            .CO(n40804));
    SB_CARRY add_6714_5 (.CI(n41262), .I0(n19392[2]), .I1(n326_adj_5095), 
            .CO(n41263));
    SB_LUT4 add_6714_4_lut (.I0(GND_net), .I1(n19392[1]), .I2(n253_adj_5097), 
            .I3(n41261), .O(n19105[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_4 (.CI(n41261), .I0(n19392[1]), .I1(n253_adj_5097), 
            .CO(n41262));
    SB_LUT4 add_6677_3_lut (.I0(GND_net), .I1(n18937[0]), .I2(n177_adj_5098), 
            .I3(n40802), .O(n18573[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6714_3_lut (.I0(GND_net), .I1(n19392[0]), .I2(n180_adj_5099), 
            .I3(n41260), .O(n19105[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_3 (.CI(n41260), .I0(n19392[0]), .I1(n180_adj_5099), 
            .CO(n41261));
    SB_CARRY add_6677_3 (.CI(n40802), .I0(n18937[0]), .I1(n177_adj_5098), 
            .CO(n40803));
    SB_LUT4 add_6677_2_lut (.I0(GND_net), .I1(n35_adj_5042), .I2(n104), 
            .I3(GND_net), .O(n18573[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6677_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6677_2 (.CI(GND_net), .I0(n35_adj_5042), .I1(n104), .CO(n40802));
    SB_LUT4 add_6714_2_lut (.I0(GND_net), .I1(n38_adj_5038), .I2(n107_adj_5037), 
            .I3(GND_net), .O(n19105[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6714_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6714_2 (.CI(GND_net), .I0(n38_adj_5038), .I1(n107_adj_5037), 
            .CO(n41260));
    SB_CARRY add_957_14 (.CI(n40567), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4230[12]), .CO(n40568));
    SB_LUT4 add_6702_13_lut (.I0(GND_net), .I1(n19249[10]), .I2(n910), 
            .I3(n40801), .O(n18937[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6702_12_lut (.I0(GND_net), .I1(n19249[9]), .I2(n837), 
            .I3(n40800), .O(n18937[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_12 (.CI(n40800), .I0(n19249[9]), .I1(n837), .CO(n40801));
    SB_LUT4 add_6736_12_lut (.I0(GND_net), .I1(n19633[9]), .I2(n840_adj_4844), 
            .I3(n41238), .O(n19392[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6736_11_lut (.I0(GND_net), .I1(n19633[8]), .I2(n767_adj_4843), 
            .I3(n41237), .O(n19392[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_11 (.CI(n41237), .I0(n19633[8]), .I1(n767_adj_4843), 
            .CO(n41238));
    SB_LUT4 add_6736_10_lut (.I0(GND_net), .I1(n19633[7]), .I2(n694_adj_4842), 
            .I3(n41236), .O(n19392[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_10 (.CI(n41236), .I0(n19633[7]), .I1(n694_adj_4842), 
            .CO(n41237));
    SB_LUT4 add_6736_9_lut (.I0(GND_net), .I1(n19633[6]), .I2(n621_adj_4840), 
            .I3(n41235), .O(n19392[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_9 (.CI(n41235), .I0(n19633[6]), .I1(n621_adj_4840), 
            .CO(n41236));
    SB_LUT4 add_6736_8_lut (.I0(GND_net), .I1(n19633[5]), .I2(n548_adj_4839), 
            .I3(n41234), .O(n19392[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6702_11_lut (.I0(GND_net), .I1(n19249[8]), .I2(n764), 
            .I3(n40799), .O(n18937[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_8 (.CI(n41234), .I0(n19633[5]), .I1(n548_adj_4839), 
            .CO(n41235));
    SB_LUT4 add_6736_7_lut (.I0(GND_net), .I1(n19633[4]), .I2(n475_adj_4838), 
            .I3(n41233), .O(n19392[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6736_7 (.CI(n41233), .I0(n19633[4]), .I1(n475_adj_4838), 
            .CO(n41234));
    SB_LUT4 add_957_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4230[11]), .I3(n40566), .O(\PID_CONTROLLER.integral_23__N_3672 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6736_6_lut (.I0(GND_net), .I1(n19633[3]), .I2(n402_adj_4836), 
            .I3(n41232), .O(n19392[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_13 (.CI(n40566), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4230[11]), .CO(n40567));
    SB_CARRY add_6736_6 (.CI(n41232), .I0(n19633[3]), .I1(n402_adj_4836), 
            .CO(n41233));
    SB_CARRY add_6702_11 (.CI(n40799), .I0(n19249[8]), .I1(n764), .CO(n40800));
    SB_LUT4 add_6736_5_lut (.I0(GND_net), .I1(n19633[2]), .I2(n329_adj_4835), 
            .I3(n41231), .O(n19392[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_5 (.CI(n41231), .I0(n19633[2]), .I1(n329_adj_4835), 
            .CO(n41232));
    SB_LUT4 add_6736_4_lut (.I0(GND_net), .I1(n19633[1]), .I2(n256_adj_4834), 
            .I3(n41230), .O(n19392[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_4 (.CI(n41230), .I0(n19633[1]), .I1(n256_adj_4834), 
            .CO(n41231));
    SB_LUT4 add_6736_3_lut (.I0(GND_net), .I1(n19633[0]), .I2(n183_adj_4833), 
            .I3(n41229), .O(n19392[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_3 (.CI(n41229), .I0(n19633[0]), .I1(n183_adj_4833), 
            .CO(n41230));
    SB_LUT4 add_6736_2_lut (.I0(GND_net), .I1(n41_adj_4832), .I2(n110_adj_4830), 
            .I3(GND_net), .O(n19392[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6736_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6736_2 (.CI(GND_net), .I0(n41_adj_4832), .I1(n110_adj_4830), 
            .CO(n41229));
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6702_10_lut (.I0(GND_net), .I1(n19249[7]), .I2(n691), 
            .I3(n40798), .O(n18937[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_10 (.CI(n40798), .I0(n19249[7]), .I1(n691), .CO(n40799));
    SB_LUT4 add_6702_9_lut (.I0(GND_net), .I1(n19249[6]), .I2(n618), .I3(n40797), 
            .O(n18937[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_957_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4230[10]), .I3(n40565), .O(\PID_CONTROLLER.integral_23__N_3672 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_9 (.CI(n40797), .I0(n19249[6]), .I1(n618), .CO(n40798));
    SB_CARRY add_957_12 (.CI(n40565), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4230[10]), .CO(n40566));
    SB_LUT4 add_6702_8_lut (.I0(GND_net), .I1(n19249[5]), .I2(n545), .I3(n40796), 
            .O(n18937[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_957_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4230[9]), .I3(n40564), .O(\PID_CONTROLLER.integral_23__N_3672 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_11 (.CI(n40564), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4230[9]), .CO(n40565));
    SB_LUT4 add_957_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4230[8]), .I3(n40563), .O(\PID_CONTROLLER.integral_23__N_3672 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_8 (.CI(n40796), .I0(n19249[5]), .I1(n545), .CO(n40797));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6702_7_lut (.I0(GND_net), .I1(n19249[4]), .I2(n472), .I3(n40795), 
            .O(n18937[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6702_7 (.CI(n40795), .I0(n19249[4]), .I1(n472), .CO(n40796));
    SB_CARRY add_957_10 (.CI(n40563), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4230[8]), .CO(n40564));
    SB_LUT4 add_957_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4230[7]), .I3(n40562), .O(\PID_CONTROLLER.integral_23__N_3672 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6702_6_lut (.I0(GND_net), .I1(n19249[3]), .I2(n399), .I3(n40794), 
            .O(n18937[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_9 (.CI(n40562), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4230[7]), .CO(n40563));
    SB_CARRY add_6702_6 (.CI(n40794), .I0(n19249[3]), .I1(n399), .CO(n40795));
    SB_LUT4 add_957_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4230[6]), .I3(n40561), .O(\PID_CONTROLLER.integral_23__N_3672 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_957_8 (.CI(n40561), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4230[6]), .CO(n40562));
    SB_LUT4 add_6702_5_lut (.I0(GND_net), .I1(n19249[2]), .I2(n326), .I3(n40793), 
            .O(n18937[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_5 (.CI(n40793), .I0(n19249[2]), .I1(n326), .CO(n40794));
    SB_LUT4 add_957_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4230[5]), .I3(n40560), .O(\PID_CONTROLLER.integral_23__N_3672 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6702_4_lut (.I0(GND_net), .I1(n19249[1]), .I2(n253), .I3(n40792), 
            .O(n18937[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6702_4 (.CI(n40792), .I0(n19249[1]), .I1(n253), .CO(n40793));
    SB_LUT4 add_6702_3_lut (.I0(GND_net), .I1(n19249[0]), .I2(n180), .I3(n40791), 
            .O(n18937[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_7 (.CI(n40560), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4230[5]), .CO(n40561));
    SB_LUT4 add_957_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4230[4]), .I3(n40559), .O(\PID_CONTROLLER.integral_23__N_3672 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_6 (.CI(n40559), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4230[4]), .CO(n40560));
    SB_CARRY add_6702_3 (.CI(n40791), .I0(n19249[0]), .I1(n180), .CO(n40792));
    SB_LUT4 add_6702_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n18937[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6702_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6702_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n40791));
    SB_LUT4 add_957_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4230[3]), .I3(n40558), .O(\PID_CONTROLLER.integral_23__N_3672 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_5 (.CI(n40558), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4230[3]), .CO(n40559));
    SB_LUT4 add_957_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4230[2]), .I3(n40557), .O(\PID_CONTROLLER.integral_23__N_3672 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6816_7_lut (.I0(GND_net), .I1(n48333), .I2(n490_adj_4799), 
            .I3(n40790), .O(n20217[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6816_6_lut (.I0(GND_net), .I1(n20288[3]), .I2(n417), .I3(n40789), 
            .O(n20217[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_4 (.CI(n40557), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4230[2]), .CO(n40558));
    SB_CARRY add_6816_6 (.CI(n40789), .I0(n20288[3]), .I1(n417), .CO(n40790));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[23]), 
            .I3(n40699), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6816_5_lut (.I0(GND_net), .I1(n20288[2]), .I2(n344), .I3(n40788), 
            .O(n20217[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[22]), 
            .I3(n40698), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_957_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4230[1]), .I3(n40556), .O(\PID_CONTROLLER.integral_23__N_3672 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_3 (.CI(n40556), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4230[1]), .CO(n40557));
    SB_CARRY add_6816_5 (.CI(n40788), .I0(n20288[2]), .I1(n344), .CO(n40789));
    SB_LUT4 add_957_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4230[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3672 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_957_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6816_4_lut (.I0(GND_net), .I1(n20288[1]), .I2(n271), .I3(n40787), 
            .O(n20217[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_957_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4230[0]), .CO(n40556));
    SB_CARRY add_6816_4 (.CI(n40787), .I0(n20288[1]), .I1(n271), .CO(n40788));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n40698), .I0(GND_net), .I1(n1_adj_5153[22]), 
            .CO(n40699));
    SB_LUT4 add_6816_3_lut (.I0(GND_net), .I1(n20288[0]), .I2(n198), .I3(n40786), 
            .O(n20217[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6816_3 (.CI(n40786), .I0(n20288[0]), .I1(n198), .CO(n40787));
    SB_LUT4 add_6816_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20217[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6816_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6816_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n40786));
    SB_LUT4 add_6725_12_lut (.I0(GND_net), .I1(n19513[9]), .I2(n840), 
            .I3(n40785), .O(n19249[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6725_11_lut (.I0(GND_net), .I1(n19513[8]), .I2(n767), 
            .I3(n40784), .O(n19249[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[21]), 
            .I3(n40697), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n40697), .I0(GND_net), .I1(n1_adj_5153[21]), 
            .CO(n40698));
    SB_CARRY add_6725_11 (.CI(n40784), .I0(n19513[8]), .I1(n767), .CO(n40785));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[20]), 
            .I3(n40696), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n40696), .I0(GND_net), .I1(n1_adj_5153[20]), 
            .CO(n40697));
    SB_LUT4 add_6725_10_lut (.I0(GND_net), .I1(n19513[7]), .I2(n694), 
            .I3(n40783), .O(n19249[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_5098));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5097));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_5096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5095));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[19]), 
            .I3(n40695), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_10 (.CI(n40783), .I0(n19513[7]), .I1(n694), .CO(n40784));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n40695), .I0(GND_net), .I1(n1_adj_5153[19]), 
            .CO(n40696));
    SB_LUT4 i26500_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n40150), .I3(n20377[0]), .O(n4_adj_4732));   // verilog/motorControl.v(34[25:36])
    defparam i26500_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_6725_9_lut (.I0(GND_net), .I1(n19513[6]), .I2(n621), .I3(n40782), 
            .O(n19249[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5094));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[18]), 
            .I3(n40694), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6725_9 (.CI(n40782), .I0(n19513[6]), .I1(n621), .CO(n40783));
    SB_CARRY unary_minus_16_add_3_20 (.CI(n40694), .I0(GND_net), .I1(n1_adj_5153[18]), 
            .CO(n40695));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[17]), 
            .I3(n40693), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6725_8_lut (.I0(GND_net), .I1(n19513[5]), .I2(n548), .I3(n40781), 
            .O(n19249[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_8 (.CI(n40781), .I0(n19513[5]), .I1(n548), .CO(n40782));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n40693), .I0(GND_net), .I1(n1_adj_5153[17]), 
            .CO(n40694));
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n10669[0]), .I2(n10138[0]), 
            .I3(n40550), .O(duty_23__N_3772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_5093));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5092));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5091));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[16]), 
            .I3(n40692), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6725_7_lut (.I0(GND_net), .I1(n19513[4]), .I2(n475), .I3(n40780), 
            .O(n19249[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n40692), .I0(GND_net), .I1(n1_adj_5153[16]), 
            .CO(n40693));
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n40549), .O(duty_23__N_3772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_7 (.CI(n40780), .I0(n19513[4]), .I1(n475), .CO(n40781));
    SB_LUT4 add_6725_6_lut (.I0(GND_net), .I1(n19513[3]), .I2(n402), .I3(n40779), 
            .O(n19249[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_6 (.CI(n40779), .I0(n19513[3]), .I1(n402), .CO(n40780));
    SB_LUT4 add_6725_5_lut (.I0(GND_net), .I1(n19513[2]), .I2(n329), .I3(n40778), 
            .O(n19249[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[15]), 
            .I3(n40691), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n40691), .I0(GND_net), .I1(n1_adj_5153[15]), 
            .CO(n40692));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[14]), 
            .I3(n40690), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_5 (.CI(n40778), .I0(n19513[2]), .I1(n329), .CO(n40779));
    SB_CARRY add_12_24 (.CI(n40549), .I0(n106[22]), .I1(n155[22]), .CO(n40550));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n40690), .I0(GND_net), .I1(n1_adj_5153[14]), 
            .CO(n40691));
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n40548), .O(duty_23__N_3772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n40548), .I0(n106[21]), .I1(n155[21]), .CO(n40549));
    SB_LUT4 add_6725_4_lut (.I0(GND_net), .I1(n19513[1]), .I2(n256), .I3(n40777), 
            .O(n19249[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[13]), 
            .I3(n40689), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_4 (.CI(n40777), .I0(n19513[1]), .I1(n256), .CO(n40778));
    SB_CARRY unary_minus_16_add_3_15 (.CI(n40689), .I0(GND_net), .I1(n1_adj_5153[13]), 
            .CO(n40690));
    SB_LUT4 add_6725_3_lut (.I0(GND_net), .I1(n19513[0]), .I2(n183), .I3(n40776), 
            .O(n19249[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_3 (.CI(n40776), .I0(n19513[0]), .I1(n183), .CO(n40777));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n40547), .O(duty_23__N_3772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[12]), 
            .I3(n40688), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n40547), .I0(n106[20]), .I1(n155[20]), .CO(n40548));
    SB_LUT4 add_6725_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n19249[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6725_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n40688), .I0(GND_net), .I1(n1_adj_5153[12]), 
            .CO(n40689));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[11]), 
            .I3(n40687), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6725_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n40776));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n40687), .I0(GND_net), .I1(n1_adj_5153[11]), 
            .CO(n40688));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[10]), 
            .I3(n40686), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n40686), .I0(GND_net), .I1(n1_adj_5153[10]), 
            .CO(n40687));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[9]), 
            .I3(n40685), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n40546), .O(duty_23__N_3772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n40546), .I0(n106[19]), .I1(n155[19]), .CO(n40547));
    SB_CARRY unary_minus_16_add_3_11 (.CI(n40685), .I0(GND_net), .I1(n1_adj_5153[9]), 
            .CO(n40686));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[8]), 
            .I3(n40684), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n40684), .I0(GND_net), .I1(n1_adj_5153[8]), 
            .CO(n40685));
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_5090));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_5101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_5103));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[7]), 
            .I3(n40683), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n40545), .O(duty_23__N_3772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n40545), .I0(n106[18]), .I1(n155[18]), .CO(n40546));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n40683), .I0(GND_net), .I1(n1_adj_5153[7]), 
            .CO(n40684));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n40544), .O(duty_23__N_3772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n40544), .I0(n106[17]), .I1(n155[17]), .CO(n40545));
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_5105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_5089));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5088));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[6]), 
            .I3(n40682), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5087));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_5086));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5085));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n20377[0]), .I3(n40150), .O(n20353[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5084));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n40543), .O(duty_23__N_3772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5083));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n34[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1521 (.I0(n62), .I1(n131), .I2(n20353[0]), 
            .I3(n204), .O(n20313[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1521.LUT_INIT = 16'h8778;
    SB_CARRY add_12_18 (.CI(n40543), .I0(n106[16]), .I1(n155[16]), .CO(n40544));
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n40542), .O(duty_23__N_3772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n40682), .I0(GND_net), .I1(n1_adj_5153[6]), 
            .CO(n40683));
    SB_LUT4 i26538_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n20353[0]), 
            .O(n4));   // verilog/motorControl.v(34[25:36])
    defparam i26538_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_12_17 (.CI(n40542), .I0(n106[15]), .I1(n155[15]), .CO(n40543));
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n40541), .O(duty_23__N_3772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n40541), .I0(n106[14]), .I1(n155[14]), .CO(n40542));
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n40540), .O(duty_23__N_3772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I1(n10645[21]), .I2(GND_net), .I3(n41033), .O(n10138[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10645[20]), .I2(GND_net), 
            .I3(n41032), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n40540), .I0(n106[13]), .I1(n155[13]), .CO(n40541));
    SB_CARRY mult_11_add_1225_23 (.CI(n41032), .I0(n10645[20]), .I1(GND_net), 
            .CO(n41033));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10645[19]), .I2(GND_net), 
            .I3(n41031), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n41031), .I0(n10645[19]), .I1(GND_net), 
            .CO(n41032));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10645[18]), .I2(GND_net), 
            .I3(n41030), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n41030), .I0(n10645[18]), .I1(GND_net), 
            .CO(n41031));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10645[17]), .I2(GND_net), 
            .I3(n41029), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n41029), .I0(n10645[17]), .I1(GND_net), 
            .CO(n41030));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10645[16]), .I2(GND_net), 
            .I3(n41028), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n41028), .I0(n10645[16]), .I1(GND_net), 
            .CO(n41029));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10645[15]), .I2(GND_net), 
            .I3(n41027), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n41027), .I0(n10645[15]), .I1(GND_net), 
            .CO(n41028));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10645[14]), .I2(GND_net), 
            .I3(n41026), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n41026), .I0(n10645[14]), .I1(GND_net), 
            .CO(n41027));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10645[13]), .I2(n1096), 
            .I3(n41025), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n41025), .I0(n10645[13]), .I1(n1096), 
            .CO(n41026));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10645[12]), .I2(n1023), 
            .I3(n41024), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n41024), .I0(n10645[12]), .I1(n1023), 
            .CO(n41025));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10645[11]), .I2(n950), 
            .I3(n41023), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n41023), .I0(n10645[11]), .I1(n950), 
            .CO(n41024));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10645[10]), .I2(n877), 
            .I3(n41022), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n41022), .I0(n10645[10]), .I1(n877), 
            .CO(n41023));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10645[9]), .I2(n804), 
            .I3(n41021), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n41021), .I0(n10645[9]), .I1(n804), 
            .CO(n41022));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10645[8]), .I2(n731), 
            .I3(n41020), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n41020), .I0(n10645[8]), .I1(n731), 
            .CO(n41021));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10645[7]), .I2(n658), 
            .I3(n41019), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n41019), .I0(n10645[7]), .I1(n658), 
            .CO(n41020));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10645[6]), .I2(n585), 
            .I3(n41018), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n41018), .I0(n10645[6]), .I1(n585), 
            .CO(n41019));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10645[5]), .I2(n512), 
            .I3(n41017), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n41017), .I0(n10645[5]), .I1(n512), 
            .CO(n41018));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10645[4]), .I2(n439), 
            .I3(n41016), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n41016), .I0(n10645[4]), .I1(n439), 
            .CO(n41017));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10645[3]), .I2(n366), 
            .I3(n41015), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n41015), .I0(n10645[3]), .I1(n366), 
            .CO(n41016));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10645[2]), .I2(n293), 
            .I3(n41014), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n41014), .I0(n10645[2]), .I1(n293), 
            .CO(n41015));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10645[1]), .I2(n220), 
            .I3(n41013), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n41013), .I0(n10645[1]), .I1(n220), 
            .CO(n41014));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10645[0]), .I2(n147), 
            .I3(n41012), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n41012), .I0(n10645[0]), .I1(n147), 
            .CO(n41013));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5082));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5081));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5080));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5079));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5078));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5077));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n41012));
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[5]), 
            .I3(n40681), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5076));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n40539), .O(duty_23__N_3772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n40539), .I0(n106[12]), .I1(n155[12]), .CO(n40540));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n40538), .O(duty_23__N_3772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5075));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_13 (.CI(n40538), .I0(n106[11]), .I1(n155[11]), .CO(n40539));
    SB_LUT4 add_4786_23_lut (.I0(GND_net), .I1(n12653[20]), .I2(GND_net), 
            .I3(n41003), .O(n10645[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_5074));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_22_lut (.I0(GND_net), .I1(n12653[19]), .I2(GND_net), 
            .I3(n41002), .O(n10645[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n40681), .I0(GND_net), .I1(n1_adj_5153[5]), 
            .CO(n40682));
    SB_CARRY add_4786_22 (.CI(n41002), .I0(n12653[19]), .I1(GND_net), 
            .CO(n41003));
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_5073));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_5072));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_21_lut (.I0(GND_net), .I1(n12653[18]), .I2(GND_net), 
            .I3(n41001), .O(n10645[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_5071));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[4]), 
            .I3(n40680), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n40680), .I0(GND_net), .I1(n1_adj_5153[4]), 
            .CO(n40681));
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_5070));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22150_2_lut (.I0(n34[12]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_5069));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_5068));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[3]), 
            .I3(n40679), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_21 (.CI(n41001), .I0(n12653[18]), .I1(GND_net), 
            .CO(n41002));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n40537), .O(duty_23__N_3772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n40537), .I0(n106[10]), .I1(n155[10]), .CO(n40538));
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_5067));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_20_lut (.I0(GND_net), .I1(n12653[17]), .I2(GND_net), 
            .I3(n41000), .O(n10645[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_20 (.CI(n41000), .I0(n12653[17]), .I1(GND_net), 
            .CO(n41001));
    SB_LUT4 add_4786_19_lut (.I0(GND_net), .I1(n12653[16]), .I2(GND_net), 
            .I3(n40999), .O(n10645[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_5066));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_5065));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_5064));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4786_19 (.CI(n40999), .I0(n12653[16]), .I1(GND_net), 
            .CO(n41000));
    SB_LUT4 add_4786_18_lut (.I0(GND_net), .I1(n12653[15]), .I2(GND_net), 
            .I3(n40998), .O(n10645[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_18 (.CI(n40998), .I0(n12653[15]), .I1(GND_net), 
            .CO(n40999));
    SB_LUT4 add_4786_17_lut (.I0(GND_net), .I1(n12653[14]), .I2(GND_net), 
            .I3(n40997), .O(n10645[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_17 (.CI(n40997), .I0(n12653[14]), .I1(GND_net), 
            .CO(n40998));
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_5063));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_16_lut (.I0(GND_net), .I1(n12653[13]), .I2(n1099_adj_5112), 
            .I3(n40996), .O(n10645[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_16 (.CI(n40996), .I0(n12653[13]), .I1(n1099_adj_5112), 
            .CO(n40997));
    SB_LUT4 add_4786_15_lut (.I0(GND_net), .I1(n12653[12]), .I2(n1026_adj_5113), 
            .I3(n40995), .O(n10645[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_15 (.CI(n40995), .I0(n12653[12]), .I1(n1026_adj_5113), 
            .CO(n40996));
    SB_LUT4 add_4786_14_lut (.I0(GND_net), .I1(n12653[11]), .I2(n953_adj_5114), 
            .I3(n40994), .O(n10645[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_14 (.CI(n40994), .I0(n12653[11]), .I1(n953_adj_5114), 
            .CO(n40995));
    SB_LUT4 add_4786_13_lut (.I0(GND_net), .I1(n12653[10]), .I2(n880_adj_5115), 
            .I3(n40993), .O(n10645[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_13 (.CI(n40993), .I0(n12653[10]), .I1(n880_adj_5115), 
            .CO(n40994));
    SB_LUT4 add_4786_12_lut (.I0(GND_net), .I1(n12653[9]), .I2(n807_adj_5116), 
            .I3(n40992), .O(n10645[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_12 (.CI(n40992), .I0(n12653[9]), .I1(n807_adj_5116), 
            .CO(n40993));
    SB_LUT4 add_4786_11_lut (.I0(GND_net), .I1(n12653[8]), .I2(n734_adj_5117), 
            .I3(n40991), .O(n10645[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_5062));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4786_11 (.CI(n40991), .I0(n12653[8]), .I1(n734_adj_5117), 
            .CO(n40992));
    SB_LUT4 add_4786_10_lut (.I0(GND_net), .I1(n12653[7]), .I2(n661_adj_5118), 
            .I3(n40990), .O(n10645[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_10 (.CI(n40990), .I0(n12653[7]), .I1(n661_adj_5118), 
            .CO(n40991));
    SB_LUT4 add_4786_9_lut (.I0(GND_net), .I1(n12653[6]), .I2(n588_adj_5119), 
            .I3(n40989), .O(n10645[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_9 (.CI(n40989), .I0(n12653[6]), .I1(n588_adj_5119), 
            .CO(n40990));
    SB_LUT4 add_4786_8_lut (.I0(GND_net), .I1(n12653[5]), .I2(n515_adj_5120), 
            .I3(n40988), .O(n10645[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_8 (.CI(n40988), .I0(n12653[5]), .I1(n515_adj_5120), 
            .CO(n40989));
    SB_LUT4 add_4786_7_lut (.I0(GND_net), .I1(n12653[4]), .I2(n442_adj_5121), 
            .I3(n40987), .O(n10645[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_7 (.CI(n40987), .I0(n12653[4]), .I1(n442_adj_5121), 
            .CO(n40988));
    SB_LUT4 add_4786_6_lut (.I0(GND_net), .I1(n12653[3]), .I2(n369_adj_5122), 
            .I3(n40986), .O(n10645[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_6 (.CI(n40986), .I0(n12653[3]), .I1(n369_adj_5122), 
            .CO(n40987));
    SB_LUT4 add_4786_5_lut (.I0(GND_net), .I1(n12653[2]), .I2(n296_adj_5123), 
            .I3(n40985), .O(n10645[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_5 (.CI(n40985), .I0(n12653[2]), .I1(n296_adj_5123), 
            .CO(n40986));
    SB_LUT4 add_4786_4_lut (.I0(GND_net), .I1(n12653[1]), .I2(n223_adj_5124), 
            .I3(n40984), .O(n10645[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_4 (.CI(n40984), .I0(n12653[1]), .I1(n223_adj_5124), 
            .CO(n40985));
    SB_LUT4 add_4786_3_lut (.I0(GND_net), .I1(n12653[0]), .I2(n150_adj_5125), 
            .I3(n40983), .O(n10645[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_3 (.CI(n40983), .I0(n12653[0]), .I1(n150_adj_5125), 
            .CO(n40984));
    SB_LUT4 add_4786_2_lut (.I0(GND_net), .I1(n8_adj_5126), .I2(n77_adj_5127), 
            .I3(GND_net), .O(n10645[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_2 (.CI(GND_net), .I0(n8_adj_5126), .I1(n77_adj_5127), 
            .CO(n40983));
    SB_LUT4 add_5749_22_lut (.I0(GND_net), .I1(n14231[19]), .I2(GND_net), 
            .I3(n40982), .O(n12653[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5749_21_lut (.I0(GND_net), .I1(n14231[18]), .I2(GND_net), 
            .I3(n40981), .O(n12653[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_21 (.CI(n40981), .I0(n14231[18]), .I1(GND_net), 
            .CO(n40982));
    SB_LUT4 add_5749_20_lut (.I0(GND_net), .I1(n14231[17]), .I2(GND_net), 
            .I3(n40980), .O(n12653[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_20 (.CI(n40980), .I0(n14231[17]), .I1(GND_net), 
            .CO(n40981));
    SB_LUT4 add_5749_19_lut (.I0(GND_net), .I1(n14231[16]), .I2(GND_net), 
            .I3(n40979), .O(n12653[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_19 (.CI(n40979), .I0(n14231[16]), .I1(GND_net), 
            .CO(n40980));
    SB_LUT4 add_5749_18_lut (.I0(GND_net), .I1(n14231[15]), .I2(GND_net), 
            .I3(n40978), .O(n12653[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_18 (.CI(n40978), .I0(n14231[15]), .I1(GND_net), 
            .CO(n40979));
    SB_LUT4 add_5749_17_lut (.I0(GND_net), .I1(n14231[14]), .I2(GND_net), 
            .I3(n40977), .O(n12653[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_17 (.CI(n40977), .I0(n14231[14]), .I1(GND_net), 
            .CO(n40978));
    SB_LUT4 add_5749_16_lut (.I0(GND_net), .I1(n14231[13]), .I2(n1102_adj_5128), 
            .I3(n40976), .O(n12653[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_16 (.CI(n40976), .I0(n14231[13]), .I1(n1102_adj_5128), 
            .CO(n40977));
    SB_LUT4 add_5749_15_lut (.I0(GND_net), .I1(n14231[12]), .I2(n1029_adj_5129), 
            .I3(n40975), .O(n12653[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_15 (.CI(n40975), .I0(n14231[12]), .I1(n1029_adj_5129), 
            .CO(n40976));
    SB_LUT4 add_5749_14_lut (.I0(GND_net), .I1(n14231[11]), .I2(n956_adj_5130), 
            .I3(n40974), .O(n12653[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_5061));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5749_14 (.CI(n40974), .I0(n14231[11]), .I1(n956_adj_5130), 
            .CO(n40975));
    SB_LUT4 add_5749_13_lut (.I0(GND_net), .I1(n14231[10]), .I2(n883_adj_5131), 
            .I3(n40973), .O(n12653[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_13 (.CI(n40973), .I0(n14231[10]), .I1(n883_adj_5131), 
            .CO(n40974));
    SB_LUT4 add_5749_12_lut (.I0(GND_net), .I1(n14231[9]), .I2(n810_adj_5132), 
            .I3(n40972), .O(n12653[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_12 (.CI(n40972), .I0(n14231[9]), .I1(n810_adj_5132), 
            .CO(n40973));
    SB_LUT4 add_5749_11_lut (.I0(GND_net), .I1(n14231[8]), .I2(n737_adj_5133), 
            .I3(n40971), .O(n12653[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_11 (.CI(n40971), .I0(n14231[8]), .I1(n737_adj_5133), 
            .CO(n40972));
    SB_LUT4 add_5749_10_lut (.I0(GND_net), .I1(n14231[7]), .I2(n664_adj_5134), 
            .I3(n40970), .O(n12653[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_10 (.CI(n40970), .I0(n14231[7]), .I1(n664_adj_5134), 
            .CO(n40971));
    SB_LUT4 add_5749_9_lut (.I0(GND_net), .I1(n14231[6]), .I2(n591_adj_5135), 
            .I3(n40969), .O(n12653[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_9 (.CI(n40969), .I0(n14231[6]), .I1(n591_adj_5135), 
            .CO(n40970));
    SB_LUT4 add_5749_8_lut (.I0(GND_net), .I1(n14231[5]), .I2(n518_adj_5136), 
            .I3(n40968), .O(n12653[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_8 (.CI(n40968), .I0(n14231[5]), .I1(n518_adj_5136), 
            .CO(n40969));
    SB_LUT4 add_5749_7_lut (.I0(GND_net), .I1(n14231[4]), .I2(n445_adj_5137), 
            .I3(n40967), .O(n12653[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_7 (.CI(n40967), .I0(n14231[4]), .I1(n445_adj_5137), 
            .CO(n40968));
    SB_LUT4 add_5749_6_lut (.I0(GND_net), .I1(n14231[3]), .I2(n372_adj_5138), 
            .I3(n40966), .O(n12653[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_6 (.CI(n40966), .I0(n14231[3]), .I1(n372_adj_5138), 
            .CO(n40967));
    SB_LUT4 add_5749_5_lut (.I0(GND_net), .I1(n14231[2]), .I2(n299_adj_5139), 
            .I3(n40965), .O(n12653[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_5 (.CI(n40965), .I0(n14231[2]), .I1(n299_adj_5139), 
            .CO(n40966));
    SB_LUT4 add_5749_4_lut (.I0(GND_net), .I1(n14231[1]), .I2(n226_adj_5140), 
            .I3(n40964), .O(n12653[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_4 (.CI(n40964), .I0(n14231[1]), .I1(n226_adj_5140), 
            .CO(n40965));
    SB_LUT4 add_5749_3_lut (.I0(GND_net), .I1(n14231[0]), .I2(n153_adj_5141), 
            .I3(n40963), .O(n12653[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_3 (.CI(n40963), .I0(n14231[0]), .I1(n153_adj_5141), 
            .CO(n40964));
    SB_LUT4 add_5749_2_lut (.I0(GND_net), .I1(n11_adj_5142), .I2(n80_adj_5143), 
            .I3(GND_net), .O(n12653[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5749_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5749_2 (.CI(GND_net), .I0(n11_adj_5142), .I1(n80_adj_5143), 
            .CO(n40963));
    SB_LUT4 add_6444_21_lut (.I0(GND_net), .I1(n15073[18]), .I2(GND_net), 
            .I3(n40962), .O(n14231[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6444_20_lut (.I0(GND_net), .I1(n15073[17]), .I2(GND_net), 
            .I3(n40961), .O(n14231[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_20 (.CI(n40961), .I0(n15073[17]), .I1(GND_net), 
            .CO(n40962));
    SB_LUT4 add_6444_19_lut (.I0(GND_net), .I1(n15073[16]), .I2(GND_net), 
            .I3(n40960), .O(n14231[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_19 (.CI(n40960), .I0(n15073[16]), .I1(GND_net), 
            .CO(n40961));
    SB_LUT4 add_6444_18_lut (.I0(GND_net), .I1(n15073[15]), .I2(GND_net), 
            .I3(n40959), .O(n14231[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_18 (.CI(n40959), .I0(n15073[15]), .I1(GND_net), 
            .CO(n40960));
    SB_LUT4 add_6444_17_lut (.I0(GND_net), .I1(n15073[14]), .I2(GND_net), 
            .I3(n40958), .O(n14231[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_17 (.CI(n40958), .I0(n15073[14]), .I1(GND_net), 
            .CO(n40959));
    SB_LUT4 add_6444_16_lut (.I0(GND_net), .I1(n15073[13]), .I2(n1105_adj_5144), 
            .I3(n40957), .O(n14231[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_16 (.CI(n40957), .I0(n15073[13]), .I1(n1105_adj_5144), 
            .CO(n40958));
    SB_LUT4 add_6444_15_lut (.I0(GND_net), .I1(n15073[12]), .I2(n1032_adj_5145), 
            .I3(n40956), .O(n14231[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_15 (.CI(n40956), .I0(n15073[12]), .I1(n1032_adj_5145), 
            .CO(n40957));
    SB_LUT4 add_6444_14_lut (.I0(GND_net), .I1(n15073[11]), .I2(n959_adj_5146), 
            .I3(n40955), .O(n14231[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_14 (.CI(n40955), .I0(n15073[11]), .I1(n959_adj_5146), 
            .CO(n40956));
    SB_LUT4 add_6444_13_lut (.I0(GND_net), .I1(n15073[10]), .I2(n886_adj_5147), 
            .I3(n40954), .O(n14231[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_13 (.CI(n40954), .I0(n15073[10]), .I1(n886_adj_5147), 
            .CO(n40955));
    SB_LUT4 add_6444_12_lut (.I0(GND_net), .I1(n15073[9]), .I2(n813_adj_5148), 
            .I3(n40953), .O(n14231[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_12 (.CI(n40953), .I0(n15073[9]), .I1(n813_adj_5148), 
            .CO(n40954));
    SB_LUT4 add_6444_11_lut (.I0(GND_net), .I1(n15073[8]), .I2(n740_adj_5149), 
            .I3(n40952), .O(n14231[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_11 (.CI(n40952), .I0(n15073[8]), .I1(n740_adj_5149), 
            .CO(n40953));
    SB_LUT4 add_6444_10_lut (.I0(GND_net), .I1(n15073[7]), .I2(n667_adj_5150), 
            .I3(n40951), .O(n14231[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n40679), .I0(GND_net), .I1(n1_adj_5153[3]), 
            .CO(n40680));
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_5060));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6444_10 (.CI(n40951), .I0(n15073[7]), .I1(n667_adj_5150), 
            .CO(n40952));
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_5059));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5058));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6444_9_lut (.I0(GND_net), .I1(n15073[6]), .I2(n594_adj_5105), 
            .I3(n40950), .O(n14231[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_9 (.CI(n40950), .I0(n15073[6]), .I1(n594_adj_5105), 
            .CO(n40951));
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_5057));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_5056));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6444_8_lut (.I0(GND_net), .I1(n15073[5]), .I2(n521_adj_5103), 
            .I3(n40949), .O(n14231[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[2]), 
            .I3(n40678), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_5055));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6444_8 (.CI(n40949), .I0(n15073[5]), .I1(n521_adj_5103), 
            .CO(n40950));
    SB_LUT4 add_6444_7_lut (.I0(GND_net), .I1(n15073[4]), .I2(n448_adj_5101), 
            .I3(n40948), .O(n14231[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_5054));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6444_7 (.CI(n40948), .I0(n15073[4]), .I1(n448_adj_5101), 
            .CO(n40949));
    SB_LUT4 add_6444_6_lut (.I0(GND_net), .I1(n15073[3]), .I2(n375_adj_5033), 
            .I3(n40947), .O(n14231[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n40678), .I0(GND_net), .I1(n1_adj_5153[2]), 
            .CO(n40679));
    SB_CARRY add_6444_6 (.CI(n40947), .I0(n15073[3]), .I1(n375_adj_5033), 
            .CO(n40948));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[1]), 
            .I3(n40677), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n40677), .I0(GND_net), .I1(n1_adj_5153[1]), 
            .CO(n40678));
    SB_LUT4 add_6444_5_lut (.I0(GND_net), .I1(n15073[2]), .I2(n302_adj_5031), 
            .I3(n40946), .O(n14231[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5153[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5153[0]), 
            .CO(n40677));
    SB_CARRY add_6444_5 (.CI(n40946), .I0(n15073[2]), .I1(n302_adj_5031), 
            .CO(n40947));
    SB_LUT4 add_6444_4_lut (.I0(GND_net), .I1(n15073[1]), .I2(n229_adj_5028), 
            .I3(n40945), .O(n14231[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_4 (.CI(n40945), .I0(n15073[1]), .I1(n229_adj_5028), 
            .CO(n40946));
    SB_LUT4 add_6444_3_lut (.I0(GND_net), .I1(n15073[0]), .I2(n156_adj_5019), 
            .I3(n40944), .O(n14231[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_3 (.CI(n40944), .I0(n15073[0]), .I1(n156_adj_5019), 
            .CO(n40945));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n40536), 
            .O(duty_23__N_3772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6444_2_lut (.I0(GND_net), .I1(n14_adj_5016), .I2(n83_adj_5007), 
            .I3(GND_net), .O(n14231[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6444_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n40676), .O(\PID_CONTROLLER.integral_23__N_3723 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6444_2 (.CI(GND_net), .I0(n14_adj_5016), .I1(n83_adj_5007), 
            .CO(n40944));
    SB_LUT4 add_6756_11_lut (.I0(GND_net), .I1(n19832[8]), .I2(n770_adj_5005), 
            .I3(n40943), .O(n19633[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6756_10_lut (.I0(GND_net), .I1(n19832[7]), .I2(n697_adj_5004), 
            .I3(n40942), .O(n19633[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_10 (.CI(n40942), .I0(n19832[7]), .I1(n697_adj_5004), 
            .CO(n40943));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n40675), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n40675), .I0(GND_net), .I1(n1[22]), 
            .CO(n40676));
    SB_CARRY add_12_11 (.CI(n40536), .I0(n106[9]), .I1(n155[9]), .CO(n40537));
    SB_LUT4 add_6756_9_lut (.I0(GND_net), .I1(n19832[6]), .I2(n624_adj_4999), 
            .I3(n40941), .O(n19633[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n40535), 
            .O(duty_23__N_3772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_9 (.CI(n40941), .I0(n19832[6]), .I1(n624_adj_4999), 
            .CO(n40942));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n40674), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6756_8_lut (.I0(GND_net), .I1(n19832[5]), .I2(n551_adj_4997), 
            .I3(n40940), .O(n19633[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_8 (.CI(n40940), .I0(n19832[5]), .I1(n551_adj_4997), 
            .CO(n40941));
    SB_LUT4 add_6756_7_lut (.I0(GND_net), .I1(n19832[4]), .I2(n478_adj_4996), 
            .I3(n40939), .O(n19633[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_7 (.CI(n40939), .I0(n19832[4]), .I1(n478_adj_4996), 
            .CO(n40940));
    SB_LUT4 add_6756_6_lut (.I0(GND_net), .I1(n19832[3]), .I2(n405_adj_4992), 
            .I3(n40938), .O(n19633[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_6 (.CI(n40938), .I0(n19832[3]), .I1(n405_adj_4992), 
            .CO(n40939));
    SB_LUT4 add_6756_5_lut (.I0(GND_net), .I1(n19832[2]), .I2(n332_adj_4991), 
            .I3(n40937), .O(n19633[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_5 (.CI(n40937), .I0(n19832[2]), .I1(n332_adj_4991), 
            .CO(n40938));
    SB_CARRY add_12_10 (.CI(n40535), .I0(n106[8]), .I1(n155[8]), .CO(n40536));
    SB_LUT4 add_6756_4_lut (.I0(GND_net), .I1(n19832[1]), .I2(n259_adj_4990), 
            .I3(n40936), .O(n19633[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_4 (.CI(n40936), .I0(n19832[1]), .I1(n259_adj_4990), 
            .CO(n40937));
    SB_LUT4 add_6756_3_lut (.I0(GND_net), .I1(n19832[0]), .I2(n186_adj_4988), 
            .I3(n40935), .O(n19633[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_3 (.CI(n40935), .I0(n19832[0]), .I1(n186_adj_4988), 
            .CO(n40936));
    SB_LUT4 add_6756_2_lut (.I0(GND_net), .I1(n44_adj_4987), .I2(n113_adj_4986), 
            .I3(GND_net), .O(n19633[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6756_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6756_2 (.CI(GND_net), .I0(n44_adj_4987), .I1(n113_adj_4986), 
            .CO(n40935));
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_5053));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6485_20_lut (.I0(GND_net), .I1(n15833[17]), .I2(GND_net), 
            .I3(n40934), .O(n15073[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_5052));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6485_19_lut (.I0(GND_net), .I1(n15833[16]), .I2(GND_net), 
            .I3(n40933), .O(n15073[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6746_11_lut (.I0(GND_net), .I1(n19733[8]), .I2(n770), 
            .I3(n40762), .O(n19513[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n40674), .I0(GND_net), .I1(n1[21]), 
            .CO(n40675));
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_5051));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_5050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6485_19 (.CI(n40933), .I0(n15833[16]), .I1(GND_net), 
            .CO(n40934));
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_5049));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6485_18_lut (.I0(GND_net), .I1(n15833[15]), .I2(GND_net), 
            .I3(n40932), .O(n15073[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_5048));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6485_18 (.CI(n40932), .I0(n15833[15]), .I1(GND_net), 
            .CO(n40933));
    SB_LUT4 add_6485_17_lut (.I0(GND_net), .I1(n15833[14]), .I2(GND_net), 
            .I3(n40931), .O(n15073[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_17 (.CI(n40931), .I0(n15833[14]), .I1(GND_net), 
            .CO(n40932));
    SB_LUT4 add_6485_16_lut (.I0(GND_net), .I1(n15833[13]), .I2(n1108_adj_4979), 
            .I3(n40930), .O(n15073[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_16 (.CI(n40930), .I0(n15833[13]), .I1(n1108_adj_4979), 
            .CO(n40931));
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6485_15_lut (.I0(GND_net), .I1(n15833[12]), .I2(n1035_adj_4978), 
            .I3(n40929), .O(n15073[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6746_10_lut (.I0(GND_net), .I1(n19733[7]), .I2(n697), 
            .I3(n40761), .O(n19513[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n40534), 
            .O(duty_23__N_3772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_15 (.CI(n40929), .I0(n15833[12]), .I1(n1035_adj_4978), 
            .CO(n40930));
    SB_LUT4 add_6485_14_lut (.I0(GND_net), .I1(n15833[11]), .I2(n962_adj_4972), 
            .I3(n40928), .O(n15073[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6746_10 (.CI(n40761), .I0(n19733[7]), .I1(n697), .CO(n40762));
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_5047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6485_14 (.CI(n40928), .I0(n15833[11]), .I1(n962_adj_4972), 
            .CO(n40929));
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_5046));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_5045));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6746_9_lut (.I0(GND_net), .I1(n19733[6]), .I2(n624), .I3(n40760), 
            .O(n19513[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6485_13_lut (.I0(GND_net), .I1(n15833[10]), .I2(n889_adj_4970), 
            .I3(n40927), .O(n15073[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_13 (.CI(n40927), .I0(n15833[10]), .I1(n889_adj_4970), 
            .CO(n40928));
    SB_LUT4 add_6485_12_lut (.I0(GND_net), .I1(n15833[9]), .I2(n816_adj_4962), 
            .I3(n40926), .O(n15073[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_12 (.CI(n40926), .I0(n15833[9]), .I1(n816_adj_4962), 
            .CO(n40927));
    SB_LUT4 add_6485_11_lut (.I0(GND_net), .I1(n15833[8]), .I2(n743_adj_4960), 
            .I3(n40925), .O(n15073[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_5044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6485_11 (.CI(n40925), .I0(n15833[8]), .I1(n743_adj_4960), 
            .CO(n40926));
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6485_10_lut (.I0(GND_net), .I1(n15833[7]), .I2(n670_adj_4959), 
            .I3(n40924), .O(n15073[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_10 (.CI(n40924), .I0(n15833[7]), .I1(n670_adj_4959), 
            .CO(n40925));
    SB_LUT4 add_6485_9_lut (.I0(GND_net), .I1(n15833[6]), .I2(n597_adj_4958), 
            .I3(n40923), .O(n15073[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n40673), .O(n41_adj_4774)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n40673), .I0(GND_net), .I1(n1[20]), 
            .CO(n40674));
    SB_CARRY add_6485_9 (.CI(n40923), .I0(n15833[6]), .I1(n597_adj_4958), 
            .CO(n40924));
    SB_LUT4 add_6485_8_lut (.I0(GND_net), .I1(n15833[5]), .I2(n524_adj_4952), 
            .I3(n40922), .O(n15073[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n40534), .I0(n106[7]), .I1(n155[7]), .CO(n40535));
    SB_CARRY add_6485_8 (.CI(n40922), .I0(n15833[5]), .I1(n524_adj_4952), 
            .CO(n40923));
    SB_LUT4 add_6485_7_lut (.I0(GND_net), .I1(n15833[4]), .I2(n451_adj_4951), 
            .I3(n40921), .O(n15073[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_7 (.CI(n40921), .I0(n15833[4]), .I1(n451_adj_4951), 
            .CO(n40922));
    SB_LUT4 add_6485_6_lut (.I0(GND_net), .I1(n15833[3]), .I2(n378_adj_4946), 
            .I3(n40920), .O(n15073[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_6 (.CI(n40920), .I0(n15833[3]), .I1(n378_adj_4946), 
            .CO(n40921));
    SB_LUT4 add_6485_5_lut (.I0(GND_net), .I1(n15833[2]), .I2(n305_adj_4939), 
            .I3(n40919), .O(n15073[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n40533), 
            .O(duty_23__N_3772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22149_2_lut (.I0(n34[13]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_8 (.CI(n40533), .I0(n106[6]), .I1(n155[6]), .CO(n40534));
    SB_CARRY add_6746_9 (.CI(n40760), .I0(n19733[6]), .I1(n624), .CO(n40761));
    SB_CARRY add_6485_5 (.CI(n40919), .I0(n15833[2]), .I1(n305_adj_4939), 
            .CO(n40920));
    SB_LUT4 add_6485_4_lut (.I0(GND_net), .I1(n15833[1]), .I2(n232_adj_4936), 
            .I3(n40918), .O(n15073[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_4 (.CI(n40918), .I0(n15833[1]), .I1(n232_adj_4936), 
            .CO(n40919));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n40672), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6485_3_lut (.I0(GND_net), .I1(n15833[0]), .I2(n159_adj_4934), 
            .I3(n40917), .O(n15073[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_3 (.CI(n40917), .I0(n15833[0]), .I1(n159_adj_4934), 
            .CO(n40918));
    SB_LUT4 add_6746_8_lut (.I0(GND_net), .I1(n19733[5]), .I2(n551), .I3(n40759), 
            .O(n19513[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6485_2_lut (.I0(GND_net), .I1(n17_adj_4933), .I2(n86_adj_4932), 
            .I3(GND_net), .O(n15073[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6485_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6485_2 (.CI(GND_net), .I0(n17_adj_4933), .I1(n86_adj_4932), 
            .CO(n40917));
    SB_LUT4 add_6522_19_lut (.I0(GND_net), .I1(n16517[16]), .I2(GND_net), 
            .I3(n40916), .O(n15833[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6522_18_lut (.I0(GND_net), .I1(n16517[15]), .I2(GND_net), 
            .I3(n40915), .O(n15833[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6746_8 (.CI(n40759), .I0(n19733[5]), .I1(n551), .CO(n40760));
    SB_CARRY add_6522_18 (.CI(n40915), .I0(n16517[15]), .I1(GND_net), 
            .CO(n40916));
    SB_LUT4 add_6522_17_lut (.I0(GND_net), .I1(n16517[14]), .I2(GND_net), 
            .I3(n40914), .O(n15833[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_17 (.CI(n40914), .I0(n16517[14]), .I1(GND_net), 
            .CO(n40915));
    SB_LUT4 add_6522_16_lut (.I0(GND_net), .I1(n16517[13]), .I2(n1111_adj_4931), 
            .I3(n40913), .O(n15833[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6746_7_lut (.I0(GND_net), .I1(n19733[4]), .I2(n478), .I3(n40758), 
            .O(n19513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35718_2_lut_4_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(duty_23__N_3772[9]), .I3(n257[9]), .O(n51352));
    defparam i35718_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6522_16 (.CI(n40913), .I0(n16517[13]), .I1(n1111_adj_4931), 
            .CO(n40914));
    SB_LUT4 add_6522_15_lut (.I0(GND_net), .I1(n16517[12]), .I2(n1038_adj_4930), 
            .I3(n40912), .O(n15833[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35731_2_lut_4_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(duty_23__N_3772[7]), .I3(n257[7]), .O(n51365));
    defparam i35731_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n40672), .I0(GND_net), .I1(n1[19]), 
            .CO(n40673));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n40532), 
            .O(duty_23__N_3772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_15 (.CI(n40912), .I0(n16517[12]), .I1(n1038_adj_4930), 
            .CO(n40913));
    SB_LUT4 add_6522_14_lut (.I0(GND_net), .I1(n16517[11]), .I2(n965_adj_4929), 
            .I3(n40911), .O(n15833[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_14 (.CI(n40911), .I0(n16517[11]), .I1(n965_adj_4929), 
            .CO(n40912));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n40671), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6746_7 (.CI(n40758), .I0(n19733[4]), .I1(n478), .CO(n40759));
    SB_LUT4 add_6746_6_lut (.I0(GND_net), .I1(n19733[3]), .I2(n405), .I3(n40757), 
            .O(n19513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n40671), .I0(GND_net), .I1(n1[18]), 
            .CO(n40672));
    SB_LUT4 add_6522_13_lut (.I0(GND_net), .I1(n16517[10]), .I2(n892_adj_4927), 
            .I3(n40910), .O(n15833[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_13 (.CI(n40910), .I0(n16517[10]), .I1(n892_adj_4927), 
            .CO(n40911));
    SB_LUT4 add_6522_12_lut (.I0(GND_net), .I1(n16517[9]), .I2(n819_adj_4926), 
            .I3(n40909), .O(n15833[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_12 (.CI(n40909), .I0(n16517[9]), .I1(n819_adj_4926), 
            .CO(n40910));
    SB_LUT4 add_6522_11_lut (.I0(GND_net), .I1(n16517[8]), .I2(n746_adj_4925), 
            .I3(n40908), .O(n15833[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_11 (.CI(n40908), .I0(n16517[8]), .I1(n746_adj_4925), 
            .CO(n40909));
    SB_LUT4 add_6522_10_lut (.I0(GND_net), .I1(n16517[7]), .I2(n673_adj_4921), 
            .I3(n40907), .O(n15833[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_10 (.CI(n40907), .I0(n16517[7]), .I1(n673_adj_4921), 
            .CO(n40908));
    SB_CARRY add_6746_6 (.CI(n40757), .I0(n19733[3]), .I1(n405), .CO(n40758));
    SB_LUT4 add_6522_9_lut (.I0(GND_net), .I1(n16517[6]), .I2(n600_adj_4920), 
            .I3(n40906), .O(n15833[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6746_5_lut (.I0(GND_net), .I1(n19733[2]), .I2(n332), .I3(n40756), 
            .O(n19513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_9 (.CI(n40906), .I0(n16517[6]), .I1(n600_adj_4920), 
            .CO(n40907));
    SB_CARRY add_6746_5 (.CI(n40756), .I0(n19733[2]), .I1(n332), .CO(n40757));
    SB_LUT4 add_6522_8_lut (.I0(GND_net), .I1(n16517[5]), .I2(n527_adj_4913), 
            .I3(n40905), .O(n15833[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_8 (.CI(n40905), .I0(n16517[5]), .I1(n527_adj_4913), 
            .CO(n40906));
    SB_LUT4 add_6522_7_lut (.I0(GND_net), .I1(n16517[4]), .I2(n454_adj_4912), 
            .I3(n40904), .O(n15833[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_7 (.CI(n40904), .I0(n16517[4]), .I1(n454_adj_4912), 
            .CO(n40905));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n40670), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n40670), .I0(GND_net), .I1(n1[17]), 
            .CO(n40671));
    SB_LUT4 add_6522_6_lut (.I0(GND_net), .I1(n16517[3]), .I2(n381_adj_4908), 
            .I3(n40903), .O(n15833[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_6 (.CI(n40903), .I0(n16517[3]), .I1(n381_adj_4908), 
            .CO(n40904));
    SB_LUT4 add_6522_5_lut (.I0(GND_net), .I1(n16517[2]), .I2(n308_adj_4907), 
            .I3(n40902), .O(n15833[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35755_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3772[9]), .O(n51389));
    defparam i35755_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i35768_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3772[7]), .O(n51402));
    defparam i35768_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_6522_5 (.CI(n40902), .I0(n16517[2]), .I1(n308_adj_4907), 
            .CO(n40903));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n40669), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6522_4_lut (.I0(GND_net), .I1(n16517[1]), .I2(n235_adj_4900), 
            .I3(n40901), .O(n15833[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_4 (.CI(n40901), .I0(n16517[1]), .I1(n235_adj_4900), 
            .CO(n40902));
    SB_LUT4 i22148_2_lut (.I0(n34[14]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6746_4_lut (.I0(GND_net), .I1(n19733[1]), .I2(n259), .I3(n40755), 
            .O(n19513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6522_3_lut (.I0(GND_net), .I1(n16517[0]), .I2(n162_adj_4894), 
            .I3(n40900), .O(n15833[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_3 (.CI(n40900), .I0(n16517[0]), .I1(n162_adj_4894), 
            .CO(n40901));
    SB_LUT4 add_6522_2_lut (.I0(GND_net), .I1(n20_adj_4893), .I2(n89_adj_4892), 
            .I3(GND_net), .O(n15833[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_2 (.CI(GND_net), .I0(n20_adj_4893), .I1(n89_adj_4892), 
            .CO(n40900));
    SB_LUT4 add_6774_10_lut (.I0(GND_net), .I1(n19993[7]), .I2(n700_adj_4890), 
            .I3(n40899), .O(n19832[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6774_9_lut (.I0(GND_net), .I1(n19993[6]), .I2(n627_adj_4885), 
            .I3(n40898), .O(n19832[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_9 (.CI(n40898), .I0(n19993[6]), .I1(n627_adj_4885), 
            .CO(n40899));
    SB_LUT4 add_6774_8_lut (.I0(GND_net), .I1(n19993[5]), .I2(n554_adj_4884), 
            .I3(n40897), .O(n19832[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_8 (.CI(n40897), .I0(n19993[5]), .I1(n554_adj_4884), 
            .CO(n40898));
    SB_LUT4 add_6774_7_lut (.I0(GND_net), .I1(n19993[4]), .I2(n481_adj_4883), 
            .I3(n40896), .O(n19832[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n40669), .I0(GND_net), .I1(n1[16]), 
            .CO(n40670));
    SB_CARRY add_6774_7 (.CI(n40896), .I0(n19993[4]), .I1(n481_adj_4883), 
            .CO(n40897));
    SB_LUT4 add_6774_6_lut (.I0(GND_net), .I1(n19993[3]), .I2(n408_adj_4882), 
            .I3(n40895), .O(n19832[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_6 (.CI(n40895), .I0(n19993[3]), .I1(n408_adj_4882), 
            .CO(n40896));
    SB_LUT4 add_6774_5_lut (.I0(GND_net), .I1(n19993[2]), .I2(n335_adj_4881), 
            .I3(n40894), .O(n19832[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_5 (.CI(n40894), .I0(n19993[2]), .I1(n335_adj_4881), 
            .CO(n40895));
    SB_LUT4 add_6774_4_lut (.I0(GND_net), .I1(n19993[1]), .I2(n262_adj_4880), 
            .I3(n40893), .O(n19832[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_4 (.CI(n40893), .I0(n19993[1]), .I1(n262_adj_4880), 
            .CO(n40894));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n40668), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6774_3_lut (.I0(GND_net), .I1(n19993[0]), .I2(n189_adj_4878), 
            .I3(n40892), .O(n19832[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_3 (.CI(n40892), .I0(n19993[0]), .I1(n189_adj_4878), 
            .CO(n40893));
    SB_LUT4 add_6774_2_lut (.I0(GND_net), .I1(n47_adj_4877), .I2(n116_adj_4876), 
            .I3(GND_net), .O(n19832[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6774_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6774_2 (.CI(GND_net), .I0(n47_adj_4877), .I1(n116_adj_4876), 
            .CO(n40892));
    SB_LUT4 add_6557_18_lut (.I0(GND_net), .I1(n17129[15]), .I2(GND_net), 
            .I3(n40891), .O(n16517[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6557_17_lut (.I0(GND_net), .I1(n17129[14]), .I2(GND_net), 
            .I3(n40890), .O(n16517[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6746_4 (.CI(n40755), .I0(n19733[1]), .I1(n259), .CO(n40756));
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4982));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6557_17 (.CI(n40890), .I0(n17129[14]), .I1(GND_net), 
            .CO(n40891));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n40668), .I0(GND_net), .I1(n1[15]), 
            .CO(n40669));
    SB_LUT4 add_6557_16_lut (.I0(GND_net), .I1(n17129[13]), .I2(n1114), 
            .I3(n40889), .O(n16517[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_16 (.CI(n40889), .I0(n17129[13]), .I1(n1114), .CO(n40890));
    SB_LUT4 add_6746_3_lut (.I0(GND_net), .I1(n19733[0]), .I2(n186), .I3(n40754), 
            .O(n19513[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6557_15_lut (.I0(GND_net), .I1(n17129[12]), .I2(n1041), 
            .I3(n40888), .O(n16517[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_15 (.CI(n40888), .I0(n17129[12]), .I1(n1041), .CO(n40889));
    SB_LUT4 add_6557_14_lut (.I0(GND_net), .I1(n17129[11]), .I2(n968), 
            .I3(n40887), .O(n16517[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_14 (.CI(n40887), .I0(n17129[11]), .I1(n968), .CO(n40888));
    SB_LUT4 add_6557_13_lut (.I0(GND_net), .I1(n17129[10]), .I2(n895), 
            .I3(n40886), .O(n16517[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_13 (.CI(n40886), .I0(n17129[10]), .I1(n895), .CO(n40887));
    SB_LUT4 add_6557_12_lut (.I0(GND_net), .I1(n17129[9]), .I2(n822), 
            .I3(n40885), .O(n16517[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_12 (.CI(n40885), .I0(n17129[9]), .I1(n822), .CO(n40886));
    SB_LUT4 add_6557_11_lut (.I0(GND_net), .I1(n17129[8]), .I2(n749), 
            .I3(n40884), .O(n16517[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_11 (.CI(n40884), .I0(n17129[8]), .I1(n749), .CO(n40885));
    SB_LUT4 add_6557_10_lut (.I0(GND_net), .I1(n17129[7]), .I2(n676), 
            .I3(n40883), .O(n16517[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_10 (.CI(n40883), .I0(n17129[7]), .I1(n676), .CO(n40884));
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4981));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6557_9_lut (.I0(GND_net), .I1(n17129[6]), .I2(n603), .I3(n40882), 
            .O(n16517[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6746_3 (.CI(n40754), .I0(n19733[0]), .I1(n186), .CO(n40755));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n40667), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6557_9 (.CI(n40882), .I0(n17129[6]), .I1(n603), .CO(n40883));
    SB_LUT4 add_6557_8_lut (.I0(GND_net), .I1(n17129[5]), .I2(n530), .I3(n40881), 
            .O(n16517[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n40667), .I0(GND_net), .I1(n1[14]), 
            .CO(n40668));
    SB_CARRY add_6557_8 (.CI(n40881), .I0(n17129[5]), .I1(n530), .CO(n40882));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n40666), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6557_7_lut (.I0(GND_net), .I1(n17129[4]), .I2(n457), .I3(n40880), 
            .O(n16517[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_7 (.CI(n40880), .I0(n17129[4]), .I1(n457), .CO(n40881));
    SB_LUT4 add_6557_6_lut (.I0(GND_net), .I1(n17129[3]), .I2(n384), .I3(n40879), 
            .O(n16517[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_6 (.CI(n40879), .I0(n17129[3]), .I1(n384), .CO(n40880));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n40666), .I0(GND_net), .I1(n1[13]), 
            .CO(n40667));
    SB_LUT4 add_6557_5_lut (.I0(GND_net), .I1(n17129[2]), .I2(n311), .I3(n40878), 
            .O(n16517[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_5 (.CI(n40878), .I0(n17129[2]), .I1(n311), .CO(n40879));
    SB_LUT4 add_6557_4_lut (.I0(GND_net), .I1(n17129[1]), .I2(n238), .I3(n40877), 
            .O(n16517[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_4 (.CI(n40877), .I0(n17129[1]), .I1(n238), .CO(n40878));
    SB_LUT4 add_6557_3_lut (.I0(GND_net), .I1(n17129[0]), .I2(n165), .I3(n40876), 
            .O(n16517[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6746_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19513[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6746_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6557_3 (.CI(n40876), .I0(n17129[0]), .I1(n165), .CO(n40877));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n40665), .O(n25_adj_4751)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_7 (.CI(n40532), .I0(n106[5]), .I1(n155[5]), .CO(n40533));
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6557_2_lut (.I0(GND_net), .I1(n23_adj_4869), .I2(n92), 
            .I3(GND_net), .O(n16517[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6557_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4967));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4961));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6557_2 (.CI(GND_net), .I0(n23_adj_4869), .I1(n92), .CO(n40876));
    SB_LUT4 add_6590_17_lut (.I0(GND_net), .I1(n17673[14]), .I2(GND_net), 
            .I3(n40875), .O(n17129[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6590_16_lut (.I0(GND_net), .I1(n17673[13]), .I2(n1117), 
            .I3(n40874), .O(n17129[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n40665), .I0(GND_net), .I1(n1[12]), 
            .CO(n40666));
    SB_CARRY add_6746_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n40754));
    SB_CARRY add_6590_16 (.CI(n40874), .I0(n17673[13]), .I1(n1117), .CO(n40875));
    SB_LUT4 add_6765_10_lut (.I0(GND_net), .I1(n19913[7]), .I2(n700), 
            .I3(n40753), .O(n19733[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6590_15_lut (.I0(GND_net), .I1(n17673[12]), .I2(n1044), 
            .I3(n40873), .O(n17129[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_15 (.CI(n40873), .I0(n17673[12]), .I1(n1044), .CO(n40874));
    SB_LUT4 add_6590_14_lut (.I0(GND_net), .I1(n17673[11]), .I2(n971), 
            .I3(n40872), .O(n17129[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6765_9_lut (.I0(GND_net), .I1(n19913[6]), .I2(n627), .I3(n40752), 
            .O(n19733[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_14 (.CI(n40872), .I0(n17673[11]), .I1(n971), .CO(n40873));
    SB_LUT4 add_6590_13_lut (.I0(GND_net), .I1(n17673[10]), .I2(n898), 
            .I3(n40871), .O(n17129[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_13 (.CI(n40871), .I0(n17673[10]), .I1(n898), .CO(n40872));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n40664), .O(n23_adj_4752)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4945));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6590_12_lut (.I0(GND_net), .I1(n17673[9]), .I2(n825), 
            .I3(n40870), .O(n17129[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_12 (.CI(n40870), .I0(n17673[9]), .I1(n825), .CO(n40871));
    SB_LUT4 add_6590_11_lut (.I0(GND_net), .I1(n17673[8]), .I2(n752), 
            .I3(n40869), .O(n17129[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6765_9 (.CI(n40752), .I0(n19913[6]), .I1(n627), .CO(n40753));
    SB_CARRY add_6590_11 (.CI(n40869), .I0(n17673[8]), .I1(n752), .CO(n40870));
    SB_LUT4 add_6590_10_lut (.I0(GND_net), .I1(n17673[7]), .I2(n679), 
            .I3(n40868), .O(n17129[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_10 (.CI(n40868), .I0(n17673[7]), .I1(n679), .CO(n40869));
    SB_LUT4 add_6590_9_lut (.I0(GND_net), .I1(n17673[6]), .I2(n606), .I3(n40867), 
            .O(n17129[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6765_8_lut (.I0(GND_net), .I1(n19913[5]), .I2(n554), .I3(n40751), 
            .O(n19733[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n40531), 
            .O(duty_23__N_3772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26595_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[21]), .I2(n34[20]), 
            .I3(\Kp[1] ), .O(n20368[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26595_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n40664), .I0(GND_net), .I1(n1[11]), 
            .CO(n40665));
    SB_CARRY add_6590_9 (.CI(n40867), .I0(n17673[6]), .I1(n606), .CO(n40868));
    SB_CARRY add_12_6 (.CI(n40531), .I0(n106[4]), .I1(n155[4]), .CO(n40532));
    SB_LUT4 add_6590_8_lut (.I0(GND_net), .I1(n17673[5]), .I2(n533), .I3(n40866), 
            .O(n17129[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n40530), 
            .O(duty_23__N_3772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4924));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_5 (.CI(n40530), .I0(n106[3]), .I1(n155[3]), .CO(n40531));
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4923));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4922));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6590_8 (.CI(n40866), .I0(n17673[5]), .I1(n533), .CO(n40867));
    SB_LUT4 i26597_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[21]), .I2(n34[20]), 
            .I3(\Kp[1] ), .O(n40268));   // verilog/motorControl.v(34[16:22])
    defparam i26597_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_6590_7_lut (.I0(GND_net), .I1(n17673[4]), .I2(n460), .I3(n40865), 
            .O(n17129[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_7 (.CI(n40865), .I0(n17673[4]), .I1(n460), .CO(n40866));
    SB_LUT4 add_6590_6_lut (.I0(GND_net), .I1(n17673[3]), .I2(n387), .I3(n40864), 
            .O(n17129[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4919));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6590_6 (.CI(n40864), .I0(n17673[3]), .I1(n387), .CO(n40865));
    SB_LUT4 add_6590_5_lut (.I0(GND_net), .I1(n17673[2]), .I2(n314), .I3(n40863), 
            .O(n17129[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_5 (.CI(n40863), .I0(n17673[2]), .I1(n314), .CO(n40864));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n40529), 
            .O(duty_23__N_3772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4918));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6590_4_lut (.I0(GND_net), .I1(n17673[1]), .I2(n241), .I3(n40862), 
            .O(n17129[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_4 (.CI(n40862), .I0(n17673[1]), .I1(n241), .CO(n40863));
    SB_LUT4 add_6590_3_lut (.I0(GND_net), .I1(n17673[0]), .I2(n168), .I3(n40861), 
            .O(n17129[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_3 (.CI(n40861), .I0(n17673[0]), .I1(n168), .CO(n40862));
    SB_LUT4 add_6590_2_lut (.I0(GND_net), .I1(n26_adj_4865), .I2(n95), 
            .I3(GND_net), .O(n17129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6590_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6590_2 (.CI(GND_net), .I0(n26_adj_4865), .I1(n95), .CO(n40861));
    SB_LUT4 add_6790_9_lut (.I0(GND_net), .I1(n20120[6]), .I2(n630_adj_4863), 
            .I3(n40860), .O(n19993[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6790_8_lut (.I0(GND_net), .I1(n20120[5]), .I2(n557_adj_4862), 
            .I3(n40859), .O(n19993[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6790_8 (.CI(n40859), .I0(n20120[5]), .I1(n557_adj_4862), 
            .CO(n40860));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n40663), .O(n21_adj_4745)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6790_7_lut (.I0(GND_net), .I1(n20120[4]), .I2(n484_adj_4860), 
            .I3(n40858), .O(n19993[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6790_7 (.CI(n40858), .I0(n20120[4]), .I1(n484_adj_4860), 
            .CO(n40859));
    SB_LUT4 add_6790_6_lut (.I0(GND_net), .I1(n20120[3]), .I2(n411_adj_4859), 
            .I3(n40857), .O(n19993[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6790_6 (.CI(n40857), .I0(n20120[3]), .I1(n411_adj_4859), 
            .CO(n40858));
    SB_LUT4 add_6790_5_lut (.I0(GND_net), .I1(n20120[2]), .I2(n338_adj_4858), 
            .I3(n40856), .O(n19993[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n40663), .I0(GND_net), .I1(n1[10]), 
            .CO(n40664));
    SB_CARRY add_6790_5 (.CI(n40856), .I0(n20120[2]), .I1(n338_adj_4858), 
            .CO(n40857));
    SB_CARRY add_12_4 (.CI(n40529), .I0(n106[2]), .I1(n155[2]), .CO(n40530));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n40662), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6790_4_lut (.I0(GND_net), .I1(n20120[1]), .I2(n265_adj_4856), 
            .I3(n40855), .O(n19993[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6790_4 (.CI(n40855), .I0(n20120[1]), .I1(n265_adj_4856), 
            .CO(n40856));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n40662), .I0(GND_net), .I1(n1[9]), 
            .CO(n40663));
    SB_LUT4 add_6790_3_lut (.I0(GND_net), .I1(n20120[0]), .I2(n192_adj_4854), 
            .I3(n40854), .O(n19993[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6790_3 (.CI(n40854), .I0(n20120[0]), .I1(n192_adj_4854), 
            .CO(n40855));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n40661), .O(n17_adj_4746)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n40528), 
            .O(duty_23__N_3772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6765_8 (.CI(n40751), .I0(n19913[5]), .I1(n554), .CO(n40752));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n40661), .I0(GND_net), .I1(n1[8]), 
            .CO(n40662));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n40660), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6790_2_lut (.I0(GND_net), .I1(n50_adj_4849), .I2(n119_adj_4848), 
            .I3(GND_net), .O(n19993[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6790_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n40660), .I0(GND_net), .I1(n1[7]), 
            .CO(n40661));
    SB_CARRY add_6790_2 (.CI(GND_net), .I0(n50_adj_4849), .I1(n119_adj_4848), 
            .CO(n40854));
    SB_LUT4 add_6765_7_lut (.I0(GND_net), .I1(n19913[4]), .I2(n481), .I3(n40750), 
            .O(n19733[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n40659), .O(n13_adj_4743)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6765_7 (.CI(n40750), .I0(n19913[4]), .I1(n481), .CO(n40751));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n40659), .I0(GND_net), .I1(n1[6]), 
            .CO(n40660));
    SB_LUT4 add_6621_16_lut (.I0(GND_net), .I1(n18153[13]), .I2(n1120), 
            .I3(n40853), .O(n17673[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6621_15_lut (.I0(GND_net), .I1(n18153[12]), .I2(n1047), 
            .I3(n40852), .O(n17673[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6621_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6765_6_lut (.I0(GND_net), .I1(n19913[3]), .I2(n408), .I3(n40749), 
            .O(n19733[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n40658), .O(n11_adj_4744)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_12_3 (.CI(n40528), .I0(n106[1]), .I1(n155[1]), .CO(n40529));
    SB_CARRY add_6765_6 (.CI(n40749), .I0(n19913[3]), .I1(n408), .CO(n40750));
    SB_CARRY add_6621_15 (.CI(n40852), .I0(n18153[12]), .I1(n1047), .CO(n40853));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n40658), .I0(GND_net), .I1(n1[5]), 
            .CO(n40659));
    SB_LUT4 add_6765_5_lut (.I0(GND_net), .I1(n19913[2]), .I2(n335), .I3(n40748), 
            .O(n19733[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6765_5 (.CI(n40748), .I0(n19913[2]), .I1(n335), .CO(n40749));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n40657), .O(n9_adj_4747)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6765_4_lut (.I0(GND_net), .I1(n19913[1]), .I2(n262), .I3(n40747), 
            .O(n19733[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6765_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26678_3_lut_4_lut (.I0(\Kp[4] ), .I1(n34[18]), .I2(n6_adj_5151), 
            .I3(n20337[2]), .O(n8_adj_4802));   // verilog/motorControl.v(34[16:22])
    defparam i26678_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(\Kp[4] ), .I1(n34[18]), .I2(n20337[2]), 
            .I3(n6_adj_5151), .O(n20288[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h8778;
    SB_LUT4 i26670_3_lut_4_lut (.I0(\Kp[3] ), .I1(n34[18]), .I2(n4_adj_5152), 
            .I3(n20337[1]), .O(n6_adj_5151));   // verilog/motorControl.v(34[16:22])
    defparam i26670_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_5150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_5149));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1523 (.I0(\Kp[3] ), .I1(n34[18]), .I2(n20337[1]), 
            .I3(n4_adj_5152), .O(n20288[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1523.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_5148));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_5147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_5146));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_5145));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_5144));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1524 (.I0(\Kp[2] ), .I1(n34[19]), .I2(n20368[0]), 
            .I3(n40293), .O(n20337[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1524.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_5143));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5142));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_5141));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_5140));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_5139));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_5138));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_5137));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_5136));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_5135));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_5134));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26631_3_lut_4_lut (.I0(\Kp[2] ), .I1(n34[19]), .I2(n40293), 
            .I3(n20368[0]), .O(n4_adj_4797));   // verilog/motorControl.v(34[16:22])
    defparam i26631_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_5133));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_5132));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26618_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[20]), .I2(n34[19]), 
            .I3(\Kp[1] ), .O(n20337[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26618_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_5131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_5130));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_5129));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_5128));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_5127));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5126));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26620_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[20]), .I2(n34[19]), 
            .I3(\Kp[1] ), .O(n40293));   // verilog/motorControl.v(34[16:22])
    defparam i26620_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_5125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_5124));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_5123));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5121));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26487_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n20353[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26487_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_5120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_5119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_5118));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_5115));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_5114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_5113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22147_2_lut (.I0(n34[15]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22147_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4917));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4916));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4915));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_5112));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4914));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\Kp[2] ), .I1(n34[18]), .I2(n20337[0]), 
            .I3(n40327), .O(n20288[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h8778;
    SB_LUT4 i26662_3_lut_4_lut (.I0(\Kp[2] ), .I1(n34[18]), .I2(n40327), 
            .I3(n20337[0]), .O(n4_adj_5152));   // verilog/motorControl.v(34[16:22])
    defparam i26662_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4909));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4906));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26649_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[19]), .I2(n34[18]), 
            .I3(\Kp[1] ), .O(n20288[0]));   // verilog/motorControl.v(34[16:22])
    defparam i26649_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4905));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4903));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4902));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26651_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n34[19]), .I2(n34[18]), 
            .I3(\Kp[1] ), .O(n40327));   // verilog/motorControl.v(34[16:22])
    defparam i26651_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4899));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4897));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4896));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4891));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4888));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4887));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3772[1]), .I1(n257[1]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3747[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3772[2]), .I1(n257[2]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3747[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3747[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3747[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26489_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n40150));   // verilog/motorControl.v(34[25:36])
    defparam i26489_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3747[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3747[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3747[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3747[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3747[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3747[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3747[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3747[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3747[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3747[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3747[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3747[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3747[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3747[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3747[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3747[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3747[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3747[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3772[23]), .I1(n257[23]), .I2(n256_adj_5043), 
            .I3(GND_net), .O(duty_23__N_3747[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3747[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22146_2_lut (.I0(n34[16]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4873));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4765));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5153[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4872));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4871));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26577_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n4_adj_4736), .I3(n20313[1]), .O(n6));   // verilog/motorControl.v(34[25:36])
    defparam i26577_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1526 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n20313[1]), .I3(n4_adj_4736), .O(n20253[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1526.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22145_2_lut (.I0(n34[17]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22145_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4867));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4866));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22144_2_lut (.I0(n34[18]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4864));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1527 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n20313[0]), .I3(n40225), .O(n20253[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1527.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22143_2_lut (.I0(n34[19]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4230[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i22143_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4855));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26525_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n20313[0]));   // verilog/motorControl.v(34[25:36])
    defparam i26525_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4853));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4852));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1528 (.I0(n6), .I1(\Ki[4] ), .I2(n20313[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n20253[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1528.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n34[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (reg_B, CLK_c, n48368, data_i, n30744, 
            data_o, n30743, n30123, GND_net, VCC_net);
    output [2:0]reg_B;
    input CLK_c;
    output n48368;
    input [2:0]data_i;
    input n30744;
    output [2:0]data_o;
    input n30743;
    input n30123;
    input GND_net;
    input VCC_net;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n16, n17, n6, cnt_next_9__N_812;
    wire [9:0]n45;
    
    wire n41801, n41800, n41799, n41798, n41797, n41796, n41795, 
        n41794, n41793;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[3]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[9]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[5]), .I2(n16), .I3(cnt_reg[6]), 
            .O(n48368));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(reg_B[1]), .I2(reg_A[0]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n48368), .I1(n6), .I2(reg_B[2]), .I3(reg_A[2]), 
            .O(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdffd;
    SB_DFFSR cnt_reg_2190__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n30744));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n30743));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_2190__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2190__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n30123));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 cnt_reg_2190_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n41801), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2190_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n41800), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_10 (.CI(n41800), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n41801));
    SB_LUT4 cnt_reg_2190_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n41799), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_9 (.CI(n41799), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n41800));
    SB_LUT4 cnt_reg_2190_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n41798), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_8 (.CI(n41798), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n41799));
    SB_LUT4 cnt_reg_2190_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n41797), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_7 (.CI(n41797), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n41798));
    SB_LUT4 cnt_reg_2190_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n41796), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_6 (.CI(n41796), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n41797));
    SB_LUT4 cnt_reg_2190_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n41795), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_5 (.CI(n41795), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n41796));
    SB_LUT4 cnt_reg_2190_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n41794), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_4 (.CI(n41794), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n41795));
    SB_LUT4 cnt_reg_2190_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n41793), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_3 (.CI(n41793), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n41794));
    SB_LUT4 cnt_reg_2190_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2190_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2190_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n41793));
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (\state[3] , n6, GND_net, CLK_c, n5608, \state[1] , 
            read, \state[0] , enable_slow_N_4190, \state[1]_adj_18 , 
            \state[2] , n7, n30170, rw, n45294, data_ready, n45186, 
            n45170, n36514, n46391, n45666, \state_7__N_4087[0] , 
            sda_enable, n4, scl_enable_N_4177, scl_enable, n6686, 
            n35782, n8, VCC_net, \state[0]_adj_19 , n4_adj_20, \saved_addr[0] , 
            n6496, n51120, n15, n10, n28421, n28416, n10_adj_21, 
            \state_7__N_4103[3] , n7227, n30174, n30159, data, n30158, 
            n30157, n30146, scl, sda_out, n30138, n30137, n30136, 
            n30135, n10_adj_22) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[3] ;
    output n6;
    input GND_net;
    input CLK_c;
    output [0:0]n5608;
    output \state[1] ;
    input read;
    output \state[0] ;
    input enable_slow_N_4190;
    output \state[1]_adj_18 ;
    output \state[2] ;
    output n7;
    input n30170;
    output rw;
    input n45294;
    output data_ready;
    input n45186;
    input n45170;
    output n36514;
    input n46391;
    output n45666;
    output \state_7__N_4087[0] ;
    output sda_enable;
    output n4;
    input scl_enable_N_4177;
    output scl_enable;
    output n6686;
    output n35782;
    input n8;
    input VCC_net;
    output \state[0]_adj_19 ;
    output n4_adj_20;
    output \saved_addr[0] ;
    input n6496;
    output n51120;
    output n15;
    output n10;
    output n28421;
    output n28416;
    output n10_adj_21;
    input \state_7__N_4103[3] ;
    input n7227;
    input n30174;
    input n30159;
    output [7:0]data;
    input n30158;
    input n30157;
    input n30146;
    output scl;
    output sda_out;
    input n30138;
    input n30137;
    input n30136;
    input n30135;
    input n10_adj_22;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n40585;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    wire [15:0]n4266;
    
    wire n40586, n28277;
    wire [15:0]delay_counter_15__N_3989;
    
    wire n29743, n30036, enable, n28, n26, n27, n25, n40599, 
        n40598, n40597, n40596, n40595, n40594, n40593, n40592, 
        n40591, n40590, n40589, n40588, n40587;
    
    SB_CARRY add_961_3 (.CI(n40585), .I0(delay_counter[1]), .I1(n4266[15]), 
            .CO(n40586));
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n28277), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[1]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[2]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[3]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[4]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[5]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[6]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[7]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[8]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[9]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[10]), .S(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[11]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[12]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[13]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[14]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[15]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_961_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4266[15]), 
            .I3(GND_net), .O(delay_counter_15__N_3989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4266[15]), 
            .CO(n40585));
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n5608[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 mux_1409_Mux_0_i1_4_lut (.I0(read), .I1(n28277), .I2(\state[0] ), 
            .I3(enable_slow_N_4190), .O(n5608[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1409_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n29743), 
            .D(delay_counter_15__N_3989[0]), .R(n30036));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut_adj_1514 (.I0(\state[1]_adj_18 ), .I1(\state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_1514.LUT_INIT = 16'heeee;
    SB_LUT4 i16360_2_lut (.I0(n29743), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n30036));   // verilog/eeprom.v(26[8] 58[4])
    defparam i16360_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n29743));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n30170));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n45294));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n28277));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36419_2_lut (.I0(n28277), .I1(enable_slow_N_4190), .I2(GND_net), 
            .I3(GND_net), .O(n4266[15]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i36419_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_961_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4266[15]), 
            .I3(n40599), .O(delay_counter_15__N_3989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_961_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4266[15]), 
            .I3(n40598), .O(delay_counter_15__N_3989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n45186));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n45170));   // verilog/eeprom.v(26[8] 58[4])
    SB_CARRY add_961_16 (.CI(n40598), .I0(delay_counter[14]), .I1(n4266[15]), 
            .CO(n40599));
    SB_LUT4 add_961_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4266[15]), 
            .I3(n40597), .O(delay_counter_15__N_3989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_15 (.CI(n40597), .I0(delay_counter[13]), .I1(n4266[15]), 
            .CO(n40598));
    SB_LUT4 add_961_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4266[15]), 
            .I3(n40596), .O(delay_counter_15__N_3989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_14 (.CI(n40596), .I0(delay_counter[12]), .I1(n4266[15]), 
            .CO(n40597));
    SB_LUT4 add_961_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4266[15]), 
            .I3(n40595), .O(delay_counter_15__N_3989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_13 (.CI(n40595), .I0(delay_counter[11]), .I1(n4266[15]), 
            .CO(n40596));
    SB_LUT4 add_961_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4266[15]), 
            .I3(n40594), .O(delay_counter_15__N_3989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_12 (.CI(n40594), .I0(delay_counter[10]), .I1(n4266[15]), 
            .CO(n40595));
    SB_LUT4 add_961_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4266[15]), 
            .I3(n40593), .O(delay_counter_15__N_3989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_11 (.CI(n40593), .I0(delay_counter[9]), .I1(n4266[15]), 
            .CO(n40594));
    SB_LUT4 add_961_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4266[15]), 
            .I3(n40592), .O(delay_counter_15__N_3989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_10 (.CI(n40592), .I0(delay_counter[8]), .I1(n4266[15]), 
            .CO(n40593));
    SB_LUT4 add_961_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4266[15]), 
            .I3(n40591), .O(delay_counter_15__N_3989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_9 (.CI(n40591), .I0(delay_counter[7]), .I1(n4266[15]), 
            .CO(n40592));
    SB_LUT4 add_961_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4266[15]), 
            .I3(n40590), .O(delay_counter_15__N_3989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_8 (.CI(n40590), .I0(delay_counter[6]), .I1(n4266[15]), 
            .CO(n40591));
    SB_LUT4 add_961_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4266[15]), 
            .I3(n40589), .O(delay_counter_15__N_3989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_7 (.CI(n40589), .I0(delay_counter[5]), .I1(n4266[15]), 
            .CO(n40590));
    SB_LUT4 add_961_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4266[15]), 
            .I3(n40588), .O(delay_counter_15__N_3989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_6 (.CI(n40588), .I0(delay_counter[4]), .I1(n4266[15]), 
            .CO(n40589));
    SB_LUT4 add_961_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4266[15]), 
            .I3(n40587), .O(delay_counter_15__N_3989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_5 (.CI(n40587), .I0(delay_counter[3]), .I1(n4266[15]), 
            .CO(n40588));
    SB_LUT4 add_961_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4266[15]), 
            .I3(n40586), .O(delay_counter_15__N_3989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_4 (.CI(n40586), .I0(delay_counter[2]), .I1(n4266[15]), 
            .CO(n40587));
    SB_LUT4 add_961_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4266[15]), 
            .I3(n40585), .O(delay_counter_15__N_3989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22834_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4190), 
            .I3(GND_net), .O(n36514));   // verilog/eeprom.v(51[5:9])
    defparam i22834_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n46391), 
            .I3(enable_slow_N_4190), .O(n45666));   // verilog/eeprom.v(51[5:9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    i2c_controller i2c (.\state_7__N_4087[0] (\state_7__N_4087[0] ), .enable_slow_N_4190(enable_slow_N_4190), 
            .GND_net(GND_net), .sda_enable(sda_enable), .n4(n4), .CLK_c(CLK_c), 
            .scl_enable_N_4177(scl_enable_N_4177), .scl_enable(scl_enable), 
            .n6686(n6686), .\state[1] (\state[1]_adj_18 ), .\state[2] (\state[2] ), 
            .\state[3] (\state[3] ), .n35782(n35782), .n8(n8), .VCC_net(VCC_net), 
            .\state[0] (\state[0]_adj_19 ), .n4_adj_15(n4_adj_20), .\saved_addr[0] (\saved_addr[0] ), 
            .n6496(n6496), .n51120(n51120), .n15(n15), .n10(n10), .n28421(n28421), 
            .n28416(n28416), .n10_adj_16(n10_adj_21), .\state_7__N_4103[3] (\state_7__N_4103[3] ), 
            .n7227(n7227), .n30174(n30174), .n30159(n30159), .data({data}), 
            .n30158(n30158), .n30157(n30157), .n30146(n30146), .scl(scl), 
            .sda_out(sda_out), .n30138(n30138), .n30137(n30137), .n30136(n30136), 
            .n30135(n30135), .n10_adj_17(n10_adj_22), .enable(enable)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state_7__N_4087[0] , enable_slow_N_4190, GND_net, 
            sda_enable, n4, CLK_c, scl_enable_N_4177, scl_enable, 
            n6686, \state[1] , \state[2] , \state[3] , n35782, n8, 
            VCC_net, \state[0] , n4_adj_15, \saved_addr[0] , n6496, 
            n51120, n15, n10, n28421, n28416, n10_adj_16, \state_7__N_4103[3] , 
            n7227, n30174, n30159, data, n30158, n30157, n30146, 
            scl, sda_out, n30138, n30137, n30136, n30135, n10_adj_17, 
            enable) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state_7__N_4087[0] ;
    input enable_slow_N_4190;
    input GND_net;
    output sda_enable;
    output n4;
    input CLK_c;
    input scl_enable_N_4177;
    output scl_enable;
    output n6686;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    output n35782;
    input n8;
    input VCC_net;
    output \state[0] ;
    output n4_adj_15;
    output \saved_addr[0] ;
    input n6496;
    output n51120;
    output n15;
    output n10;
    output n28421;
    output n28416;
    output n10_adj_16;
    input \state_7__N_4103[3] ;
    input n7227;
    input n30174;
    input n30159;
    output [7:0]data;
    input n30158;
    input n30157;
    input n30146;
    output scl;
    output sda_out;
    input n30138;
    input n30137;
    input n30136;
    input n30135;
    input n10_adj_17;
    input enable;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire enable_slow_N_4189;
    wire [7:0]n119;
    
    wire n29828;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n29967, n20868, n7130, n29971;
    wire [0:0]n6532;
    
    wire n29968, sda_out_adj_4715;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n30055, i2c_clk_N_4176;
    wire [5:0]n29;
    
    wire n29709, n5, n36484, n35997, n36482, n45344, n47238, n51106, 
        n51051, n7, n4_adj_4717, n33, n37, n34, n11, n11_adj_4718, 
        n29561, n9, n12, n6679, n46397, n40769, n40768, n40767, 
        n40766, n40765, n35779, n11_adj_4721, n40764, n11_adj_4722, 
        n40763, n41907, n41906, n41905, n41904, n41903, n51137;
    
    SB_LUT4 i36376_2_lut (.I0(\state_7__N_4087[0] ), .I1(enable_slow_N_4190), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4189));   // verilog/i2c_controller.v(62[6:32])
    defparam i36376_2_lut.LUT_INIT = 16'h7777;
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n29828), .D(n119[7]), 
            .R(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n29828), .D(n119[6]), 
            .R(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n29828), .D(n119[5]), 
            .R(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n29828), .D(n119[4]), 
            .R(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n29828), .D(n119[3]), 
            .R(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n29828), .D(n119[2]), 
            .S(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n29828), .D(n119[1]), 
            .S(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7130), 
            .D(n20868), .S(n29971));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4715), .C(i2c_clk), .E(n29968), 
            .D(n6532[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n29828), .D(n119[0]), 
            .S(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_339_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_339_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n30055));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n30055), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4176));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4176));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4177));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFSR counter2_2202_2203__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4087[0] ), .C(CLK_c), .E(n29709), 
            .D(enable_slow_N_4189));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6686), .D(n5), 
            .S(n36484));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6686), .D(n35997), 
            .S(n36482));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6686), .D(n45344), 
            .S(n47238));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i22106_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35782));
    defparam i22106_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_338_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_15));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_338_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i35560_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n51106));   // verilog/i2c_controller.v(198[28:35])
    defparam i35560_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i35534_4_lut (.I0(n51106), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n51051));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i35534_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1620_i1_4_lut (.I0(n51051), .I1(\state[0] ), .I2(n6496), 
            .I3(\state[2] ), .O(n6532[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1620_i1_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(\state[1] ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4717));
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n29971));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i36421_4_lut (.I0(n6496), .I1(n34), .I2(n4_adj_4717), .I3(n37), 
            .O(n7130));
    defparam i36421_4_lut.LUT_INIT = 16'haf8c;
    SB_LUT4 i36392_2_lut (.I0(\state[0] ), .I1(n6496), .I2(GND_net), .I3(GND_net), 
            .O(n20868));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i36392_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i35556_3_lut_4_lut (.I0(n11), .I1(n11_adj_4718), .I2(enable_slow_N_4190), 
            .I3(\state_7__N_4087[0] ), .O(n51120));
    defparam i35556_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i36408_3_lut_4_lut (.I0(n11), .I1(n11_adj_4718), .I2(n15), 
            .I3(n6686), .O(n36484));
    defparam i36408_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n29561));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i36406_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4718), 
            .I3(n6686), .O(n36482));   // verilog/i2c_controller.v(151[5:14])
    defparam i36406_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n28421));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1510 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n28416));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1510.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_16));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_16), 
            .O(n6679));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30831_2_lut (.I0(\state_7__N_4103[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n46397));
    defparam i30831_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n6679), .I1(n46397), .I2(n7227), .I3(n37), 
            .O(n29828));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n40769), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n40768), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n40768), .I0(counter[6]), .I1(VCC_net), 
            .CO(n40769));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n40767), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n40767), .I0(counter[5]), .I1(VCC_net), 
            .CO(n40768));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n40766), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n40766), .I0(counter[4]), .I1(VCC_net), 
            .CO(n40767));
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n30174));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n30159));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30158));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30157));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n30146));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n40765), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i22831_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n35779));
    defparam i22831_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i36404_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6686), .O(n47238));
    defparam i36404_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 equal_263_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_263_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4721));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i30755_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n46397), .O(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i30755_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i22079_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i22079_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2565_2_lut (.I0(sda_out_adj_4715), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_39_add_2_5 (.CI(n40765), .I0(counter[3]), .I1(VCC_net), 
            .CO(n40766));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n40764), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4722));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_CARRY sub_39_add_2_4 (.CI(n40764), .I0(counter[2]), .I1(VCC_net), 
            .CO(n40765));
    SB_LUT4 i1_4_lut_4_lut_adj_1511 (.I0(\state[0] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(\state[2] ), .O(n29968));
    defparam i1_4_lut_4_lut_adj_1511.LUT_INIT = 16'h0316;
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n40763), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n40763), .I0(counter[1]), .I1(VCC_net), 
            .CO(n40764));
    SB_LUT4 counter2_2202_2203_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n41907), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2202_2203_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n41906), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2202_2203_add_4_6 (.CI(n41906), .I0(GND_net), .I1(counter2[4]), 
            .CO(n41907));
    SB_LUT4 counter2_2202_2203_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n41905), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2202_2203_add_4_5 (.CI(n41905), .I0(GND_net), .I1(counter2[3]), 
            .CO(n41906));
    SB_LUT4 counter2_2202_2203_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n41904), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2202_2203_add_4_4 (.CI(n41904), .I0(GND_net), .I1(counter2[2]), 
            .CO(n41905));
    SB_LUT4 counter2_2202_2203_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n41903), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2202_2203_add_4_3 (.CI(n41903), .I0(GND_net), .I1(counter2[1]), 
            .CO(n41904));
    SB_LUT4 counter2_2202_2203_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2202_2203_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n30138));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n30137));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30136));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n30135));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2202_2203__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2202_2203__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2202_2203__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2202_2203__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2202_2203__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n30055));   // verilog/i2c_controller.v(69[20:35])
    SB_CARRY counter2_2202_2203_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n41903));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n40763));
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4718));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i35685_4_lut (.I0(n10_adj_17), .I1(n10), .I2(\state_7__N_4103[3] ), 
            .I3(enable), .O(n51137));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i35685_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n7), .I2(n51137), .I3(\state[0] ), 
            .O(n45344));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i36489_2_lut (.I0(\state_7__N_4103[3] ), .I1(n11_adj_4722), 
            .I2(GND_net), .I3(GND_net), .O(n35997));
    defparam i36489_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i36390_4_lut (.I0(n29561), .I1(n6679), .I2(n11), .I3(n35779), 
            .O(n6686));
    defparam i36390_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_1512 (.I0(n11_adj_4721), .I1(n11_adj_4722), .I2(\state_7__N_4103[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1512.LUT_INIT = 16'h5755;
    SB_LUT4 i1_2_lut_3_lut_adj_1513 (.I0(enable), .I1(\state_7__N_4087[0] ), 
            .I2(enable_slow_N_4190), .I3(GND_net), .O(n29709));
    defparam i1_2_lut_3_lut_adj_1513.LUT_INIT = 16'heaea;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\data[15] , \state[1] , \state[0] , n47264, GND_net, 
            n6, n15, n5, n5_adj_13, n35840, CLK_c, n30212, current, 
            n30211, n30210, n30209, n30208, n30207, n30206, n30205, 
            n30204, n30203, n30202, n30201, n30198, \data[0] , n10, 
            n9, n11, state_7__N_4293, n9_adj_14, clk_out, n30171, 
            CS_c, n30168, n30148, n30147, \data[12] , n30145, \data[11] , 
            n30144, \data[10] , n30143, \data[9] , n28429, n28432, 
            n30142, \data[8] , n30141, \data[7] , n28437, n30140, 
            \data[6] , n30139, \data[5] , n30134, \data[4] , n30133, 
            \data[3] , n30132, \data[2] , n30131, \data[1] , n28444, 
            VCC_net, CS_CLK_c, n28440) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \data[15] ;
    output \state[1] ;
    output \state[0] ;
    output n47264;
    input GND_net;
    output n6;
    output n15;
    output n5;
    output n5_adj_13;
    output n35840;
    input CLK_c;
    input n30212;
    output [12:0]current;
    input n30211;
    input n30210;
    input n30209;
    input n30208;
    input n30207;
    input n30206;
    input n30205;
    input n30204;
    input n30203;
    input n30202;
    input n30201;
    input n30198;
    output \data[0] ;
    output n10;
    output n9;
    output n11;
    output state_7__N_4293;
    input n9_adj_14;
    output clk_out;
    input n30171;
    output CS_c;
    input n30168;
    input n30148;
    input n30147;
    output \data[12] ;
    input n30145;
    output \data[11] ;
    input n30144;
    output \data[10] ;
    input n30143;
    output \data[9] ;
    output n28429;
    output n28432;
    input n30142;
    output \data[8] ;
    input n30141;
    output \data[7] ;
    output n28437;
    input n30140;
    output \data[6] ;
    input n30139;
    output \data[5] ;
    input n30134;
    output \data[4] ;
    input n30133;
    output \data[3] ;
    input n30132;
    output \data[2] ;
    input n30131;
    output \data[1] ;
    output n28444;
    input VCC_net;
    output CS_CLK_c;
    output n28440;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n35883;
    wire [7:0]n37;
    
    wire n29788, n30103, n11284, n29725, n29952, clk_slow_N_4206, 
        n51069, n25309;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n6_adj_4711, clk_slow_N_4207, n1;
    wire [13:0]n61;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4288;
    wire [4:0]n25;
    
    wire n51099, n25320, n51100, n25318, n51104, n25316, n6_adj_4712, 
        n6_adj_4713, n47467, n47406, n47375, n41856, n41855, n41854, 
        n41853, n41852, n41851, n41850, n41849, n41848, n41847, 
        n41846, n41845, n41844, n41843, n41842, n41841, n41840, 
        n41808, n41807, n41806, n41805, n41804, n41803, n41802;
    
    SB_LUT4 i2_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n47264));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_319_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(52[9:26])
    defparam equal_319_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i36426_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n35883));
    defparam i36426_2_lut.LUT_INIT = 16'h1111;
    SB_DFFNESR bit_counter_2191__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n29788), 
            .D(n37[7]), .R(n30103));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2191__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n29788), 
            .D(n37[6]), .R(n30103));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2191__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n29788), 
            .D(n37[5]), .R(n30103));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2191__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n29788), 
            .D(n37[4]), .R(n30103));   // verilog/tli4970.v(53[24:39])
    SB_LUT4 equal_313_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(52[9:26])
    defparam equal_313_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_312_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_13));   // verilog/tli4970.v(52[9:26])
    defparam equal_312_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n29725), .D(n11284), 
            .R(n29952));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i22164_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n35840));
    defparam i22164_2_lut.LUT_INIT = 16'h8888;
    SB_DFF clk_slow_62 (.Q(clk_slow), .C(CLK_c), .D(clk_slow_N_4206));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 i11661_3_lut (.I0(\state[0] ), .I1(n51069), .I2(\state[1] ), 
            .I3(GND_net), .O(n25309));   // verilog/tli4970.v(53[24:39])
    defparam i11661_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n29725), .D(n35883), 
            .S(n29952));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i1 (.Q(current[1]), .C(clk_slow), .D(n30212));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i2 (.Q(current[2]), .C(clk_slow), .D(n30211));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i3 (.Q(current[3]), .C(clk_slow), .D(n30210));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i4 (.Q(current[4]), .C(clk_slow), .D(n30209));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i5 (.Q(current[5]), .C(clk_slow), .D(n30208));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i2_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4711));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2297_4_lut (.I0(counter[0]), .I1(counter[4]), .I2(n6_adj_4711), 
            .I3(counter[3]), .O(clk_slow_N_4207));
    defparam i2297_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 clk_slow_I_0_71_2_lut (.I0(clk_slow), .I1(clk_slow_N_4207), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4206));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_71_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4759_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // verilog/tli4970.v(41[5] 65[12])
    defparam i4759_1_lut.LUT_INIT = 16'h5555;
    SB_DFFN current_i0_i6 (.Q(current[6]), .C(clk_slow), .D(n30207));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i7 (.Q(current[7]), .C(clk_slow), .D(n30206));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i8 (.Q(current[8]), .C(clk_slow), .D(n30205));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i9 (.Q(current[9]), .C(clk_slow), .D(n30204));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i10 (.Q(current[10]), .C(clk_slow), .D(n30203));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i11 (.Q(current[11]), .C(clk_slow), .D(n30202));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i12 (.Q(current[12]), .C(clk_slow), .D(n30201));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30198));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNE bit_counter_2191__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n29788), 
            .D(n25309));   // verilog/tli4970.v(53[24:39])
    SB_DFFNSR delay_counter_2193_2194__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n61[0]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFSR counter_2195_2196__i1 (.Q(counter[0]), .C(CLK_c), .D(n25[0]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i11672_3_lut (.I0(\state[0] ), .I1(n51099), .I2(\state[1] ), 
            .I3(GND_net), .O(n25320));   // verilog/tli4970.v(53[24:39])
    defparam i11672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11670_3_lut (.I0(\state[0] ), .I1(n51100), .I2(\state[1] ), 
            .I3(GND_net), .O(n25318));   // verilog/tli4970.v(53[24:39])
    defparam i11670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11668_3_lut (.I0(\state[0] ), .I1(n51104), .I2(\state[1] ), 
            .I3(GND_net), .O(n25316));   // verilog/tli4970.v(53[24:39])
    defparam i11668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_256_i10_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/tli4970.v(54[12:26])
    defparam equal_256_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_256_i9_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/tli4970.v(54[12:26])
    defparam equal_256_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4712));   // verilog/tli4970.v(54[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_4712), .O(n15));   // verilog/tli4970.v(54[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1501 (.I0(delay_counter[5]), .I1(delay_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4713));
    defparam i2_2_lut_adj_1501.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(delay_counter[0]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[2]), .O(n47467));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1502 (.I0(n47467), .I1(n6_adj_4713), .I2(delay_counter[7]), 
            .I3(delay_counter[4]), .O(n47406));
    defparam i3_4_lut_adj_1502.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_1503 (.I0(n47406), .I1(delay_counter[8]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n47375));
    defparam i3_4_lut_adj_1503.LUT_INIT = 16'h8000;
    SB_LUT4 i2302_4_lut (.I0(n47375), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(delay_counter_15__N_4288));
    defparam i2302_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 mux_2294_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n11284));
    defparam mux_2294_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 state_7__I_0_76_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4293));   // verilog/tli4970.v(51[7:17])
    defparam state_7__I_0_76_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16192_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29788));
    defparam i16192_2_lut.LUT_INIT = 16'h6666;
    SB_DFFN clk_out_66 (.Q(clk_out), .C(clk_slow), .D(n9_adj_14));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN slave_select_65 (.Q(CS_c), .C(clk_slow), .D(n30171));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i0 (.Q(current[0]), .C(clk_slow), .D(n30168));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n30148));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n30147));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n30145));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n30144));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n30143));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[3]), 
            .I3(bit_counter[2]), .O(n28429));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1504 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n28432));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1504.LUT_INIT = 16'hffbf;
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n30142));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n30141));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i16414_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n30103));   // verilog/tli4970.v(53[24:39])
    defparam i16414_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 equal_256_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(54[12:26])
    defparam equal_256_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n28437));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n30140));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNE bit_counter_2191__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n29788), 
            .D(n25316));   // verilog/tli4970.v(53[24:39])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n30139));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNE bit_counter_2191__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n29788), 
            .D(n25318));   // verilog/tli4970.v(53[24:39])
    SB_DFFNE bit_counter_2191__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n29788), 
            .D(n25320));   // verilog/tli4970.v(53[24:39])
    SB_DFFNSR delay_counter_2193_2194__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n61[1]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n61[2]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n61[3]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n61[4]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n61[5]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n61[6]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n61[7]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n61[8]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n61[9]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n61[10]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n61[11]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i13 (.Q(delay_counter[12]), .C(clk_slow), 
            .D(n61[12]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2193_2194__i14 (.Q(delay_counter[13]), .C(clk_slow), 
            .D(n61[13]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFSR counter_2195_2196__i2 (.Q(counter[1]), .C(CLK_c), .D(n25[1]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2195_2196__i3 (.Q(counter[2]), .C(CLK_c), .D(n25[2]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2195_2196__i4 (.Q(counter[3]), .C(CLK_c), .D(n25[3]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2195_2196__i5 (.Q(counter[4]), .C(CLK_c), .D(n25[4]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n30134));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n30133));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n30132));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n30131));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1505 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n28444));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_4_lut_adj_1505.LUT_INIT = 16'hfffb;
    SB_LUT4 counter_2195_2196_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n41856), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2195_2196_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2195_2196_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n41855), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2195_2196_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2195_2196_add_4_5 (.CI(n41855), .I0(GND_net), .I1(counter[3]), 
            .CO(n41856));
    SB_LUT4 counter_2195_2196_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n41854), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2195_2196_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2195_2196_add_4_4 (.CI(n41854), .I0(GND_net), .I1(counter[2]), 
            .CO(n41855));
    SB_LUT4 counter_2195_2196_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n41853), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2195_2196_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2195_2196_add_4_3 (.CI(n41853), .I0(GND_net), .I1(counter[1]), 
            .CO(n41854));
    SB_LUT4 counter_2195_2196_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2195_2196_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2195_2196_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n41853));
    SB_LUT4 delay_counter_2193_2194_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n41852), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2193_2194_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n41851), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_14 (.CI(n41851), .I0(GND_net), 
            .I1(delay_counter[12]), .CO(n41852));
    SB_LUT4 delay_counter_2193_2194_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n41850), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_13 (.CI(n41850), .I0(GND_net), 
            .I1(delay_counter[11]), .CO(n41851));
    SB_LUT4 delay_counter_2193_2194_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n41849), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_12 (.CI(n41849), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n41850));
    SB_LUT4 delay_counter_2193_2194_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n41848), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_11 (.CI(n41848), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n41849));
    SB_LUT4 delay_counter_2193_2194_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n41847), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_10 (.CI(n41847), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n41848));
    SB_LUT4 delay_counter_2193_2194_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n41846), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_9 (.CI(n41846), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n41847));
    SB_LUT4 delay_counter_2193_2194_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n41845), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_8 (.CI(n41845), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n41846));
    SB_LUT4 delay_counter_2193_2194_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n41844), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_7 (.CI(n41844), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n41845));
    SB_LUT4 delay_counter_2193_2194_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n41843), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_6 (.CI(n41843), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n41844));
    SB_LUT4 delay_counter_2193_2194_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n41842), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_5 (.CI(n41842), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n41843));
    SB_LUT4 delay_counter_2193_2194_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n41841), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_4 (.CI(n41841), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n41842));
    SB_LUT4 delay_counter_2193_2194_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n41840), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2193_2194_add_4_3 (.CI(n41840), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n41841));
    SB_LUT4 delay_counter_2193_2194_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2193_2194_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY delay_counter_2193_2194_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n41840));
    SB_LUT4 bit_counter_2191_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n41808), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2191_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n41807), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2191_add_4_8 (.CI(n41807), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n41808));
    SB_LUT4 bit_counter_2191_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n41806), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2191_add_4_7 (.CI(n41806), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n41807));
    SB_LUT4 bit_counter_2191_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n41805), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2191_add_4_6 (.CI(n41805), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n41806));
    SB_LUT4 bit_counter_2191_add_4_5_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n41804), .O(n51099)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2191_add_4_5 (.CI(n41804), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n41805));
    SB_LUT4 bit_counter_2191_add_4_4_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n41803), .O(n51100)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2191_add_4_4 (.CI(n41803), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n41804));
    SB_LUT4 bit_counter_2191_add_4_3_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n41802), .O(n51104)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2191_add_4_3 (.CI(n41802), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n41803));
    SB_LUT4 bit_counter_2191_add_4_2_lut (.I0(n1), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n51069)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2191_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n41802));
    SB_LUT4 i1_2_lut_4_lut_adj_1506 (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4288), .O(n29725));
    defparam i1_2_lut_4_lut_adj_1506.LUT_INIT = 16'hfff4;
    SB_LUT4 i16263_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4288), .O(n29952));
    defparam i16263_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_LUT4 i1_2_lut_4_lut_adj_1507 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n28440));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_4_lut_adj_1507.LUT_INIT = 16'hffbf;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (b_prev, GND_net, a_new, direction_N_3907, 
            ENCODER0_B_N_keep, n1668, ENCODER0_A_N_keep, n30218, n1632, 
            encoder0_position, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3907;
    input ENCODER0_B_N_keep;
    input n1668;
    input ENCODER0_A_N_keep;
    input n30218;
    output n1632;
    output [31:0]encoder0_position;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3910, debounce_cnt, a_prev, direction_N_3906;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_3913, n30217, n30213;
    wire [31:0]n133;
    
    wire n41902, n41901, n41900, n41899, n41898, n41897, n41896, 
        n41895, n41894, n41893, n41892, n41891, n41890, n41889, 
        n41888, n41887, n41886, n41885, n41884, n41883, n41882, 
        n41881, n41880, n41879, n41878, n41877, n41876, n41875, 
        n41874, n41873, n41872;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36411_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i36411_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1632), .C(n1668), .D(n30218));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n30217));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n30213));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2201__i0 (.Q(encoder0_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i1 (.Q(encoder0_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i2 (.Q(encoder0_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i3 (.Q(encoder0_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i4 (.Q(encoder0_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i5 (.Q(encoder0_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i6 (.Q(encoder0_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i7 (.Q(encoder0_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i8 (.Q(encoder0_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i9 (.Q(encoder0_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i10 (.Q(encoder0_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i11 (.Q(encoder0_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i12 (.Q(encoder0_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i13 (.Q(encoder0_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i14 (.Q(encoder0_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i15 (.Q(encoder0_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i16 (.Q(encoder0_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i17 (.Q(encoder0_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i18 (.Q(encoder0_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i19 (.Q(encoder0_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i20 (.Q(encoder0_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i21 (.Q(encoder0_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i22 (.Q(encoder0_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i23 (.Q(encoder0_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i24 (.Q(encoder0_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i25 (.Q(encoder0_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i26 (.Q(encoder0_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i27 (.Q(encoder0_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i28 (.Q(encoder0_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i29 (.Q(encoder0_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i30 (.Q(encoder0_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2201__i31 (.Q(encoder0_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_2201_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[31]), .I3(n41902), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2201_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[30]), .I3(n41901), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_32 (.CI(n41901), .I0(direction_N_3906), 
            .I1(encoder0_position[30]), .CO(n41902));
    SB_LUT4 position_2201_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[29]), .I3(n41900), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_31 (.CI(n41900), .I0(direction_N_3906), 
            .I1(encoder0_position[29]), .CO(n41901));
    SB_LUT4 position_2201_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[28]), .I3(n41899), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_30 (.CI(n41899), .I0(direction_N_3906), 
            .I1(encoder0_position[28]), .CO(n41900));
    SB_LUT4 position_2201_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[27]), .I3(n41898), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_29 (.CI(n41898), .I0(direction_N_3906), 
            .I1(encoder0_position[27]), .CO(n41899));
    SB_LUT4 position_2201_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[26]), .I3(n41897), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_28 (.CI(n41897), .I0(direction_N_3906), 
            .I1(encoder0_position[26]), .CO(n41898));
    SB_LUT4 position_2201_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[25]), .I3(n41896), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_27 (.CI(n41896), .I0(direction_N_3906), 
            .I1(encoder0_position[25]), .CO(n41897));
    SB_LUT4 position_2201_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[24]), .I3(n41895), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_26 (.CI(n41895), .I0(direction_N_3906), 
            .I1(encoder0_position[24]), .CO(n41896));
    SB_LUT4 position_2201_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[23]), .I3(n41894), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_25 (.CI(n41894), .I0(direction_N_3906), 
            .I1(encoder0_position[23]), .CO(n41895));
    SB_LUT4 position_2201_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[22]), .I3(n41893), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_24 (.CI(n41893), .I0(direction_N_3906), 
            .I1(encoder0_position[22]), .CO(n41894));
    SB_LUT4 position_2201_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[21]), .I3(n41892), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_23 (.CI(n41892), .I0(direction_N_3906), 
            .I1(encoder0_position[21]), .CO(n41893));
    SB_LUT4 position_2201_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[20]), .I3(n41891), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_22 (.CI(n41891), .I0(direction_N_3906), 
            .I1(encoder0_position[20]), .CO(n41892));
    SB_LUT4 position_2201_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[19]), .I3(n41890), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_21 (.CI(n41890), .I0(direction_N_3906), 
            .I1(encoder0_position[19]), .CO(n41891));
    SB_LUT4 position_2201_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[18]), .I3(n41889), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_20 (.CI(n41889), .I0(direction_N_3906), 
            .I1(encoder0_position[18]), .CO(n41890));
    SB_LUT4 position_2201_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[17]), .I3(n41888), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_19 (.CI(n41888), .I0(direction_N_3906), 
            .I1(encoder0_position[17]), .CO(n41889));
    SB_LUT4 position_2201_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[16]), .I3(n41887), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_18 (.CI(n41887), .I0(direction_N_3906), 
            .I1(encoder0_position[16]), .CO(n41888));
    SB_LUT4 position_2201_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[15]), .I3(n41886), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_17 (.CI(n41886), .I0(direction_N_3906), 
            .I1(encoder0_position[15]), .CO(n41887));
    SB_LUT4 position_2201_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[14]), .I3(n41885), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_16 (.CI(n41885), .I0(direction_N_3906), 
            .I1(encoder0_position[14]), .CO(n41886));
    SB_LUT4 position_2201_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[13]), .I3(n41884), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_15 (.CI(n41884), .I0(direction_N_3906), 
            .I1(encoder0_position[13]), .CO(n41885));
    SB_LUT4 position_2201_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[12]), .I3(n41883), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_14 (.CI(n41883), .I0(direction_N_3906), 
            .I1(encoder0_position[12]), .CO(n41884));
    SB_LUT4 position_2201_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[11]), .I3(n41882), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_13 (.CI(n41882), .I0(direction_N_3906), 
            .I1(encoder0_position[11]), .CO(n41883));
    SB_LUT4 position_2201_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[10]), .I3(n41881), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_12 (.CI(n41881), .I0(direction_N_3906), 
            .I1(encoder0_position[10]), .CO(n41882));
    SB_LUT4 position_2201_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[9]), .I3(n41880), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_11 (.CI(n41880), .I0(direction_N_3906), 
            .I1(encoder0_position[9]), .CO(n41881));
    SB_LUT4 position_2201_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[8]), .I3(n41879), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_10 (.CI(n41879), .I0(direction_N_3906), 
            .I1(encoder0_position[8]), .CO(n41880));
    SB_LUT4 position_2201_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[7]), .I3(n41878), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_9 (.CI(n41878), .I0(direction_N_3906), 
            .I1(encoder0_position[7]), .CO(n41879));
    SB_LUT4 position_2201_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[6]), .I3(n41877), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_8 (.CI(n41877), .I0(direction_N_3906), 
            .I1(encoder0_position[6]), .CO(n41878));
    SB_LUT4 position_2201_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[5]), .I3(n41876), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_7 (.CI(n41876), .I0(direction_N_3906), 
            .I1(encoder0_position[5]), .CO(n41877));
    SB_LUT4 position_2201_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[4]), .I3(n41875), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_6 (.CI(n41875), .I0(direction_N_3906), 
            .I1(encoder0_position[4]), .CO(n41876));
    SB_LUT4 position_2201_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[3]), .I3(n41874), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_5 (.CI(n41874), .I0(direction_N_3906), 
            .I1(encoder0_position[3]), .CO(n41875));
    SB_LUT4 position_2201_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[2]), .I3(n41873), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_4 (.CI(n41873), .I0(direction_N_3906), 
            .I1(encoder0_position[2]), .CO(n41874));
    SB_LUT4 position_2201_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[1]), .I3(n41872), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_3 (.CI(n41872), .I0(direction_N_3906), 
            .I1(encoder0_position[1]), .CO(n41873));
    SB_LUT4 position_2201_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2201_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2201_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n41872));
    SB_LUT4 i16528_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n30217));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16524_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n30213));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16524_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (b_prev, GND_net, a_new, direction_N_3907, 
            ENCODER1_B_N_keep, n1668, ENCODER1_A_N_keep, n30219, n1673, 
            encoder1_position, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3907;
    input ENCODER1_B_N_keep;
    input n1668;
    input ENCODER1_A_N_keep;
    input n30219;
    output n1673;
    output [31:0]encoder1_position;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3910, debounce_cnt, a_prev, direction_N_3906;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_3913, n30220, n30199;
    wire [31:0]n133;
    
    wire n41839, n41838, n41837, n41836, n41835, n41834, n41833, 
        n41832, n41831, n41830, n41829, n41828, n41827, n41826, 
        n41825, n41824, n41823, n41822, n41821, n41820, n41819, 
        n41818, n41817, n41816, n41815, n41814, n41813, n41812, 
        n41811, n41810, n41809;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36414_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i36414_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n30220));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1673), .C(n1668), .D(n30219));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n30199));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2192__i0 (.Q(encoder1_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i1 (.Q(encoder1_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i2 (.Q(encoder1_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i3 (.Q(encoder1_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i4 (.Q(encoder1_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i5 (.Q(encoder1_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i6 (.Q(encoder1_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i7 (.Q(encoder1_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i8 (.Q(encoder1_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i9 (.Q(encoder1_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i10 (.Q(encoder1_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i11 (.Q(encoder1_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i12 (.Q(encoder1_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i13 (.Q(encoder1_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i14 (.Q(encoder1_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i15 (.Q(encoder1_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i16 (.Q(encoder1_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i17 (.Q(encoder1_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i18 (.Q(encoder1_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i19 (.Q(encoder1_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i20 (.Q(encoder1_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i21 (.Q(encoder1_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i22 (.Q(encoder1_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i23 (.Q(encoder1_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i24 (.Q(encoder1_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i25 (.Q(encoder1_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i26 (.Q(encoder1_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i27 (.Q(encoder1_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i28 (.Q(encoder1_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i29 (.Q(encoder1_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i30 (.Q(encoder1_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2192__i31 (.Q(encoder1_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_2192_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[31]), .I3(n41839), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2192_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[30]), .I3(n41838), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_32 (.CI(n41838), .I0(direction_N_3906), 
            .I1(encoder1_position[30]), .CO(n41839));
    SB_LUT4 position_2192_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[29]), .I3(n41837), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_31 (.CI(n41837), .I0(direction_N_3906), 
            .I1(encoder1_position[29]), .CO(n41838));
    SB_LUT4 position_2192_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[28]), .I3(n41836), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_30 (.CI(n41836), .I0(direction_N_3906), 
            .I1(encoder1_position[28]), .CO(n41837));
    SB_LUT4 position_2192_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[27]), .I3(n41835), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_29 (.CI(n41835), .I0(direction_N_3906), 
            .I1(encoder1_position[27]), .CO(n41836));
    SB_LUT4 position_2192_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[26]), .I3(n41834), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_28 (.CI(n41834), .I0(direction_N_3906), 
            .I1(encoder1_position[26]), .CO(n41835));
    SB_LUT4 position_2192_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[25]), .I3(n41833), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_27 (.CI(n41833), .I0(direction_N_3906), 
            .I1(encoder1_position[25]), .CO(n41834));
    SB_LUT4 position_2192_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[24]), .I3(n41832), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_26 (.CI(n41832), .I0(direction_N_3906), 
            .I1(encoder1_position[24]), .CO(n41833));
    SB_LUT4 position_2192_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[23]), .I3(n41831), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_25 (.CI(n41831), .I0(direction_N_3906), 
            .I1(encoder1_position[23]), .CO(n41832));
    SB_LUT4 position_2192_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[22]), .I3(n41830), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_24 (.CI(n41830), .I0(direction_N_3906), 
            .I1(encoder1_position[22]), .CO(n41831));
    SB_LUT4 position_2192_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[21]), .I3(n41829), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_23 (.CI(n41829), .I0(direction_N_3906), 
            .I1(encoder1_position[21]), .CO(n41830));
    SB_LUT4 position_2192_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[20]), .I3(n41828), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_22 (.CI(n41828), .I0(direction_N_3906), 
            .I1(encoder1_position[20]), .CO(n41829));
    SB_LUT4 position_2192_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[19]), .I3(n41827), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_21 (.CI(n41827), .I0(direction_N_3906), 
            .I1(encoder1_position[19]), .CO(n41828));
    SB_LUT4 position_2192_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[18]), .I3(n41826), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_20 (.CI(n41826), .I0(direction_N_3906), 
            .I1(encoder1_position[18]), .CO(n41827));
    SB_LUT4 position_2192_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[17]), .I3(n41825), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_19 (.CI(n41825), .I0(direction_N_3906), 
            .I1(encoder1_position[17]), .CO(n41826));
    SB_LUT4 position_2192_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[16]), .I3(n41824), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_18 (.CI(n41824), .I0(direction_N_3906), 
            .I1(encoder1_position[16]), .CO(n41825));
    SB_LUT4 position_2192_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[15]), .I3(n41823), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_17 (.CI(n41823), .I0(direction_N_3906), 
            .I1(encoder1_position[15]), .CO(n41824));
    SB_LUT4 position_2192_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[14]), .I3(n41822), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_16 (.CI(n41822), .I0(direction_N_3906), 
            .I1(encoder1_position[14]), .CO(n41823));
    SB_LUT4 position_2192_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[13]), .I3(n41821), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_15 (.CI(n41821), .I0(direction_N_3906), 
            .I1(encoder1_position[13]), .CO(n41822));
    SB_LUT4 position_2192_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[12]), .I3(n41820), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_14 (.CI(n41820), .I0(direction_N_3906), 
            .I1(encoder1_position[12]), .CO(n41821));
    SB_LUT4 position_2192_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[11]), .I3(n41819), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_13 (.CI(n41819), .I0(direction_N_3906), 
            .I1(encoder1_position[11]), .CO(n41820));
    SB_LUT4 position_2192_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[10]), .I3(n41818), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_12 (.CI(n41818), .I0(direction_N_3906), 
            .I1(encoder1_position[10]), .CO(n41819));
    SB_LUT4 position_2192_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[9]), .I3(n41817), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_11 (.CI(n41817), .I0(direction_N_3906), 
            .I1(encoder1_position[9]), .CO(n41818));
    SB_LUT4 position_2192_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[8]), .I3(n41816), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_10 (.CI(n41816), .I0(direction_N_3906), 
            .I1(encoder1_position[8]), .CO(n41817));
    SB_LUT4 position_2192_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[7]), .I3(n41815), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_9 (.CI(n41815), .I0(direction_N_3906), 
            .I1(encoder1_position[7]), .CO(n41816));
    SB_LUT4 position_2192_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[6]), .I3(n41814), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_8 (.CI(n41814), .I0(direction_N_3906), 
            .I1(encoder1_position[6]), .CO(n41815));
    SB_LUT4 position_2192_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[5]), .I3(n41813), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_7 (.CI(n41813), .I0(direction_N_3906), 
            .I1(encoder1_position[5]), .CO(n41814));
    SB_LUT4 position_2192_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[4]), .I3(n41812), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_6 (.CI(n41812), .I0(direction_N_3906), 
            .I1(encoder1_position[4]), .CO(n41813));
    SB_LUT4 position_2192_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[3]), .I3(n41811), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_5 (.CI(n41811), .I0(direction_N_3906), 
            .I1(encoder1_position[3]), .CO(n41812));
    SB_LUT4 position_2192_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[2]), .I3(n41810), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_4 (.CI(n41810), .I0(direction_N_3906), 
            .I1(encoder1_position[2]), .CO(n41811));
    SB_LUT4 position_2192_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[1]), .I3(n41809), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_3 (.CI(n41809), .I0(direction_N_3906), 
            .I1(encoder1_position[1]), .CO(n41810));
    SB_LUT4 position_2192_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2192_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2192_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n41809));
    SB_LUT4 i16531_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n30220));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16531_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16510_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n30199));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16510_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n30269, PWMLimit, CLK_c, n30268, n30267, n30266, n30265, 
            n30264, GND_net, \data_in_frame[1] , \data_in_frame[2] , 
            \FRAME_MATCHER.state , \FRAME_MATCHER.state[2] , \FRAME_MATCHER.state[3] , 
            n30263, n30262, n30261, rx_data_ready, \data_out_frame[16] , 
            \data_out_frame[18] , \data_out_frame[6] , \data_out_frame[7] , 
            \data_out_frame[4] , \data_out_frame[5] , n30260, n30259, 
            \data_out_frame[8] , \data_out_frame[9] , \data_out_frame[10] , 
            \data_out_frame[11] , \data_out_frame[14] , \data_out_frame[15] , 
            \data_out_frame[12] , \data_out_frame[13] , n30258, \data_out_frame[20] , 
            \data_out_frame[22] , \data_in[1] , \data_in[0] , \data_in[3] , 
            \data_in[2] , n771, \data_in_frame[3] , n4452, n28383, 
            n63, n3807, setpoint, n30257, n63_adj_3, n3303, n122, 
            n42261, n5, n53135, n30256, n30255, n30254, n30253, 
            \data_in_frame[9] , \data_in_frame[11] , \data_in_frame[13] , 
            \data_in_frame[5] , \data_in_frame[10] , n52967, \data_out_frame[23] , 
            tx_transmit_N_3513, \data_in_frame[12] , \data_in_frame[8] , 
            \data_out_frame[17] , \data_out_frame[19] , \data_out_frame[21][4] , 
            \data_out_frame[20][1] , \data_out_frame[21][1] , \data_out_frame[21][2] , 
            ID, DE_c, LED_c, \data_in_frame[4] , \data_in_frame[6] , 
            \data_out_frame[25] , \data_out_frame[24] , n47698, \data_out_frame[21][0] , 
            \data_out_frame[27][1] , n29783, \data_out_frame[20][0] , 
            \data_out_frame[21][3] , n25438, n42259, rx_data, tx_active, 
            n2025, n54, n46, n46338, \state[2] , \state[3] , n10, 
            n44944, n30166, n30165, control_mode, n30163, neopxl_color, 
            n30162, \Ki[0] , n30161, \Kp[0] , n30160, n30742, IntegralLimit, 
            n30741, n30740, n30739, n30738, n30737, n30736, n30735, 
            n30734, n30733, n30732, n30731, \state[0] , \state[1] , 
            enable_slow_N_4190, n7227, n30730, n30729, n30728, n30727, 
            n30726, n30725, n30724, n30723, n30722, n30721, n30719, 
            n30718, n30717, n30716, n30715, n30714, n30713, n30712, 
            n30711, n30710, n30709, n30708, n30707, n30706, n30705, 
            n30704, n30703, n30702, n30701, n30700, n30699, n30698, 
            n30697, n30696, n30695, n30694, n30693, n30692, n30691, 
            n30690, n30689, n30688, n30687, \Kp[1] , n30686, \Kp[2] , 
            n30685, \Kp[3] , n30684, \Kp[4] , n30683, \Kp[5] , n30682, 
            \Kp[6] , n30681, \Kp[7] , n30680, \Kp[8] , n30679, \Kp[9] , 
            n30678, \Kp[10] , n30677, \Kp[11] , n30676, \Kp[12] , 
            n30675, \Kp[13] , n30674, \Kp[14] , n30673, \Kp[15] , 
            n30671, \Ki[1] , n30670, \Ki[2] , n30669, \Ki[3] , n30668, 
            \Ki[4] , n30667, \Ki[5] , n30666, \Ki[6] , n30665, \Ki[7] , 
            n30664, \Ki[8] , n30663, \Ki[9] , n30662, \Ki[10] , 
            n30661, \Ki[11] , n30660, \Ki[12] , n30659, \Ki[13] , 
            n30658, \Ki[14] , n30657, \Ki[15] , n30656, n30655, 
            n30654, n30653, n30652, n30651, n30650, n30649, n30648, 
            n30647, n30646, n30645, n30644, n30643, n30642, n30641, 
            n30640, n30639, n30638, n30637, n30636, n30635, n30634, 
            n30633, n30632, n30631, n30630, n30629, n30628, n30627, 
            n30626, n30625, n30624, n30623, n30622, n30621, n30620, 
            n30619, n30618, n30617, n30616, n30615, n30614, n30613, 
            n30612, n30611, n30610, n30609, n30608, n30607, n30606, 
            n30605, n30604, n30603, n30602, n30601, n30600, n30599, 
            n30598, n30597, n30596, n30595, n30594, n30593, n30592, 
            n30591, n30590, n30589, n30588, n30587, n30586, n30585, 
            n30584, n30583, n30582, n30581, n30580, n30579, n30578, 
            n30577, n30576, n30575, n30574, n30573, n30572, n30571, 
            n30570, n30569, n30568, n30567, n30566, n30565, n30564, 
            n30563, n30562, n30561, n30560, n30559, n30558, n30557, 
            n30556, n30555, n30554, n30553, n30552, n30551, n30550, 
            n30549, n30548, n30547, n30546, n30545, n30544, n30543, 
            n30542, n30541, n30540, n30539, n30538, n30537, n30536, 
            n30535, n30534, n30533, n30532, n30531, n30530, n30529, 
            n30528, n30527, n30526, n30525, n30523, n30522, n30521, 
            n30520, n30519, n30518, n30517, n30516, n30515, n30514, 
            n30513, n30512, n30511, n30510, n30509, n30508, n30507, 
            n30505, n30504, n30503, n30502, n30500, n30499, n30498, 
            n30497, n30496, n30495, n30494, n30493, n30492, n30491, 
            n30490, n30489, n30488, n30487, n30486, n30485, n30484, 
            n30483, n30482, n30481, n30480, n30479, n30478, n30477, 
            n30476, n30475, n30474, n30473, n30472, n30471, n30470, 
            n30469, n30468, n30467, n30466, n30465, n30464, n30463, 
            n30462, n30461, n30460, n30459, n30458, n30124, n30282, 
            n30281, n30280, n30279, n30278, n30277, n30276, n30275, 
            n30274, n30273, n30272, n29618, n30271, n30270, n15, 
            scl_enable_N_4177, n6496, n5_adj_4, n45649, \displacement[4] , 
            n25701, n47127, n46329, r_SM_Main, n20694, \r_Bit_Index[0] , 
            tx_o, n29684, n45512, \r_SM_Main_2__N_3613[1] , n53023, 
            n30173, n4, n30186, VCC_net, tx_enable, n29701, n4_adj_5, 
            n4_adj_6, \r_Bit_Index[0]_adj_7 , n28484, n35741, r_SM_Main_adj_12, 
            r_Rx_Data, \r_SM_Main_2__N_3542[2] , RX_N_10, n28489, n4_adj_11, 
            n30197, n45507, n30156, n30155, n30154, n30153, n30152, 
            n30151, n30150, n45602, n29660, n30189, n45162) /* synthesis syn_module_defined=1 */ ;
    input n30269;
    output [23:0]PWMLimit;
    input CLK_c;
    input n30268;
    input n30267;
    input n30266;
    input n30265;
    input n30264;
    input GND_net;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output [31:0]\FRAME_MATCHER.state ;
    output \FRAME_MATCHER.state[2] ;
    output \FRAME_MATCHER.state[3] ;
    input n30263;
    input n30262;
    input n30261;
    output rx_data_ready;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    input n30260;
    input n30259;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    input n30258;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[2] ;
    output n771;
    output [7:0]\data_in_frame[3] ;
    output n4452;
    output n28383;
    output n63;
    output n3807;
    output [23:0]setpoint;
    input n30257;
    output n63_adj_3;
    output n3303;
    output n122;
    output n42261;
    output n5;
    output n53135;
    input n30256;
    input n30255;
    input n30254;
    input n30253;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[10] ;
    input n52967;
    output [7:0]\data_out_frame[23] ;
    output tx_transmit_N_3513;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[19] ;
    output \data_out_frame[21][4] ;
    output \data_out_frame[20][1] ;
    output \data_out_frame[21][1] ;
    output \data_out_frame[21][2] ;
    input [7:0]ID;
    output DE_c;
    output LED_c;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    output n47698;
    output \data_out_frame[21][0] ;
    output \data_out_frame[27][1] ;
    output n29783;
    output \data_out_frame[20][0] ;
    output \data_out_frame[21][3] ;
    output n25438;
    output n42259;
    output [7:0]rx_data;
    output tx_active;
    output n2025;
    output n54;
    output n46;
    output n46338;
    input \state[2] ;
    input \state[3] ;
    output n10;
    input n44944;
    input n30166;
    input n30165;
    output [7:0]control_mode;
    input n30163;
    output [23:0]neopxl_color;
    input n30162;
    output \Ki[0] ;
    input n30161;
    output \Kp[0] ;
    input n30160;
    input n30742;
    output [23:0]IntegralLimit;
    input n30741;
    input n30740;
    input n30739;
    input n30738;
    input n30737;
    input n30736;
    input n30735;
    input n30734;
    input n30733;
    input n30732;
    input n30731;
    input \state[0] ;
    input \state[1] ;
    output enable_slow_N_4190;
    output n7227;
    input n30730;
    input n30729;
    input n30728;
    input n30727;
    input n30726;
    input n30725;
    input n30724;
    input n30723;
    input n30722;
    input n30721;
    input n30719;
    input n30718;
    input n30717;
    input n30716;
    input n30715;
    input n30714;
    input n30713;
    input n30712;
    input n30711;
    input n30710;
    input n30709;
    input n30708;
    input n30707;
    input n30706;
    input n30705;
    input n30704;
    input n30703;
    input n30702;
    input n30701;
    input n30700;
    input n30699;
    input n30698;
    input n30697;
    input n30696;
    input n30695;
    input n30694;
    input n30693;
    input n30692;
    input n30691;
    input n30690;
    input n30689;
    input n30688;
    input n30687;
    output \Kp[1] ;
    input n30686;
    output \Kp[2] ;
    input n30685;
    output \Kp[3] ;
    input n30684;
    output \Kp[4] ;
    input n30683;
    output \Kp[5] ;
    input n30682;
    output \Kp[6] ;
    input n30681;
    output \Kp[7] ;
    input n30680;
    output \Kp[8] ;
    input n30679;
    output \Kp[9] ;
    input n30678;
    output \Kp[10] ;
    input n30677;
    output \Kp[11] ;
    input n30676;
    output \Kp[12] ;
    input n30675;
    output \Kp[13] ;
    input n30674;
    output \Kp[14] ;
    input n30673;
    output \Kp[15] ;
    input n30671;
    output \Ki[1] ;
    input n30670;
    output \Ki[2] ;
    input n30669;
    output \Ki[3] ;
    input n30668;
    output \Ki[4] ;
    input n30667;
    output \Ki[5] ;
    input n30666;
    output \Ki[6] ;
    input n30665;
    output \Ki[7] ;
    input n30664;
    output \Ki[8] ;
    input n30663;
    output \Ki[9] ;
    input n30662;
    output \Ki[10] ;
    input n30661;
    output \Ki[11] ;
    input n30660;
    output \Ki[12] ;
    input n30659;
    output \Ki[13] ;
    input n30658;
    output \Ki[14] ;
    input n30657;
    output \Ki[15] ;
    input n30656;
    input n30655;
    input n30654;
    input n30653;
    input n30652;
    input n30651;
    input n30650;
    input n30649;
    input n30648;
    input n30647;
    input n30646;
    input n30645;
    input n30644;
    input n30643;
    input n30642;
    input n30641;
    input n30640;
    input n30639;
    input n30638;
    input n30637;
    input n30636;
    input n30635;
    input n30634;
    input n30633;
    input n30632;
    input n30631;
    input n30630;
    input n30629;
    input n30628;
    input n30627;
    input n30626;
    input n30625;
    input n30624;
    input n30623;
    input n30622;
    input n30621;
    input n30620;
    input n30619;
    input n30618;
    input n30617;
    input n30616;
    input n30615;
    input n30614;
    input n30613;
    input n30612;
    input n30611;
    input n30610;
    input n30609;
    input n30608;
    input n30607;
    input n30606;
    input n30605;
    input n30604;
    input n30603;
    input n30602;
    input n30601;
    input n30600;
    input n30599;
    input n30598;
    input n30597;
    input n30596;
    input n30595;
    input n30594;
    input n30593;
    input n30592;
    input n30591;
    input n30590;
    input n30589;
    input n30588;
    input n30587;
    input n30586;
    input n30585;
    input n30584;
    input n30583;
    input n30582;
    input n30581;
    input n30580;
    input n30579;
    input n30578;
    input n30577;
    input n30576;
    input n30575;
    input n30574;
    input n30573;
    input n30572;
    input n30571;
    input n30570;
    input n30569;
    input n30568;
    input n30567;
    input n30566;
    input n30565;
    input n30564;
    input n30563;
    input n30562;
    input n30561;
    input n30560;
    input n30559;
    input n30558;
    input n30557;
    input n30556;
    input n30555;
    input n30554;
    input n30553;
    input n30552;
    input n30551;
    input n30550;
    input n30549;
    input n30548;
    input n30547;
    input n30546;
    input n30545;
    input n30544;
    input n30543;
    input n30542;
    input n30541;
    input n30540;
    input n30539;
    input n30538;
    input n30537;
    input n30536;
    input n30535;
    input n30534;
    input n30533;
    input n30532;
    input n30531;
    input n30530;
    input n30529;
    input n30528;
    input n30527;
    input n30526;
    input n30525;
    input n30523;
    input n30522;
    input n30521;
    input n30520;
    input n30519;
    input n30518;
    input n30517;
    input n30516;
    input n30515;
    input n30514;
    input n30513;
    input n30512;
    input n30511;
    input n30510;
    input n30509;
    input n30508;
    input n30507;
    input n30505;
    input n30504;
    input n30503;
    input n30502;
    input n30500;
    input n30499;
    input n30498;
    input n30497;
    input n30496;
    input n30495;
    input n30494;
    input n30493;
    input n30492;
    input n30491;
    input n30490;
    input n30489;
    input n30488;
    input n30487;
    input n30486;
    input n30485;
    input n30484;
    input n30483;
    input n30482;
    input n30481;
    input n30480;
    input n30479;
    input n30478;
    input n30477;
    input n30476;
    input n30475;
    input n30474;
    input n30473;
    input n30472;
    input n30471;
    input n30470;
    input n30469;
    input n30468;
    input n30467;
    input n30466;
    input n30465;
    input n30464;
    input n30463;
    input n30462;
    input n30461;
    input n30460;
    input n30459;
    input n30458;
    input n30124;
    input n30282;
    input n30281;
    input n30280;
    input n30279;
    input n30278;
    input n30277;
    input n30276;
    input n30275;
    input n30274;
    input n30273;
    input n30272;
    output n29618;
    input n30271;
    input n30270;
    input n15;
    output scl_enable_N_4177;
    output n6496;
    output n5_adj_4;
    input n45649;
    input \displacement[4] ;
    output n25701;
    output n47127;
    input n46329;
    output [2:0]r_SM_Main;
    output n20694;
    output \r_Bit_Index[0] ;
    output tx_o;
    output n29684;
    output n45512;
    output \r_SM_Main_2__N_3613[1] ;
    input n53023;
    input n30173;
    output n4;
    input n30186;
    input VCC_net;
    output tx_enable;
    output n29701;
    output n4_adj_5;
    output n4_adj_6;
    output \r_Bit_Index[0]_adj_7 ;
    output n28484;
    output n35741;
    output [2:0]r_SM_Main_adj_12;
    output r_Rx_Data;
    output \r_SM_Main_2__N_3542[2] ;
    input RX_N_10;
    output n28489;
    output n4_adj_11;
    input n30197;
    output n45507;
    input n30156;
    input n30155;
    input n30154;
    input n30153;
    input n30152;
    input n30151;
    input n30150;
    input n45602;
    output n29660;
    input n30189;
    input n45162;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire Kp_23__N_969, n45804, n45767, n16, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n46249, n21, n17, n28750, n61, n24, n29147, n50003, 
        n20, n6;
    wire [31:0]\FRAME_MATCHER.state_31__N_2724 ;
    
    wire n43663, n46468, n43664, n47799, n63_c;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(112[11:16])
    
    wire n15_c, n67, n4_c, n48237;
    wire [7:0]n8825;
    
    wire n29645;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n39711, n36474, n3059, \FRAME_MATCHER.rx_data_ready_prev , 
        n161, n42875, n46187, n28663, n28910, n42894, n50179, 
        n50180, n50178, n52927, n51118, n50173, n50174, n50172, 
        n52939, n51122, n52903, n52765, n51822, n50283, n50284, 
        n50305, n50304, n50220, n50221, n50299, n50298, n50301, 
        n50302, n50224, n50223, n40527, n40526, n45947, n43975, 
        n43038, n46098, n50289, n50290, n50275, n50274, n50235, 
        n50236, n50263, n50262, n50244, n50245, n50227, n50226, 
        n50250, n50251, n50197, n50196, n50271, n50272, n50164, 
        n50163, n50167, n50168, n50166, n52945, n51117, n50159, 
        n50157;
    wire [0:0]n4882;
    wire [2:0]r_SM_Main_2__N_3616;
    
    wire n7099, n52951, n51116, n16_adj_4408, n17_adj_4409, n28397, 
        n28295, n16_adj_4410, n17_adj_4411, n63_adj_4412, n28472, 
        n28478, n18, n20_adj_4413, n15_adj_4414, n63_adj_4415, n6_adj_4416, 
        n28274, n42507, n62;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n6997, n8, n28400, n40525, n28386, n8_adj_4418, n36220, 
        n28426, n45, n38, n10_c, n6998, n6996, n29629, n44, 
        n42, n43, n41, n40, n39, n50, n6999, n45_adj_4419, n10_adj_4420, 
        n14, n14_adj_4421, n7000, n15_adj_4422, n20_adj_4423, n19, 
        n50065, n7001, n7002, n40524, n28276, n7003, n40523, n40522, 
        n45955, n45944, n29261, n45865, n28835, n46163, n46107;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n45750, n14_adj_4425, n46260, n46025, n15_adj_4426, n28776, 
        Kp_23__N_1803, n29105, n45853, n28861, n4_adj_4427, n46209, 
        n46101, n16_adj_4428, n46919, n8_adj_4429, n43827, n17_adj_4430, 
        n43836, n46269, n43800;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n45764, n48165, n46008, n46011;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n46030, n29210, n46014, n46160, n8_adj_4431;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n7004, n29195, n46042, n46219, n47604, n42975, n72, n45913, 
        n46166, n46036, n45996, n78, n50188, n52921, n51136, n40521;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire Kp_23__N_1321, n76, n50143, n46282, n46266, n77, n20_adj_4432, 
        n45724, n75, n46064, n74, n50189, n46216, n45987, n47973, 
        n73, n90, n50187, n43017, n10_adj_4433, n46285, n83, n7005, 
        n42954, n82, n42873, n80, n29188, n43915, n81, n45961, 
        n79, n52747, n50144, n50131, n92, n6_adj_4434, n91, n7, 
        n52843, n50130;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n47090, n47108, n47097, n47333, n29, n5_adj_4435, n7006, 
        n10_adj_4436, n45718, n45706, n46196, n6_adj_4437, n52915, 
        n51134, n50146, n20_adj_4438, n46089, n29255, n43889, n27975, 
        n43795, n12, n45885, n6_adj_4439, n50195, n28674, n50193, 
        n28809, n52777, n50147, n50137, n7_adj_4440, n52837, n50136, 
        Kp_23__N_1195, n6_adj_4441, n46240, n10_adj_4442, n46092, 
        n6_adj_4443, n28892, n46020, n28827, n42988, n46203, n12_adj_4444, 
        n42892, n45999, n43606, n52909, n51132, n50149, n10_adj_4445, 
        n14_adj_4446, n20_adj_4447, n50204, n50202, n52783, n50150, 
        n50140, n7_adj_4448, n52825, n50139, n46279, n46193, n46273, 
        n10_adj_4449, n45875, n14_adj_4450, n46225, n45973, n46184, 
        n45715, n10_adj_4451, n45910, n43430, n46049, n42921, n12_adj_4452, 
        n7007, n45930, n43899, n6_adj_4453, Kp_23__N_1285, n29226, 
        n29505, n7008, n7009, n29268, n46054, n6_adj_4454, n7010, 
        n2_adj_4455, n40520, n46257, n14_adj_4456, n10_adj_4457, n45936, 
        n28565, n6_adj_4458, n43811, n28815, n34, n50027, n24_adj_4459, 
        n54_c, n2_adj_4460, n40519, n42655, n18_adj_4461, n46136, 
        n19_adj_4462, n45991, n12_adj_4463, n46228, n45827, n14_adj_4464, 
        n10_adj_4465, n45817, n2_adj_4466, n40518, n14_adj_4467, n13, 
        n50238, n50239, n50242;
    wire [7:0]\data_out_frame[20]_c ;   // verilog/coms.v(97[12:26])
    
    wire n50241, n50277, n50278, n50281, n50280, n50256, n50257, 
        n50269, n50268, n7011, n9, n8_adj_4468, n2_adj_4469, n40517, 
        n7_adj_4470, n9_adj_4471, n49, n35937, n46478, n36742, n29930, 
        n28791, n45781, n10_adj_4472, n45795, n45958, n12_adj_4473, 
        n46130, n14_adj_4474, n10_adj_4475, n11, Kp_23__N_1020, n28870, 
        n13_adj_4476, n7012, Kp_23__N_1093, n7_adj_4477, n28761, n8_adj_4478, 
        n6_adj_4479, n29223, n45916, n28578, n48160, n46002, n10_adj_4480, 
        n47661, n43816, n47627, n2134, n43832, n6_adj_4481, n47566, 
        n46061, n43803, n46181, n10_adj_4482, n47422, n2_adj_4483, 
        n40516, n7013, n42864, n47800, n45801, n7014, n29481, 
        n46046, n10_adj_4484, n47041, n48100, n45841, n12_adj_4485, 
        n46148, n29389, n45733, n2_adj_4486, n40515, n43906, n12_adj_4487, 
        n46222, n48133, n47769, n46033, n28003, n12_adj_4488, n46095, 
        n46928, n43860, n10_adj_4489, n7019, n7018, n7017, n7016, 
        n7015, n45721, n45676, n15_adj_4490, n6_adj_4491, n14_adj_4492, 
        n47644, n45952, n45821, n28981, Kp_23__N_988, n28977, n45580, 
        n44886, n45830, n6_adj_4493, n45696, n42909, n14_adj_4494, 
        n28990, n10_adj_4495, n45777, n6_adj_4496, n29502, n29529, 
        n10_adj_4497, n27216, n46139, n10_adj_4498, n29171, n45862, 
        n46124, n45689, n27979, n29134, n45693, n45859, n29137, 
        n28702, n46142, n45967, n10_adj_4499, n45919, n28997, n45729, 
        n46071, n16_adj_4500, n45678, n46104, n17_adj_4501, n4_adj_4502, 
        n45787, n45983, n45673, n62_adj_4503, n12_adj_4504, n45907, 
        n47414, n28741, n43910, n45784, n28, n43007, n26, n27, 
        n43846, n43805, n1563, n45752, n25, n46246, n28941, n29044, 
        n10_adj_4505, n29164, n2_adj_4506, n40514, n46263, n48327, 
        n26683, n40_adj_4507, n48347, n38_adj_4508, n28595, n39_adj_4509, 
        n37, n45872, n42_adj_4510, n46_c, n41_adj_4511, n46077, 
        n6_adj_4512, n6_adj_4513, n46119, n46127, n12_adj_4514, n46213, 
        n46058, n60, n45893, n48336, n43_adj_4515, n45674, n70, 
        n47706, n68, n42936, n45939, n69, n45758, n25_adj_4516, 
        n42930, n67_adj_4517, n11_adj_4518, n48, n46206, n64, n42898, 
        n66, n6_adj_4519, n47199, n30, n45881, n45970, n45755, 
        n65, n28_adj_4520, n76_adj_4521, n29_adj_4522, n71, n27_adj_4523, 
        n43858, n43834, n45635, n32424, n45761, n46112, n29034, 
        n15_adj_4524, n14_adj_4525, n27987, n7_adj_4526, n8_adj_4527, 
        n48169, n10_adj_4528, n25_adj_4529, n11_adj_4530, n45882, 
        n46157, n46253, n10_adj_4531, n45850, n46005, n12_adj_4532, 
        n43854, n8_adj_4533, n51996, n45933, n10_adj_4534, n47476, 
        n46908, n6_adj_4535, n46175, n6_adj_4536, n29296, n46154, 
        n46145, n10_adj_4537, n8_adj_4538, n45856, n12_adj_4539, n26646, 
        n47315, n45770, n12_adj_4540, n46115, n28719, n46039, n10_adj_4541, 
        n28127, n47174, n29020, n10_adj_4542, n48173, n4_adj_4543, 
        n29458, n45896, n15_adj_4544, n45712, n14_adj_4545, n29380, 
        n8_adj_4546, n45964, n46231, n48076, n2_adj_4547, n40513, 
        n2_adj_4548, n40512, n20_adj_4549, n19_adj_4550, n21_adj_4551, 
        n45486, n160, n45614, n2_adj_4552, n40511, n2_adj_4553, 
        n40510, n6_adj_4554, n7_adj_4555, n45670, n7_adj_4556, n44942, 
        n4_adj_4557, n51760, n51114, n52960, n52819, n7_adj_4558;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n52954, n52957, n45102, n44946, n45040, n42278, n45098, 
        n44910, n45094, n44948, n7_adj_4559, n35660, n7_adj_4560, 
        n8_adj_4561, n45090, n44950, n35658, n36461, n45086, n44952, 
        n7_adj_4562, n8_adj_4563, n45082, n44954, n7_adj_4564, n8_adj_4565, 
        n7_adj_4566, n8_adj_4567, n45078, n42276, n35656, n8_adj_4568, 
        n45012, n44884, n45074, n44956, n45010, n44902, n35650, 
        n8_adj_4569, n6_adj_4570, n51044, n36547, n58, n8_adj_4571, 
        n45491, n45070, n44958, n52948, n45066, n44960, n45062, 
        n44962, n45058, n44964, n45054, n44966, n45006, n44968, 
        n45050, n44892, n44896, n10_adj_4572, n44890, n52972, n45745, 
        n2_adj_4573, n40509, n35635, n45616, n48289, n52942, n1519, 
        n28528, n1516, n1168, n45703, n29293, n45837, n46086, 
        n46237, n52936, n52924, n52918, n52912, n52906, n52900, 
        n43979, n16_adj_4574, n17_adj_4575, n45685, n3_adj_4576, n3_adj_4577, 
        n3_adj_4578, n3_adj_4579, n3_adj_4580, n3_adj_4581, n3_adj_4582, 
        n3_adj_4583, n3_adj_4584, n3_adj_4585, n3_adj_4586, n3_adj_4587, 
        n2_adj_4588, n3_adj_4589, n2_adj_4590, n3_adj_4591, n2_adj_4592, 
        n3_adj_4593, n2_adj_4594, n3_adj_4595, n2_adj_4596, n3_adj_4597, 
        n2_adj_4598, n3_adj_4599, n2_adj_4600, n3_adj_4601, n2_adj_4602, 
        n3_adj_4603, n2_adj_4604, n3_adj_4605, n18_adj_4606, n2_adj_4607, 
        n3_adj_4608, n2_adj_4609, n3_adj_4610, n2_adj_4611, n3_adj_4612, 
        n2_adj_4613, n3_adj_4614, n2_adj_4615, n3_adj_4616, n2_adj_4617, 
        n3_adj_4618, n2_adj_4619, n3_adj_4620, n2_adj_4621, n3_adj_4622, 
        n2_adj_4623, n3_adj_4624, n2_adj_4625, n3_adj_4626, Kp_23__N_993, 
        n16_adj_4627, n45737, n20_adj_4628, n46178, n28113, n45869, 
        n40508, n45901, n6_adj_4629, n6_adj_4630, n12_adj_4631, n45824, 
        n6_adj_4632, n45846, n46151, n10_adj_4633, n1668, n45976, 
        n28510, n46169, n1247, n12_adj_4634, n46074, n28519, n46017, 
        n12_adj_4635, n6_adj_4636, n40507, n40506, n43121, n6_adj_4637, 
        n46172, n10_adj_4638, n45709, n6_adj_4639, n1537, n46234, 
        n1191, n45925, n28500, n40505, n52876, n45790, n18_adj_4640, 
        n40504, n20_adj_4641, n16_adj_4642, n47801, n18_adj_4643, 
        n30_adj_4644, n28_adj_4645, n40503, n45888, n29_adj_4646, 
        n46082, n27_adj_4647, n43887, n14_adj_4648, n13_adj_4649, 
        n9_adj_4650, n40502, n40501, n52879, n12_adj_4651, n45743, 
        n43025, n45699, n28542, n40500, n4_adj_4652, n10_adj_4653, 
        n52753, n52870, n52807, n7_adj_4654, n52759, n52864, n52861, 
        n7_adj_4655, n52858, n52852, n14_adj_4656, n52846, n14_adj_4657, 
        n52840, n52834, n14_adj_4658, n45814, n29091, n43940, n8_adj_4659, 
        n48270, n46276, n47669;
    wire [31:0]n1;
    
    wire n47182, n40499, n43862, n45642, n10_adj_4660, n3_adj_4661, 
        n18_adj_4662, n45651, n46495, n11_adj_4663, n6_adj_4664, n16_adj_4665, 
        n20_adj_4666, n40498, n52822, n40497, n40496, n46133, n8_adj_4667, 
        n45626, n30443, n40495, n52816, n52804, n52798, n7_adj_4668, 
        n52792, n52795, n40494, n30444, n40493, n30445, n30446, 
        n30447, n30448, n30449, n30450, n8_adj_4670, n30435, n30436, 
        n52741, n52786, n30437, n30438, n30439, n30440, n5_adj_4672, 
        n30441, n40492, n6_adj_4673;
    wire [31:0]\FRAME_MATCHER.state_31__N_2692 ;
    
    wire n30442, n8_adj_4674, n30427, n30428, n94, n94_adj_4675, 
        n28494, n30429, n7_adj_4676, n7_adj_4677, n25525, n30430, 
        n30431, n40491, n30432, n28389, n30433, n30434, n30164, 
        n40490, n18_adj_4679, n24_adj_4680, n22, n26_adj_4681, n8_adj_4682, 
        n45904, n10_adj_4683, n14_adj_4684, n43222, n53051, n12_adj_4685, 
        n43797;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n10_adj_4686, n43876, n47755, n6_adj_4687;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n6_adj_4688, n7_adj_4689, n47169, n50156, n50154, n7_adj_4690, 
        n117, n50155, n6_adj_4691, n46949, n8_adj_4692, n30524, 
        n30457, n30456, n30455, n30454, n30453, n30452, n30451, 
        n30426, n30425, n30424, n30423, n30422, n30421, n30420, 
        n30419, n30418, n30417, n30416, n30415, n30414, n30413, 
        n30412, n30411, n30410, n52780, n52774, n30409, n30408, 
        n30407, n30406, n30405, n30404, n30403, n30402, n30401, 
        n30400, n30399, n30398, n30397, n30396, n30395, n30394, 
        n30393, n30392, n30391, n30390, n30389, n30388, n30387, 
        n30386, n30385, n30384, n30383, n30382, n30381, n30380, 
        n30379, n30378, n30377, n30376, n30375, n30374, n30373, 
        n30372, n30371, n30370, n30369, n30368, n30367, n30366, 
        n30365, n30364, n30363, n30362, n30361, n30360, n30359, 
        n30358, n30357, n30356, n30355, n30354, n30353, n30352, 
        n30351, n30350, n30349, n30348, n30347, n30346, n30345, 
        n30344, n30343, n30342, n30341, n30340, n30339, n30338, 
        n30337, n30336, n30335, n30334, n30333, n30332, n30331, 
        n30330, n30329, n30328, n30327, n30326, n30325, n30324, 
        n30323, n30322, n30321, n30320, n30319, n30318, n30317, 
        n30316, n30315, n30314, n30313, n30312, n30311, n30310, 
        n30309, n30308, n30307, n30306, n30305, n30304, n30303, 
        n30302, n30301, n30300, n30299, n30298, n30297, n30296, 
        n30295, n30294, n30293, n30292, n30291, n30290, n30289, 
        n30288, n30287, n30286, n30285, n30284, n30283, n8_adj_4693, 
        n53041, n6_adj_4694, n47172, n8_adj_4695, n50031, n47094, 
        n36526, n50025, n46996, n8_adj_4697, n26_adj_4699, n32, 
        n47851, n45654, n52762, n52756, n52750, n52744, n7_adj_4700, 
        n52738;
    
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n30269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n30268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n30267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n30266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n30265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n30264));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_969), .I2(GND_net), 
            .I3(GND_net), .O(n45804));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(n45767), .I3(n45804), .O(n16));
    defparam i3_4_lut.LUT_INIT = 16'h1248;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut (.I0(n46249), .I1(n16), .I2(\data_in_frame[2] [0]), 
            .I3(n45804), .O(n21));
    defparam i8_4_lut.LUT_INIT = 16'h4004;
    SB_LUT4 i11_4_lut (.I0(n21), .I1(n17), .I2(n28750), .I3(n61), .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i34427_4_lut (.I0(\data_in_frame[0] [6]), .I1(n29147), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[0] [5]), .O(n50003));
    defparam i34427_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i1_4_lut (.I0(n50003), .I1(\data_in_frame[1] [6]), .I2(n24), 
            .I3(n20), .O(n6));
    defparam i1_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(n6), .O(\FRAME_MATCHER.state_31__N_2724 [3]));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i36384_4_lut (.I0(n43663), .I1(n46468), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n43664), .O(n47799));
    defparam i36384_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_867 (.I0(n63_c), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .O(n15_c));
    defparam i1_4_lut_adj_867.LUT_INIT = 16'ha0ac;
    SB_LUT4 i37079_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n15_c), .I2(n67), 
            .I3(n4_c), .O(n48237));
    defparam i37079_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 i2_3_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n46468));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n30263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n30262));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n29645), .D(n8825[1]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n29645), .D(n8825[2]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n29645), .D(n8825[3]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n29645), .D(n8825[4]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n29645), .D(n8825[5]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n29645), .D(n8825[6]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n29645), .D(n8825[7]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i22796_1_lut (.I0(n36474), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n3059));
    defparam i22796_1_lut.LUT_INIT = 16'h5555;
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n30261));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[16] [2]), .I1(n42875), .I2(\data_out_frame[16] [1]), 
            .I3(n46187), .O(n28663));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_868 (.I0(\data_out_frame[16] [2]), .I1(n42875), 
            .I2(\data_out_frame[18] [4]), .I3(n28910), .O(n42894));
    defparam i2_3_lut_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i34545_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50179));
    defparam i34545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34546_4_lut (.I0(n50179), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50180));
    defparam i34546_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i34544_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50178));
    defparam i34544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35679_2_lut (.I0(n52927), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51118));
    defparam i35679_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34539_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50173));
    defparam i34539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34540_4_lut (.I0(n50173), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50174));
    defparam i34540_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i34538_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50172));
    defparam i34538_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n30260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n30259));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i35571_2_lut (.I0(n52939), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51122));
    defparam i35571_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i36187_3_lut (.I0(n52903), .I1(n52765), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n51822));
    defparam i36187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34649_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50283));
    defparam i34649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34650_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50284));
    defparam i34650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34671_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50305));
    defparam i34671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34670_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50304));
    defparam i34670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34586_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50220));
    defparam i34586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34587_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50221));
    defparam i34587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34665_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50299));
    defparam i34665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34664_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50298));
    defparam i34664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34667_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50301));
    defparam i34667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34668_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50302));
    defparam i34668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34590_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50224));
    defparam i34590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34589_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50223));
    defparam i34589_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n30258));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n40527), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n40526), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_8 (.CI(n40526), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n40527));
    SB_LUT4 i1_2_lut_4_lut (.I0(n45947), .I1(\data_out_frame[20] [3]), .I2(n43975), 
            .I3(\data_out_frame[20] [2]), .O(n43038));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_869 (.I0(n45947), .I1(\data_out_frame[20] [3]), 
            .I2(n43975), .I3(\data_out_frame[22] [5]), .O(n46098));
    defparam i1_2_lut_4_lut_adj_869.LUT_INIT = 16'h9669;
    SB_LUT4 i34655_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50289));
    defparam i34655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34656_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50290));
    defparam i34656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34641_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50275));
    defparam i34641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34640_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50274));
    defparam i34640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34601_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50235));
    defparam i34601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34602_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50236));
    defparam i34602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34629_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50263));
    defparam i34629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34628_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50262));
    defparam i34628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34610_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50244));
    defparam i34610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34611_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50245));
    defparam i34611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34593_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50227));
    defparam i34593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34592_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50226));
    defparam i34592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34616_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50250));
    defparam i34616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34617_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50251));
    defparam i34617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34563_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50197));
    defparam i34563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34562_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50196));
    defparam i34562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34637_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50271));
    defparam i34637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34638_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50272));
    defparam i34638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34530_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50164));
    defparam i34530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34529_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50163));
    defparam i34529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34533_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50167));
    defparam i34533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34534_4_lut (.I0(n50167), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n50168));
    defparam i34534_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i34532_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50166));
    defparam i34532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35662_2_lut (.I0(n52945), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51117));
    defparam i35662_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34525_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n50159));
    defparam i34525_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34523_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50157));
    defparam i34523_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3616[0]), .C(CLK_c), .D(n4882[0]), 
            .R(n7099));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i35627_2_lut (.I0(n52951), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51116));
    defparam i35627_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n16_adj_4408));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [2]), .O(n17_adj_4409));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(n17_adj_4409), .I1(\data_in[1] [6]), .I2(n16_adj_4408), 
            .I3(\data_in[3] [7]), .O(n28397));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_870 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n28295), .O(n16_adj_4410));
    defparam i6_4_lut_adj_870.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_871 (.I0(n28397), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4411));
    defparam i7_4_lut_adj_871.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_872 (.I0(n17_adj_4411), .I1(\data_in[3] [5]), .I2(n16_adj_4410), 
            .I3(\data_in[3] [3]), .O(n63_adj_4412));
    defparam i9_4_lut_adj_872.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_873 (.I0(\data_in[2] [4]), .I1(n28472), .I2(\data_in[1] [5]), 
            .I3(n28478), .O(n18));
    defparam i7_4_lut_adj_873.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_874 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n28397), .O(n20_adj_4413));
    defparam i9_4_lut_adj_874.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4414));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4414), .I1(n20_adj_4413), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_4415));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4416));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_875 (.I0(\FRAME_MATCHER.i [0]), .I1(n6_adj_4416), 
            .I2(n28274), .I3(\FRAME_MATCHER.i [1]), .O(n42507));
    defparam i3_4_lut_adj_875.LUT_INIT = 16'hfefc;
    SB_LUT4 i22244_2_lut (.I0(n42507), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i22244_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_2021_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n6997));
    defparam mux_2021_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22250_4_lut (.I0(n8), .I1(\FRAME_MATCHER.i [31]), .I2(n28400), 
            .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i22250_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n40525), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_876 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n28386));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_876.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_3_lut (.I0(n36474), .I1(n28383), .I2(n63), .I3(GND_net), 
            .O(n8_adj_4418));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut_adj_877 (.I0(n36220), .I1(n8_adj_4418), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n28426), .O(n3807));
    defparam i4_4_lut_adj_877.LUT_INIT = 16'h8808;
    SB_LUT4 i1_2_lut_adj_878 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n45), 
            .I2(GND_net), .I3(GND_net), .O(n38));
    defparam i1_2_lut_adj_878.LUT_INIT = 16'heeee;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_7 (.CI(n40525), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n40526));
    SB_LUT4 i4_4_lut_adj_879 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_c));
    defparam i4_4_lut_adj_879.LUT_INIT = 16'hfdff;
    SB_LUT4 mux_2021_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n6998));
    defparam mux_2021_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut (.I0(\data_in[3] [4]), .I1(n10_c), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n28478));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n29629), .D(n6996));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_2021_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n6999));
    defparam mux_2021_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_4419));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45_adj_4419), .I1(n50), .I2(n39), .I3(n40), 
            .O(n28400));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_880 (.I0(\FRAME_MATCHER.i [4]), .I1(n28400), .I2(GND_net), 
            .I3(GND_net), .O(n28274));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_880.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_881 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4420));
    defparam i2_2_lut_adj_881.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_882 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14));
    defparam i6_4_lut_adj_882.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_883 (.I0(\data_in[3] [6]), .I1(n14), .I2(n10_adj_4420), 
            .I3(\data_in[2] [1]), .O(n28472));
    defparam i7_4_lut_adj_883.LUT_INIT = 16'hfffd;
    SB_LUT4 i5_3_lut_adj_884 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4421));
    defparam i5_3_lut_adj_884.LUT_INIT = 16'hdfdf;
    SB_LUT4 mux_2021_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n7000));
    defparam mux_2021_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_885 (.I0(\data_in[0] [6]), .I1(n28478), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4422));
    defparam i6_4_lut_adj_885.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_886 (.I0(n15_adj_4422), .I1(\data_in[3] [0]), .I2(n14_adj_4421), 
            .I3(\data_in[2] [2]), .O(n28295));
    defparam i8_4_lut_adj_886.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_887 (.I0(n28295), .I1(n28472), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [5]), .O(n20_adj_4423));
    defparam i8_4_lut_adj_887.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_888 (.I0(\data_in[2] [5]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[2] [6]), .O(n19));
    defparam i7_4_lut_adj_888.LUT_INIT = 16'hfffd;
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n30257));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34488_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[1] [2]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [1]), .O(n50065));
    defparam i34488_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mux_2021_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n7001));
    defparam mux_2021_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2021_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n7002));
    defparam mux_2021_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_3_lut (.I0(n50065), .I1(n19), .I2(n20_adj_4423), .I3(GND_net), 
            .O(n63_adj_3));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n40524), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22249_2_lut (.I0(n28276), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i22249_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i22339_3_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_4415), 
            .I2(n63_adj_4412), .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i22339_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_685_Select_2_i5_4_lut (.I0(n122), .I1(n42261), .I2(n3303), 
            .I3(n63_adj_3), .O(n5));
    defparam select_685_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i22335_rep_158_2_lut (.I0(n122), .I1(n63_adj_3), .I2(GND_net), 
            .I3(GND_net), .O(n53135));   // verilog/coms.v(142[4] 144[7])
    defparam i22335_rep_158_2_lut.LUT_INIT = 16'h8888;
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n30256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n30255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n30254));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_2021_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n7003));
    defparam mux_2021_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n30253));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_6 (.CI(n40524), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n40525));
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n40523), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_5 (.CI(n40523), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n40524));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n40522), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_4 (.CI(n40522), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n40523));
    SB_LUT4 i3_4_lut_adj_889 (.I0(n45955), .I1(\data_in_frame[9] [3]), .I2(\data_in_frame[11] [4]), 
            .I3(n45944), .O(n29261));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_in_frame[9] [5]), .I1(n45865), .I2(n28835), 
            .I3(\data_in_frame[9] [4]), .O(n46163));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_891 (.I0(n46107), .I1(\data_in_frame[16] [3]), 
            .I2(n45750), .I3(GND_net), .O(n14_adj_4425));
    defparam i5_3_lut_adj_891.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_892 (.I0(\data_in_frame[16] [2]), .I1(n46260), 
            .I2(n46025), .I3(\data_in_frame[11] [4]), .O(n15_adj_4426));
    defparam i6_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_893 (.I0(n15_adj_4426), .I1(n46163), .I2(n14_adj_4425), 
            .I3(n28776), .O(Kp_23__N_1803));
    defparam i8_4_lut_adj_893.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_894 (.I0(\data_in_frame[13] [4]), .I1(n29105), 
            .I2(n45853), .I3(\data_in_frame[11] [3]), .O(n28861));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_895 (.I0(\data_in_frame[13] [3]), .I1(n4_adj_4427), 
            .I2(n46209), .I3(n46101), .O(n16_adj_4428));
    defparam i6_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_896 (.I0(n46919), .I1(\data_in_frame[11] [0]), 
            .I2(n8_adj_4429), .I3(n43827), .O(n17_adj_4430));
    defparam i7_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_897 (.I0(n17_adj_4430), .I1(n43836), .I2(n16_adj_4428), 
            .I3(n46269), .O(n43800));
    defparam i9_4_lut_adj_897.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45865));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_899 (.I0(\data_in_frame[5] [2]), .I1(n46249), .I2(\data_in_frame[3] [1]), 
            .I3(GND_net), .O(n45764));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_899.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46269));
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_in_frame[16] [3]), .I1(n48165), 
            .I2(GND_net), .I3(GND_net), .O(n46008));
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_902 (.I0(\data_in_frame[10] [7]), .I1(n43827), 
            .I2(GND_net), .I3(GND_net), .O(n46011));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_903 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n46030));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_904 (.I0(\data_in_frame[9] [2]), .I1(n29210), .I2(n28776), 
            .I3(GND_net), .O(n45853));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_904.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_905 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[11] [4]), 
            .I2(n46014), .I3(n46160), .O(n8_adj_4431));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_905.LUT_INIT = 16'h9669;
    SB_LUT4 mux_2021_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n7004));
    defparam mux_2021_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_3_lut (.I0(\data_in_frame[16] [0]), .I1(n8_adj_4431), .I2(n45853), 
            .I3(GND_net), .O(n29195));   // verilog/coms.v(75[16:43])
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_in_frame[18] [0]), .I1(n28861), 
            .I2(GND_net), .I3(GND_net), .O(n46042));
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(CLK_c), 
           .D(n52967));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_907 (.I0(n46042), .I1(\data_in_frame[15] [7]), 
            .I2(n29195), .I3(\data_in_frame[15] [6]), .O(n46219));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_908 (.I0(\data_in_frame[9] [2]), .I1(n47604), 
            .I2(n46030), .I3(n42975), .O(n72));
    defparam i25_4_lut_adj_908.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45913));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i31_4_lut (.I0(n46166), .I1(n46011), .I2(n46036), .I3(n45996), 
            .O(n78));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34554_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50188));
    defparam i34554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35631_2_lut (.I0(n52921), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51136));
    defparam i35631_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n40521), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29_4_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[7] [5]), 
            .I2(Kp_23__N_1321), .I3(\data_in_frame[13] [0]), .O(n76));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34509_4_lut (.I0(byte_transmit_counter[0]), .I1(n51136), .I2(byte_transmit_counter[3]), 
            .I3(\data_out_frame[20] [5]), .O(n50143));
    defparam i34509_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i30_4_lut (.I0(\data_in_frame[17] [3]), .I1(n46282), .I2(\data_in_frame[16] [5]), 
            .I3(n46266), .O(n77));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i20_3_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\data_out_frame[23] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4432));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3971_3 (.CI(n40521), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n40522));
    SB_LUT4 i28_4_lut (.I0(n46008), .I1(n45724), .I2(n45913), .I3(\data_in_frame[10] [1]), 
            .O(n75));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(\data_in_frame[17] [4]), .I1(n46269), .I2(\data_in_frame[18] [1]), 
            .I3(n46064), .O(n74));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34555_4_lut (.I0(n50188), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50189));
    defparam i34555_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i26_4_lut (.I0(n46216), .I1(\data_in_frame[7] [4]), .I2(n45987), 
            .I3(n47973), .O(n73));
    defparam i26_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i43_4_lut (.I0(n75), .I1(n77), .I2(n76), .I3(n78), .O(n90));
    defparam i43_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34553_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50187));
    defparam i34553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36_4_lut (.I0(n43017), .I1(n72), .I2(n10_adj_4433), .I3(n46285), 
            .O(n83));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2021_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n7005));
    defparam mux_2021_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i35_4_lut (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(n42954), .O(n82));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n42873), .I1(\data_in_frame[15] [1]), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[13] [6]), .O(n80));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34_4_lut (.I0(n29188), .I1(\data_in_frame[11] [7]), .I2(n43915), 
            .I3(\data_in_frame[17] [2]), .O(n81));
    defparam i34_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i32_4_lut (.I0(n45961), .I1(n45764), .I2(n45865), .I3(\data_in_frame[3] [0]), 
            .O(n79));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34497_4_lut (.I0(n52747), .I1(n50144), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n50131));
    defparam i34497_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i45_4_lut (.I0(n83), .I1(n90), .I2(n73), .I3(n74), .O(n92));
    defparam i45_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [5]), .I3(\data_in_frame[19] [2]), .O(n6_adj_4434));   // verilog/coms.v(85[17:28])
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i44_4_lut (.I0(n79), .I1(n81), .I2(n80), .I3(n82), .O(n91));
    defparam i44_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34496_3_lut (.I0(n7), .I1(n52843), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n50130));
    defparam i34496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34498_3_lut (.I0(n50130), .I1(n50131), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[5]));
    defparam i34498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3513), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut_adj_910 (.I0(n47090), .I1(n47108), .I2(n47097), 
            .I3(n47333), .O(n29));
    defparam i11_4_lut_adj_910.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[19] [7]), .I3(GND_net), .O(n5_adj_4435));   // verilog/coms.v(85[17:28])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_2021_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n7006));
    defparam mux_2021_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_911 (.I0(n5_adj_4435), .I1(n91), .I2(n6_adj_4434), 
            .I3(n92), .O(n10_adj_4436));
    defparam i3_4_lut_adj_911.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_912 (.I0(\data_in_frame[17] [5]), .I1(n43800), 
            .I2(\data_in_frame[15] [4]), .I3(n45718), .O(n43017));
    defparam i1_4_lut_adj_912.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_913 (.I0(n45706), .I1(n46196), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4437));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i35686_2_lut (.I0(n52915), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51134));
    defparam i35686_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34512_4_lut (.I0(byte_transmit_counter[0]), .I1(n51134), .I2(byte_transmit_counter[3]), 
            .I3(\data_out_frame[20] [6]), .O(n50146));
    defparam i34512_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i20_3_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\data_out_frame[23] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4438));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_914 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[14] [7]), 
            .I2(n46089), .I3(n6_adj_4437), .O(n29255));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n43889), .I1(n27975), .I2(n43795), .I3(n29255), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_915 (.I0(n43017), .I1(n12), .I2(n10_adj_4436), 
            .I3(n46219), .O(n45885));
    defparam i6_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_916 (.I0(n43836), .I1(\data_in_frame[10] [7]), 
            .I2(n8_adj_4429), .I3(n43827), .O(n46919));
    defparam i3_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_917 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4439));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h6666;
    SB_LUT4 i34561_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n50195));
    defparam i34561_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i4_4_lut_adj_918 (.I0(n28674), .I1(n46919), .I2(\data_in_frame[11] [1]), 
            .I3(n6_adj_4439), .O(n45724));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_918.LUT_INIT = 16'h9669;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3513), 
            .CO(n40521));
    SB_LUT4 i34559_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50193));
    defparam i34559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_919 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46101));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_920 (.I0(n28809), .I1(n46101), .I2(n45724), .I3(\data_in_frame[10] [5]), 
            .O(n42975));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46285));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_922 (.I0(n42975), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45718));
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h6666;
    SB_LUT4 i34503_4_lut (.I0(n52777), .I1(n50147), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n50137));
    defparam i34503_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34502_3_lut (.I0(n7_adj_4440), .I1(n52837), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n50136));
    defparam i34502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34504_3_lut (.I0(n50136), .I1(n50137), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[6]));
    defparam i34504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_923 (.I0(Kp_23__N_1195), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[11] [0]), .I3(n6_adj_4441), .O(n46089));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_924 (.I0(n46240), .I1(n46089), .I2(\data_in_frame[17] [4]), 
            .I3(n45718), .O(n10_adj_4442));
    defparam i4_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46092));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4443));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_927 (.I0(n28674), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [7]), .I3(n6_adj_4443), .O(n45706));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_928 (.I0(n28892), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46240));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46216));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_930 (.I0(\data_in_frame[10] [2]), .I1(n42873), 
            .I2(n46020), .I3(n28827), .O(n42988));
    defparam i3_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_931 (.I0(n46203), .I1(n42988), .I2(\data_in_frame[16] [6]), 
            .I3(n46216), .O(n12_adj_4444));
    defparam i5_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_932 (.I0(n42892), .I1(n12_adj_4444), .I2(\data_in_frame[14] [4]), 
            .I3(n45999), .O(n43606));
    defparam i6_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i35689_2_lut (.I0(n52909), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51132));
    defparam i35689_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34515_4_lut (.I0(\data_out_frame[20] [7]), .I1(n51132), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[0]), .O(n50149));
    defparam i34515_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_933 (.I0(n43606), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43915));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_934 (.I0(n45706), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4445));
    defparam i2_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_935 (.I0(n46092), .I1(n42988), .I2(\data_in_frame[14] [6]), 
            .I3(\data_in_frame[15] [0]), .O(n14_adj_4446));
    defparam i6_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_936 (.I0(\data_in_frame[17] [2]), .I1(n14_adj_4446), 
            .I2(n10_adj_4445), .I3(n4_adj_4427), .O(n43795));
    defparam i7_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i20_3_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\data_out_frame[23] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4447));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34570_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n50204));
    defparam i34570_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34568_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50202));
    defparam i34568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34506_4_lut (.I0(n52783), .I1(n50150), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n50140));
    defparam i34506_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34505_3_lut (.I0(n7_adj_4448), .I1(n52825), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n50139));
    defparam i34505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34507_3_lut (.I0(n50139), .I1(n50140), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[7]));
    defparam i34507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n46279));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_938 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n46193));
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_939 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n46273));
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_940 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4449));
    defparam i2_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_941 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[8] [0]), 
            .I2(n45875), .I3(\data_in_frame[1] [4]), .O(n14_adj_4450));
    defparam i6_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_942 (.I0(\data_in_frame[10] [1]), .I1(n14_adj_4450), 
            .I2(n10_adj_4449), .I3(n46166), .O(n46225));
    defparam i7_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_943 (.I0(\data_in_frame[12] [3]), .I1(n46225), 
            .I2(\data_in_frame[14] [5]), .I3(GND_net), .O(n45973));
    defparam i2_3_lut_adj_943.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_944 (.I0(\data_in_frame[10] [3]), .I1(n46184), 
            .I2(n45715), .I3(\data_in_frame[8] [1]), .O(n10_adj_4451));   // verilog/coms.v(96[12:25])
    defparam i4_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_945 (.I0(n45910), .I1(n10_adj_4451), .I2(\data_in_frame[7] [7]), 
            .I3(GND_net), .O(n46196));   // verilog/coms.v(96[12:25])
    defparam i5_3_lut_adj_945.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_946 (.I0(n43430), .I1(n46049), .I2(\data_in_frame[12] [2]), 
            .I3(n42921), .O(n12_adj_4452));
    defparam i5_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2021_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n7007));
    defparam mux_2021_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_947 (.I0(n46279), .I1(n12_adj_4452), .I2(\data_in_frame[14] [3]), 
            .I3(n46225), .O(n48165));
    defparam i6_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_948 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n45930));
    defparam i2_3_lut_adj_948.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_949 (.I0(n48165), .I1(n46196), .I2(n45973), .I3(\data_in_frame[12] [4]), 
            .O(n43899));
    defparam i3_4_lut_adj_949.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_950 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(n46273), .I3(\data_in_frame[17] [1]), .O(n6_adj_4453));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_951 (.I0(n45973), .I1(Kp_23__N_1285), .I2(n46193), 
            .I3(n6_adj_4453), .O(n47973));
    defparam i4_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_952 (.I0(n43430), .I1(n29226), .I2(GND_net), 
            .I3(GND_net), .O(n46014));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29505));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2021_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n7008));
    defparam mux_2021_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2021_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n7009));
    defparam mux_2021_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_954 (.I0(\data_in_frame[7] [7]), .I1(n29268), .I2(n46054), 
            .I3(n6_adj_4454), .O(n42873));   // verilog/coms.v(96[12:25])
    defparam i4_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2021_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n7010));
    defparam mux_2021_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_adj_955 (.I0(n28809), .I1(n4_adj_4427), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1285));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_33_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n40520), .O(n2_adj_4455)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_956 (.I0(n29226), .I1(n29210), .I2(GND_net), 
            .I3(GND_net), .O(n45944));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_957 (.I0(n46257), .I1(n28674), .I2(n45944), .I3(Kp_23__N_1285), 
            .O(n14_adj_4456));
    defparam i6_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_958 (.I0(n42873), .I1(n14_adj_4456), .I2(n10_adj_4457), 
            .I3(n45936), .O(n43827));
    defparam i7_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_959 (.I0(n28674), .I1(\data_in_frame[9] [0]), .I2(n43827), 
            .I3(GND_net), .O(n43836));
    defparam i1_3_lut_adj_959.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_960 (.I0(n43836), .I1(n28565), .I2(\data_in_frame[9] [5]), 
            .I3(n6_adj_4458), .O(n43811));
    defparam i4_4_lut_adj_960.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_961 (.I0(\data_in_frame[8] [6]), .I1(n8_adj_4429), 
            .I2(GND_net), .I3(GND_net), .O(n28815));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_962 (.I0(n29), .I1(n34), .I2(n50027), .I3(n24_adj_4459), 
            .O(n54_c));
    defparam i17_4_lut_adj_962.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_963 (.I0(Kp_23__N_1195), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n46036));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_964 (.I0(n28776), .I1(\data_in_frame[9] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n46209));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_32_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n40519), .O(n2_adj_4460)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_965 (.I0(\data_in_frame[8] [0]), .I1(n42655), .I2(n46036), 
            .I3(\data_in_frame[8] [3]), .O(n18_adj_4461));
    defparam i7_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_966 (.I0(n46136), .I1(n28815), .I2(\data_in_frame[8] [1]), 
            .I3(n43811), .O(n19_adj_4462));
    defparam i8_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_967 (.I0(n19_adj_4462), .I1(n45991), .I2(n18_adj_4461), 
            .I3(n12_adj_4463), .O(n47604));
    defparam i10_4_lut_adj_967.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_968 (.I0(\data_in_frame[9] [0]), .I1(n47604), .I2(\data_in_frame[7] [7]), 
            .I3(\data_in_frame[12] [0]), .O(n46228));
    defparam i3_4_lut_adj_968.LUT_INIT = 16'h9669;
    SB_CARRY add_43_32 (.CI(n40519), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n40520));
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46049));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_970 (.I0(\data_in_frame[13] [7]), .I1(n45827), 
            .I2(n46049), .I3(\data_in_frame[11] [5]), .O(n14_adj_4464));
    defparam i6_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_971 (.I0(\data_in_frame[14] [1]), .I1(n14_adj_4464), 
            .I2(n10_adj_4465), .I3(n46228), .O(n46107));
    defparam i7_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28565));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_973 (.I0(n28776), .I1(n8_adj_4429), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1321));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_adj_973.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_974 (.I0(n45817), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n45955));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_974.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_975 (.I0(n28776), .I1(n43430), .I2(GND_net), 
            .I3(GND_net), .O(n46257));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_976 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n46160));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_31_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n40518), .O(n2_adj_4466)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_977 (.I0(n46260), .I1(\data_in_frame[9] [4]), .I2(n46160), 
            .I3(\data_in_frame[15] [7]), .O(n14_adj_4467));
    defparam i6_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_978 (.I0(\data_in_frame[16] [1]), .I1(n46257), 
            .I2(n45955), .I3(\data_in_frame[16] [2]), .O(n13));
    defparam i5_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_979 (.I0(\data_in_frame[18] [3]), .I1(n13), .I2(n14_adj_4467), 
            .I3(GND_net), .O(n45987));
    defparam i1_3_lut_adj_979.LUT_INIT = 16'h6969;
    SB_LUT4 i34604_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50238));
    defparam i34604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34605_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50239));
    defparam i34605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34608_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50242));
    defparam i34608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34607_3_lut (.I0(\data_out_frame[20]_c [4]), .I1(\data_out_frame[21][4] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50241));
    defparam i34607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34643_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50277));
    defparam i34643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34644_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50278));
    defparam i34644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34647_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50281));
    defparam i34647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34646_3_lut (.I0(\data_out_frame[20][1] ), .I1(\data_out_frame[21][1] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50280));
    defparam i34646_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n29645), .D(n8825[0]), .R(n39711));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i34622_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50256));
    defparam i34622_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_31 (.CI(n40518), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n40519));
    SB_LUT4 i34623_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50257));
    defparam i34623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34635_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50269));
    defparam i34635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34634_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21][2] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50268));
    defparam i34634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2021_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n7011));
    defparam mux_2021_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_980 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [4]), 
            .I2(ID[0]), .I3(ID[4]), .O(n9));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_980.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_981 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [1]), 
            .I2(ID[7]), .I3(ID[1]), .O(n8_adj_4468));
    defparam i2_4_lut_adj_981.LUT_INIT = 16'h7bde;
    SB_LUT4 add_43_30_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n40517), .O(n2_adj_4469)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_982 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[5]), .I3(ID[3]), .O(n7_adj_4470));
    defparam i1_4_lut_adj_982.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_983 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[2]), .I3(ID[6]), .O(n9_adj_4471));
    defparam i3_4_lut_adj_983.LUT_INIT = 16'h7bde;
    SB_LUT4 i5_3_lut_adj_984 (.I0(n9_adj_4471), .I1(n7_adj_4470), .I2(n8_adj_4468), 
            .I3(GND_net), .O(n49));
    defparam i5_3_lut_adj_984.LUT_INIT = 16'hfefe;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n46478), .D(n35937), 
            .R(n36742));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n48237), .D(n29930), 
            .R(n47799));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_985 (.I0(\data_in_frame[4] [3]), .I1(n28791), .I2(\data_in_frame[8] [7]), 
            .I3(n45781), .O(n10_adj_4472));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_986 (.I0(n45795), .I1(n45958), .I2(\data_in_frame[6] [1]), 
            .I3(\data_in_frame[5] [7]), .O(n12_adj_4473));
    defparam i5_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_987 (.I0(\data_in_frame[8] [3]), .I1(n12_adj_4473), 
            .I2(n46130), .I3(\data_in_frame[6] [2]), .O(n28809));
    defparam i6_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_988 (.I0(n29147), .I1(\data_in_frame[4] [4]), .I2(\data_in_frame[6] [6]), 
            .I3(\data_in_frame[7] [0]), .O(n14_adj_4474));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_989 (.I0(\data_in_frame[4] [6]), .I1(n14_adj_4474), 
            .I2(n10_adj_4475), .I3(\data_in_frame[6] [7]), .O(n28776));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n45958));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 i3_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/coms.v(78[16:27])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_991 (.I0(\data_in_frame[8] [0]), .I1(Kp_23__N_1020), 
            .I2(\data_in_frame[4] [5]), .I3(n28870), .O(n13_adj_4476));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_992 (.I0(n13_adj_4476), .I1(n11), .I2(n45991), 
            .I3(n45958), .O(n46054));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_992.LUT_INIT = 16'h9669;
    SB_CARRY add_43_30 (.CI(n40517), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n40518));
    SB_LUT4 mux_2021_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[17] [0]), .O(n7012));
    defparam mux_2021_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_adj_993 (.I0(Kp_23__N_1093), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4477));   // verilog/coms.v(78[16:27])
    defparam i2_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_994 (.I0(n28761), .I1(n7_adj_4477), .I2(\data_in_frame[8] [4]), 
            .I3(n8_adj_4478), .O(n4_adj_4427));   // verilog/coms.v(74[16:43])
    defparam i2_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_in_frame[4] [7]), .I1(n6_adj_4479), 
            .I2(GND_net), .I3(GND_net), .O(n29223));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_996 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[6] [7]), 
            .I2(n29223), .I3(\data_in_frame[7] [1]), .O(n45916));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_997 (.I0(\data_out_frame[25] [6]), .I1(n28578), 
            .I2(n48160), .I3(n46002), .O(n10_adj_4480));
    defparam i4_4_lut_adj_997.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_998 (.I0(\data_out_frame[23] [6]), .I1(n10_adj_4480), 
            .I2(\data_out_frame[23] [4]), .I3(GND_net), .O(n47661));
    defparam i5_3_lut_adj_998.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_999 (.I0(n43816), .I1(n47627), .I2(\data_out_frame[25] [7]), 
            .I3(GND_net), .O(n46002));
    defparam i2_3_lut_adj_999.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1000 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n46130));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1000.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1001 (.I0(\data_out_frame[24] [0]), .I1(n2134), 
            .I2(n43832), .I3(n6_adj_4481), .O(n47566));
    defparam i4_4_lut_adj_1001.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1002 (.I0(n46061), .I1(n43803), .I2(n48160), 
            .I3(n46181), .O(n10_adj_4482));
    defparam i4_4_lut_adj_1002.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1003 (.I0(n47627), .I1(n10_adj_4482), .I2(n2134), 
            .I3(GND_net), .O(n47422));
    defparam i5_3_lut_adj_1003.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_29_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n40516), .O(n2_adj_4483)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_2021_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n7013));
    defparam mux_2021_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1004 (.I0(\data_out_frame[19] [4]), .I1(n42864), 
            .I2(\data_out_frame[19] [3]), .I3(n47800), .O(n48160));
    defparam i3_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1005 (.I0(\data_in_frame[0] [0]), .I1(n46130), 
            .I2(n45801), .I3(\data_in_frame[2] [1]), .O(Kp_23__N_1093));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1093), 
            .I2(GND_net), .I3(GND_net), .O(n46136));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2021_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n7014));
    defparam mux_2021_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_43_29 (.CI(n40516), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n40517));
    SB_LUT4 i2_3_lut_adj_1007 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n46282));
    defparam i2_3_lut_adj_1007.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29268));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(n48160), .I1(\data_out_frame[23] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43832));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n29481), .I1(\data_out_frame[24] [1]), 
            .I2(n43832), .I3(n46046), .O(n10_adj_4484));
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1011 (.I0(n47041), .I1(n10_adj_4484), .I2(\data_out_frame[22] [1]), 
            .I3(GND_net), .O(n48100));
    defparam i5_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1012 (.I0(\data_out_frame[19] [5]), .I1(n45841), 
            .I2(\data_out_frame[19] [4]), .I3(\data_out_frame[17] [4]), 
            .O(n12_adj_4485));
    defparam i5_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1013 (.I0(\data_out_frame[17] [2]), .I1(n12_adj_4485), 
            .I2(n46148), .I3(n29389), .O(n2134));
    defparam i6_4_lut_adj_1013.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45733));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_28_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n40515), .O(n2_adj_4486)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_out_frame[24] [2]), .I1(n2134), 
            .I2(GND_net), .I3(GND_net), .O(n46046));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_CARRY add_43_28 (.CI(n40515), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n40516));
    SB_LUT4 i5_4_lut_adj_1016 (.I0(\data_out_frame[20][1] ), .I1(n46046), 
            .I2(\data_out_frame[24] [3]), .I3(n43906), .O(n12_adj_4487));
    defparam i5_4_lut_adj_1016.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1017 (.I0(n43803), .I1(n12_adj_4487), .I2(n46222), 
            .I3(n48133), .O(n47769));
    defparam i6_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1018 (.I0(\data_out_frame[20]_c [4]), .I1(n46033), 
            .I2(n28003), .I3(n43906), .O(n12_adj_4488));
    defparam i5_4_lut_adj_1018.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1019 (.I0(n47041), .I1(n12_adj_4488), .I2(n46095), 
            .I3(\data_out_frame[24] [4]), .O(n46928));
    defparam i6_4_lut_adj_1019.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1020 (.I0(n43860), .I1(n43038), .I2(\data_out_frame[22] [4]), 
            .I3(\data_out_frame[20][1] ), .O(n10_adj_4489));
    defparam i4_4_lut_adj_1020.LUT_INIT = 16'h9669;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n29629), .D(n7019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n29629), .D(n7018));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n29629), .D(n7017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n29629), .D(n7016));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n29629), .D(n7015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n29629), .D(n7014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n29629), .D(n7013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n29629), .D(n7012));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n29629), .D(n7011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n29629), .D(n7010));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n29629), .D(n7009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n29629), .D(n7008));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n29629), .D(n7007));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n29629), .D(n7006));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n29629), .D(n7005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n29629), .D(n7004));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n29629), .D(n7003));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n29629), .D(n7002));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n29629), .D(n7001));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n29629), .D(n7000));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n29629), .D(n6999));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n29629), .D(n6998));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n29629), .D(n6997));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1021 (.I0(n45721), .I1(n46098), .I2(n28003), 
            .I3(n45676), .O(n15_adj_4490));
    defparam i6_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2021_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n7015));
    defparam mux_2021_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1022 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [4]), 
            .I2(\data_in_frame[5] [3]), .I3(n6_adj_4491), .O(n45875));
    defparam i4_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1023 (.I0(n15_adj_4490), .I1(n28663), .I2(n14_adj_4492), 
            .I3(\data_out_frame[24] [6]), .O(n47644));
    defparam i8_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1024 (.I0(n45733), .I1(n45952), .I2(n46184), 
            .I3(n46266), .O(n28892));
    defparam i3_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1025 (.I0(\data_out_frame[20][1] ), .I1(\data_out_frame[20] [2]), 
            .I2(\data_out_frame[20]_c [4]), .I3(GND_net), .O(n45721));
    defparam i2_3_lut_adj_1025.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(n45721), .I1(n46095), .I2(GND_net), 
            .I3(GND_net), .O(n29481));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1027 (.I0(n45821), .I1(n46136), .I2(\data_in_frame[8] [5]), 
            .I3(GND_net), .O(n28674));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1027.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1028 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[22] [1]), 
            .I2(\data_out_frame[22] [3]), .I3(GND_net), .O(n46033));
    defparam i2_3_lut_adj_1028.LUT_INIT = 16'h9696;
    SB_LUT4 equal_2184_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4433));   // verilog/coms.v(166[9:87])
    defparam equal_2184_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45952));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\data_out_frame[24] [4]), .I1(n48133), 
            .I2(GND_net), .I3(GND_net), .O(n43860));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(n28870), .I1(n45910), .I2(GND_net), 
            .I3(GND_net), .O(n28981));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_988), .I3(\data_in_frame[0] [5]), .O(n28977));
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n46249));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(CLK_c), 
            .D(n45580), .S(n44886));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\data_in_frame[3] [2]), .I1(n45830), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4493));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1035 (.I0(\data_out_frame[17] [6]), .I1(n29389), 
            .I2(n45696), .I3(n42909), .O(n14_adj_4494));
    defparam i6_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1036 (.I0(n28990), .I1(n14_adj_4494), .I2(n10_adj_4495), 
            .I3(\data_out_frame[19] [7]), .O(n45777));
    defparam i7_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1037 (.I0(n6_adj_4496), .I1(n29502), .I2(\data_out_frame[17] [3]), 
            .I3(n29529), .O(n10_adj_4497));
    defparam i4_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1038 (.I0(\data_out_frame[15] [1]), .I1(n10_adj_4497), 
            .I2(\data_out_frame[15] [2]), .I3(GND_net), .O(n42864));
    defparam i5_3_lut_adj_1038.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1039 (.I0(\data_in_frame[7] [4]), .I1(n27216), 
            .I2(n28977), .I3(n6_adj_4493), .O(n46139));
    defparam i4_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1040 (.I0(n42864), .I1(\data_out_frame[17] [5]), 
            .I2(n45777), .I3(\data_out_frame[19] [5]), .O(n10_adj_4498));
    defparam i4_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1041 (.I0(n29171), .I1(n10_adj_4498), .I2(n45862), 
            .I3(GND_net), .O(n43803));
    defparam i5_3_lut_adj_1041.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(n46139), .I1(n46249), .I2(GND_net), 
            .I3(GND_net), .O(n28835));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\data_in_frame[7] [7]), .I1(n42954), 
            .I2(GND_net), .I3(GND_net), .O(n46020));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_in_frame[4] [5]), .I1(n28750), 
            .I2(GND_net), .I3(GND_net), .O(n46124));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n45689));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1046 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n28750));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1046.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_out_frame[13] [1]), .I1(n27979), 
            .I2(GND_net), .I3(GND_net), .O(n29529));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29134));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n45693));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45767));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45859));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_in_frame[2] [1]), .I1(n29137), 
            .I2(GND_net), .I3(GND_net), .O(n28702));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1053 (.I0(\data_in_frame[0] [5]), .I1(n45859), 
            .I2(n45767), .I3(n45693), .O(Kp_23__N_969));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1054 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n46142));
    defparam i2_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1055 (.I0(n45862), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[17] [5]), .I3(n45967), .O(n10_adj_4499));
    defparam i4_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1056 (.I0(\data_out_frame[19] [7]), .I1(n10_adj_4499), 
            .I2(\data_out_frame[18] [0]), .I3(GND_net), .O(n43906));
    defparam i5_3_lut_adj_1056.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\data_out_frame[24] [5]), .I1(n43906), 
            .I2(GND_net), .I3(GND_net), .O(n45676));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45919));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46181));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1060 (.I0(n28997), .I1(n45729), .I2(n46071), 
            .I3(\data_out_frame[5] [7]), .O(n16_adj_4500));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1061 (.I0(\data_out_frame[12] [7]), .I1(n45678), 
            .I2(n46104), .I3(\data_out_frame[10] [7]), .O(n17_adj_4501));   // verilog/coms.v(85[17:70])
    defparam i7_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1062 (.I0(n17_adj_4501), .I1(\data_out_frame[11] [0]), 
            .I2(n16_adj_4500), .I3(n4_adj_4502), .O(n27979));   // verilog/coms.v(85[17:70])
    defparam i9_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n46187), .I1(n45787), .I2(n45983), .I3(n45673), 
            .O(n62_adj_4503));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2021_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n7016));
    defparam mux_2021_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_4_lut_adj_1063 (.I0(n27979), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[18] [1]), .I3(\data_out_frame[20] [6]), 
            .O(n12_adj_4504));
    defparam i5_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1064 (.I0(\data_out_frame[22] [5]), .I1(n46181), 
            .I2(n45907), .I3(\data_out_frame[23] [7]), .O(n47414));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28761));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1066 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n45961));
    defparam i2_3_lut_adj_1066.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28741));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[14] [4]), .I1(n43910), .I2(n42909), 
            .I3(n45784), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1068 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[5] [7]), .O(n45715));   // verilog/coms.v(96[12:25])
    defparam i3_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1069 (.I0(n45729), .I1(\data_out_frame[5] [7]), 
            .I2(n43007), .I3(n29171), .O(n26));
    defparam i10_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1070 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[8] [3]), .I3(n29529), .O(n27));
    defparam i11_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1071 (.I0(n43846), .I1(n43805), .I2(n1563), .I3(n45752), 
            .O(n25));
    defparam i9_4_lut_adj_1071.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1072 (.I0(n46246), .I1(n28941), .I2(n29044), 
            .I3(\data_out_frame[14] [6]), .O(n10_adj_4505));
    defparam i4_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28791));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n29164));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_27_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n40514), .O(n2_adj_4506)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_adj_1075 (.I0(\data_out_frame[14] [7]), .I1(n10_adj_4505), 
            .I2(n46263), .I3(GND_net), .O(n48327));
    defparam i5_3_lut_adj_1075.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1076 (.I0(\data_in_frame[3] [0]), .I1(n26683), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[5] [3]), .O(n45830));
    defparam i3_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1077 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [1]), 
            .I2(n45830), .I3(\data_in_frame[3] [4]), .O(n40_adj_4507));
    defparam i16_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1078 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n48347));
    defparam i15_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1079 (.I0(\data_in_frame[6] [7]), .I1(n29164), 
            .I2(n28791), .I3(\data_in_frame[3] [3]), .O(n38_adj_4508));
    defparam i14_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1080 (.I0(n28595), .I1(\data_in_frame[3] [6]), 
            .I2(n45715), .I3(n28741), .O(n39_adj_4509));
    defparam i15_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n28761), .I1(\data_in_frame[6] [1]), .I2(n46142), 
            .I3(\data_in_frame[6] [4]), .O(n37));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1081 (.I0(n45872), .I1(Kp_23__N_969), .I2(n28702), 
            .I3(n29147), .O(n42_adj_4510));
    defparam i18_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39_adj_4509), .I2(n38_adj_4508), 
            .I3(n40_adj_4507), .O(n46_c));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1082 (.I0(n29134), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [7]), .I3(Kp_23__N_1020), .O(n41_adj_4511));
    defparam i17_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1083 (.I0(\data_in_frame[3] [5]), .I1(n45689), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[8] [1]), .O(n46077));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45781));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4512));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1086 (.I0(n29147), .I1(\data_in_frame[2] [0]), 
            .I2(n45801), .I3(n6_adj_4512), .O(n45821));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_in_frame[0] [0]), .I1(n45821), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4513));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1088 (.I0(n48347), .I1(n46119), .I2(n48327), 
            .I3(n46127), .O(n12_adj_4514));
    defparam i5_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n46213), .I1(\data_out_frame[24] [2]), .I2(\data_out_frame[15] [3]), 
            .I3(n46058), .O(n60));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1089 (.I0(n45919), .I1(n12_adj_4514), .I2(n45893), 
            .I3(n45841), .O(n48336));
    defparam i6_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut_adj_1090 (.I0(n43_adj_4515), .I1(n62_adj_4503), .I2(\data_out_frame[19] [4]), 
            .I3(n45674), .O(n70));
    defparam i31_4_lut_adj_1090.LUT_INIT = 16'h9669;
    SB_LUT4 i29_4_lut_adj_1091 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[19] [7]), 
            .I2(n47706), .I3(n43803), .O(n68));
    defparam i29_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1092 (.I0(n42936), .I1(n60), .I2(n43860), .I3(n45939), 
            .O(n69));
    defparam i30_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1093 (.I0(\data_in_frame[6] [5]), .I1(n29164), 
            .I2(n45758), .I3(n6_adj_4513), .O(Kp_23__N_1195));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(n43430), .I1(Kp_23__N_1195), .I2(\data_in_frame[8] [6]), 
            .I3(GND_net), .O(n25_adj_4516));
    defparam i8_3_lut.LUT_INIT = 16'h7d7d;
    SB_LUT4 i28_4_lut_adj_1094 (.I0(\data_out_frame[16] [4]), .I1(n45676), 
            .I2(n48336), .I3(n42930), .O(n67_adj_4517));
    defparam i28_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1095 (.I0(\data_out_frame[22] [4]), .I1(n11_adj_4518), 
            .I2(n47414), .I3(n12_adj_4504), .O(n48));
    defparam i9_4_lut_adj_1095.LUT_INIT = 16'h9669;
    SB_LUT4 i25_4_lut_adj_1096 (.I0(\data_out_frame[25] [7]), .I1(n46206), 
            .I2(\data_out_frame[18] [4]), .I3(n46061), .O(n64));
    defparam i25_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_1097 (.I0(n45696), .I1(n42898), .I2(\data_out_frame[16] [2]), 
            .I3(\data_out_frame[16] [7]), .O(n66));
    defparam i27_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1098 (.I0(\data_in_frame[3] [6]), .I1(n29137), 
            .I2(n46124), .I3(n6_adj_4519), .O(n47199));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1099 (.I0(n25_adj_4516), .I1(n46020), .I2(n29226), 
            .I3(n28835), .O(n30));
    defparam i13_4_lut_adj_1099.LUT_INIT = 16'hfbff;
    SB_LUT4 i26_4_lut_adj_1100 (.I0(n46033), .I1(n45881), .I2(n45970), 
            .I3(n45755), .O(n65));
    defparam i26_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1101 (.I0(n29210), .I1(n28674), .I2(n28892), 
            .I3(n42921), .O(n28_adj_4520));
    defparam i11_4_lut_adj_1101.LUT_INIT = 16'hfffe;
    SB_LUT4 i37_4_lut (.I0(n67_adj_4517), .I1(n69), .I2(n68), .I3(n70), 
            .O(n76_adj_4521));
    defparam i37_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1102 (.I0(n4_adj_4427), .I1(n28827), .I2(n47199), 
            .I3(n46054), .O(n29_adj_4522));
    defparam i12_4_lut_adj_1102.LUT_INIT = 16'hfbff;
    SB_LUT4 i32_4_lut_adj_1103 (.I0(n29481), .I1(n64), .I2(n48), .I3(n43007), 
            .O(n71));
    defparam i32_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1104 (.I0(n28776), .I1(n28809), .I2(n8_adj_4429), 
            .I3(n61), .O(n27_adj_4523));
    defparam i10_4_lut_adj_1104.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1105 (.I0(n27_adj_4523), .I1(n29_adj_4522), .I2(n28_adj_4520), 
            .I3(n30), .O(n62));
    defparam i16_4_lut_adj_1105.LUT_INIT = 16'hfffe;
    SB_LUT4 i38_4_lut (.I0(n71), .I1(n76_adj_4521), .I2(n65), .I3(n66), 
            .O(n47698));
    defparam i38_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24283_3_lut (.I0(n54_c), .I1(n62), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n63_c));   // verilog/coms.v(112[11:16])
    defparam i24283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(n47698), .I1(n43858), .I2(GND_net), 
            .I3(GND_net), .O(n43834));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i37075_4_lut (.I0(n63_c), .I1(n45635), .I2(n32424), .I3(\FRAME_MATCHER.state[2] ), 
            .O(n29629));
    defparam i37075_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_2021_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n7017));
    defparam mux_2021_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1107 (.I0(n45761), .I1(n46112), .I2(\data_out_frame[9] [0]), 
            .I3(n29034), .O(n15_adj_4524));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1108 (.I0(n15_adj_4524), .I1(\data_out_frame[4] [0]), 
            .I2(n14_adj_4525), .I3(\data_out_frame[8] [5]), .O(n29389));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_CARRY add_43_27 (.CI(n40514), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n40515));
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_out_frame[17] [6]), .I1(n27987), 
            .I2(GND_net), .I3(GND_net), .O(n42936));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(n29389), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4526));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1111 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n43007), .I3(GND_net), .O(n45967));
    defparam i2_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1112 (.I0(n29171), .I1(n7_adj_4526), .I2(n42936), 
            .I3(n8_adj_4527), .O(n47706));
    defparam i5_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1113 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n45907));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1114 (.I0(n47706), .I1(\data_out_frame[18] [0]), 
            .I2(n43975), .I3(GND_net), .O(n28003));
    defparam i2_3_lut_adj_1114.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1115 (.I0(n48169), .I1(n28003), .I2(n43038), 
            .I3(GND_net), .O(n10_adj_4528));
    defparam i3_3_lut_adj_1115.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1116 (.I0(n45674), .I1(n45907), .I2(n28663), 
            .I3(n25_adj_4529), .O(n11_adj_4530));
    defparam i4_4_lut_adj_1116.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1117 (.I0(n11_adj_4530), .I1(\data_out_frame[22] [4]), 
            .I2(n10_adj_4528), .I3(\data_out_frame[25] [0]), .O(n43858));
    defparam i6_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(n43858), .I1(n45881), .I2(GND_net), 
            .I3(GND_net), .O(n45882));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1119 (.I0(n42894), .I1(n45947), .I2(\data_out_frame[22] [6]), 
            .I3(\data_out_frame[22] [7]), .O(n45673));
    defparam i3_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(n46157), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[13] [3]), .I3(n46253), .O(n10_adj_4531));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1121 (.I0(n45850), .I1(n10_adj_4531), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n29171));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1122 (.I0(n42875), .I1(n46005), .I2(n29171), 
            .I3(\data_out_frame[15] [5]), .O(n12_adj_4532));
    defparam i5_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1123 (.I0(\data_out_frame[18] [1]), .I1(n43854), 
            .I2(n12_adj_4532), .I3(n8_adj_4533), .O(n43975));
    defparam i1_4_lut_adj_1123.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1124 (.I0(\data_out_frame[20]_c [4]), .I1(n45673), 
            .I2(n28663), .I3(n48169), .O(n45674));
    defparam i3_4_lut_adj_1124.LUT_INIT = 16'h9669;
    SB_LUT4 i36361_2_lut (.I0(n45674), .I1(\data_out_frame[23] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n51996));   // verilog/coms.v(97[12:26])
    defparam i36361_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1125 (.I0(n45933), .I1(n28663), .I2(\data_out_frame[24] [7]), 
            .I3(n46098), .O(n10_adj_4534));
    defparam i4_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1126 (.I0(\data_out_frame[25] [1]), .I1(n42894), 
            .I2(n10_adj_4534), .I3(n51996), .O(n45881));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(n47476), .I1(n45881), .I2(\data_out_frame[25] [2]), 
            .I3(GND_net), .O(n46908));
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4502));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1129 (.I0(\data_out_frame[8] [7]), .I1(n4_adj_4502), 
            .I2(\data_out_frame[11] [2]), .I3(n6_adj_4535), .O(n45850));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(n45850), .I1(n46175), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4536));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(\data_out_frame[9] [0]), .I1(n29296), 
            .I2(n46154), .I3(n6_adj_4536), .O(n27987));
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[13] [4]), .I1(n27987), 
            .I2(GND_net), .I3(GND_net), .O(n28990));
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(n46112), .I1(n46145), .I2(\data_out_frame[13] [6]), 
            .I3(\data_out_frame[9] [2]), .O(n10_adj_4537));
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1134 (.I0(\data_out_frame[15] [6]), .I1(n42930), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n8_adj_4538));   // verilog/coms.v(71[16:27])
    defparam i3_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1135 (.I0(\data_out_frame[18] [2]), .I1(n46005), 
            .I2(n8_adj_4538), .I3(\data_out_frame[15] [7]), .O(n45947));
    defparam i1_4_lut_adj_1135.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45933));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45787));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1138 (.I0(n45856), .I1(n45933), .I2(\data_out_frame[23] [1]), 
            .I3(\data_out_frame[23] [0]), .O(n12_adj_4539));
    defparam i5_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1139 (.I0(\data_out_frame[21][0] ), .I1(n12_adj_4539), 
            .I2(n45947), .I3(\data_out_frame[20]_c [4]), .O(n47476));
    defparam i6_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1140 (.I0(n47476), .I1(n45787), .I2(n26646), 
            .I3(GND_net), .O(n47315));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1141 (.I0(n46145), .I1(\data_out_frame[11] [3]), 
            .I2(n28997), .I3(GND_net), .O(n46154));
    defparam i3_3_lut_adj_1141.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1142 (.I0(\data_out_frame[9] [3]), .I1(n46154), 
            .I2(\data_out_frame[8] [7]), .I3(n45770), .O(n12_adj_4540));
    defparam i5_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1143 (.I0(\data_out_frame[9] [1]), .I1(n12_adj_4540), 
            .I2(\data_out_frame[13] [5]), .I3(n46115), .O(n43007));
    defparam i6_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1144 (.I0(\data_out_frame[14] [0]), .I1(n28719), 
            .I2(n43007), .I3(n46039), .O(n10_adj_4541));
    defparam i4_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1145 (.I0(\data_out_frame[11] [6]), .I1(n10_adj_4541), 
            .I2(n28127), .I3(GND_net), .O(n43846));
    defparam i5_3_lut_adj_1145.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1146 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n43846), .I3(GND_net), .O(n47174));
    defparam i2_3_lut_adj_1146.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4529));   // verilog/coms.v(97[12:26])
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1148 (.I0(n25_adj_4529), .I1(n29020), .I2(n28663), 
            .I3(n45939), .O(n10_adj_4542));
    defparam i4_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1149 (.I0(\data_out_frame[21][1] ), .I1(n10_adj_4542), 
            .I2(\data_out_frame[23] [2]), .I3(GND_net), .O(n26646));
    defparam i5_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1150 (.I0(\data_out_frame[25] [3]), .I1(n45983), 
            .I2(n26646), .I3(GND_net), .O(n48173));
    defparam i2_3_lut_adj_1150.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_adj_1151 (.I0(\data_out_frame[9] [2]), .I1(n4_adj_4543), 
            .I2(GND_net), .I3(GND_net), .O(n29296));
    defparam i2_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(n29458), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46115));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1153 (.I0(n46115), .I1(\data_out_frame[14] [1]), 
            .I2(n29296), .I3(n45896), .O(n15_adj_4544));
    defparam i6_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1154 (.I0(n15_adj_4544), .I1(n45712), .I2(n14_adj_4545), 
            .I3(\data_out_frame[13] [6]), .O(n42875));
    defparam i8_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1155 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n29020));
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(\data_out_frame[16] [6]), .I1(n29020), 
            .I2(n29380), .I3(n42898), .O(n45856));
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n46058));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1158 (.I0(n45856), .I1(n42894), .I2(\data_out_frame[21][0] ), 
            .I3(GND_net), .O(n8_adj_4546));
    defparam i3_3_lut_adj_1158.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1159 (.I0(\data_out_frame[25] [4]), .I1(n45964), 
            .I2(n8_adj_4546), .I3(\data_out_frame[23] [2]), .O(n45983));
    defparam i1_4_lut_adj_1159.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1160 (.I0(n45983), .I1(\data_out_frame[25] [5]), 
            .I2(n46058), .I3(n46231), .O(n48076));
    defparam i3_4_lut_adj_1160.LUT_INIT = 16'h9669;
    SB_LUT4 mux_2021_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17] [6]), .O(n7018));
    defparam mux_2021_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2021_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n7019));
    defparam mux_2021_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_2021_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n62), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n6996));
    defparam mux_2021_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_43_26_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n40513), .O(n2_adj_4547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n40513), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n40514));
    SB_LUT4 add_43_25_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n40512), .O(n2_adj_4548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1161 (.I0(\FRAME_MATCHER.state_c [21]), .I1(\FRAME_MATCHER.state_c [25]), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(\FRAME_MATCHER.state_c [28]), 
            .O(n20_adj_4549));   // verilog/coms.v(127[12] 300[6])
    defparam i8_4_lut_adj_1161.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1162 (.I0(\FRAME_MATCHER.state_c [19]), .I1(\FRAME_MATCHER.state_c [7]), 
            .I2(\FRAME_MATCHER.state_c [6]), .I3(\FRAME_MATCHER.state_c [29]), 
            .O(n19_adj_4550));   // verilog/coms.v(127[12] 300[6])
    defparam i7_4_lut_adj_1162.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1163 (.I0(\FRAME_MATCHER.state_c [12]), .I1(\FRAME_MATCHER.state_c [11]), 
            .I2(\FRAME_MATCHER.state_c [30]), .I3(\FRAME_MATCHER.state_c [5]), 
            .O(n21_adj_4551));   // verilog/coms.v(127[12] 300[6])
    defparam i9_4_lut_adj_1163.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut_adj_1164 (.I0(n21_adj_4551), .I1(n19_adj_4550), .I2(n20_adj_4549), 
            .I3(GND_net), .O(n45486));   // verilog/coms.v(127[12] 300[6])
    defparam i11_3_lut_adj_1164.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1165 (.I0(\FRAME_MATCHER.state_c [16]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(\FRAME_MATCHER.state_c [18]), 
            .O(n160));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1165.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1166 (.I0(\FRAME_MATCHER.state_c [9]), .I1(\FRAME_MATCHER.state_c [10]), 
            .I2(\FRAME_MATCHER.state_c [14]), .I3(\FRAME_MATCHER.state_c [13]), 
            .O(n45614));
    defparam i3_4_lut_adj_1166.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_25 (.CI(n40512), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n40513));
    SB_LUT4 add_43_24_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n40511), .O(n2_adj_4552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n40511), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n40512));
    SB_LUT4 add_43_23_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n40510), .O(n2_adj_4553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_adj_1167 (.I0(\FRAME_MATCHER.state_c [26]), .I1(\FRAME_MATCHER.state_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4554));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_adj_1167.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1168 (.I0(\FRAME_MATCHER.state_c [27]), .I1(\FRAME_MATCHER.state_c [17]), 
            .I2(n6_adj_4554), .I3(\FRAME_MATCHER.state_c [8]), .O(n7_adj_4555));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1168.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state_c [15]), 
            .I2(GND_net), .I3(GND_net), .O(n45670));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1170 (.I0(n41_adj_4511), .I1(n46_c), .I2(n42_adj_4510), 
            .I3(\data_in_frame[6] [0]), .O(n45991));
    defparam i1_2_lut_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(CLK_c), 
            .D(n7_adj_4556), .S(n44942));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1171 (.I0(n160), .I1(n45614), .I2(GND_net), .I3(GND_net), 
            .O(n43664));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1172 (.I0(n7_adj_4555), .I1(\FRAME_MATCHER.state_c [23]), 
            .I2(n45486), .I3(n45670), .O(n43663));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1172.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1173 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_4557));
    defparam i1_4_lut_adj_1173.LUT_INIT = 16'ha8a0;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n51760), .I2(n51114), .I3(byte_transmit_counter[4]), .O(n52960));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n52960_bdd_4_lut (.I0(n52960), .I1(n52819), .I2(n7_adj_4558), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n52960_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n52954));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n52954_bdd_4_lut (.I0(n52954), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n52957));
    defparam n52954_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(CLK_c), 
            .D(n45102), .S(n44946));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(CLK_c), 
            .D(n45040), .S(n42278));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(CLK_c), 
            .D(n45098), .S(n44910));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(CLK_c), 
            .D(n45094), .S(n44948));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(CLK_c), 
            .D(n7_adj_4559), .S(n35660));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(CLK_c), 
            .D(n7_adj_4560), .S(n8_adj_4561));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(CLK_c), 
            .D(n45090), .S(n44950));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(CLK_c), 
            .D(n35658), .S(n36461));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(CLK_c), 
            .D(n45086), .S(n44952));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(CLK_c), 
            .D(n7_adj_4562), .S(n8_adj_4563));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(CLK_c), 
            .D(n45082), .S(n44954));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(CLK_c), 
            .D(n7_adj_4564), .S(n8_adj_4565));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(CLK_c), 
            .D(n7_adj_4566), .S(n8_adj_4567));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(CLK_c), 
            .D(n45078), .S(n42276));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(CLK_c), 
            .D(n35656), .S(n8_adj_4568));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(CLK_c), 
            .D(n45012), .S(n44884));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(CLK_c), 
            .D(n45074), .S(n44956));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(CLK_c), 
            .D(n45010), .S(n44902));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(CLK_c), 
            .D(n35650), .S(n8_adj_4569));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_23 (.CI(n40510), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n40511));
    SB_LUT4 i2_2_lut_adj_1174 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4570));
    defparam i2_2_lut_adj_1174.LUT_INIT = 16'heeee;
    SB_LUT4 i36480_4_lut (.I0(byte_transmit_counter[3]), .I1(n6_adj_4570), 
            .I2(byte_transmit_counter[7]), .I3(n4_adj_4557), .O(tx_transmit_N_3513));
    defparam i36480_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i36485_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n35937));
    defparam i36485_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(\FRAME_MATCHER.state [0]), .I1(n32424), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n35937), .O(n7099));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'hecfc;
    SB_LUT4 mux_1377_i1_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n51044), 
            .I2(n36547), .I3(n58), .O(n4882[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_1377_i1_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i5_4_lut_adj_1176 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n7_adj_4555), 
            .I2(n45614), .I3(n8_adj_4571), .O(n45491));   // verilog/coms.v(127[12] 300[6])
    defparam i5_4_lut_adj_1176.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1177 (.I0(n41_adj_4511), .I1(n46_c), .I2(n42_adj_4510), 
            .I3(n46077), .O(n6_adj_4519));
    defparam i1_2_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n10_adj_4495));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(CLK_c), 
            .D(n45070), .S(n44958));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37277 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27][1] ), 
            .I3(byte_transmit_counter[1]), .O(n52948));
    defparam byte_transmit_counter_0__bdd_4_lut_37277.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(CLK_c), 
            .D(n45066), .S(n44960));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(CLK_c), 
            .D(n45062), .S(n44962));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(CLK_c), 
            .D(n45058), .S(n44964));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(CLK_c), 
            .D(n45054), .S(n44966));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(CLK_c), 
            .D(n45006), .S(n44968));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(CLK_c), 
            .D(n45050), .S(n44892));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(CLK_c), 
            .D(n44896), .S(n10_adj_4572));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state_c [1]), .C(CLK_c), 
            .D(n44890), .S(n52972));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n52948_bdd_4_lut (.I0(n52948), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n52951));
    defparam n52948_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n29783), .D(n45745));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_22_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n40509), .O(n2_adj_4573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1178 (.I0(n35635), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n45616));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1178.LUT_INIT = 16'hffdf;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n29783), .D(n48076));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n29783), .D(n48173));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n29783), .D(n47315));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n29783), .D(n46908));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n29783), .D(n45882));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n29783), .D(n43834));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n29783), .D(n47644));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n29783), .D(n48289));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n29783), .D(n46928));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n29783), .D(n47769));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n29783), .D(n48100));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n29783), .D(n47422));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n29783), .D(n47566));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n29783), .D(n47661));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37272 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n52942));
    defparam byte_transmit_counter_0__bdd_4_lut_37272.LUT_INIT = 16'he4aa;
    SB_LUT4 n52942_bdd_4_lut (.I0(n52942), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n52945));
    defparam n52942_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1179 (.I0(n1519), .I1(n28528), .I2(\data_out_frame[14] [6]), 
            .I3(n1516), .O(n46148));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[19] [6]), .I1(n45777), .I2(\data_out_frame[22] [0]), 
            .I3(GND_net), .O(n46222));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45635));   // verilog/coms.v(231[5:23])
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1181 (.I0(\data_out_frame[7] [1]), .I1(n1168), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n46145));
    defparam i1_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n45703));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1183 (.I0(n29293), .I1(n46253), .I2(n46145), 
            .I3(n45837), .O(n28127));
    defparam i3_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1184 (.I0(n28127), .I1(n45703), .I2(n46086), 
            .I3(n46237), .O(n43910));
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37267 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n52936));
    defparam byte_transmit_counter_0__bdd_4_lut_37267.LUT_INIT = 16'he4aa;
    SB_LUT4 n52936_bdd_4_lut (.I0(n52936), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n52939));
    defparam n52936_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37262 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n52924));
    defparam byte_transmit_counter_0__bdd_4_lut_37262.LUT_INIT = 16'he4aa;
    SB_LUT4 n52924_bdd_4_lut (.I0(n52924), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n52927));
    defparam n52924_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37252 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n52918));
    defparam byte_transmit_counter_0__bdd_4_lut_37252.LUT_INIT = 16'he4aa;
    SB_LUT4 n52918_bdd_4_lut (.I0(n52918), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n52921));
    defparam n52918_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37247 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n52912));
    defparam byte_transmit_counter_0__bdd_4_lut_37247.LUT_INIT = 16'he4aa;
    SB_LUT4 n52912_bdd_4_lut (.I0(n52912), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n52915));
    defparam n52912_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37242 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n52906));
    defparam byte_transmit_counter_0__bdd_4_lut_37242.LUT_INIT = 16'he4aa;
    SB_LUT4 n52906_bdd_4_lut (.I0(n52906), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n52909));
    defparam n52906_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37237 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n52900));
    defparam byte_transmit_counter_0__bdd_4_lut_37237.LUT_INIT = 16'he4aa;
    SB_LUT4 n52900_bdd_4_lut (.I0(n52900), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n52903));
    defparam n52900_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28528));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1186 (.I0(n46246), .I1(\data_out_frame[12] [1]), 
            .I2(n43979), .I3(\data_out_frame[11] [2]), .O(n16_adj_4574));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_1186.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1187 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[11] [4]), 
            .O(n17_adj_4575));   // verilog/coms.v(85[17:63])
    defparam i7_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1188 (.I0(n17_adj_4575), .I1(n45685), .I2(n16_adj_4574), 
            .I3(n28528), .O(n46086));   // verilog/coms.v(85[17:63])
    defparam i9_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4455), .S(n3_adj_4576));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4460), .S(n3_adj_4577));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4466), .S(n3_adj_4578));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4469), .S(n3_adj_4579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4483), .S(n3_adj_4580));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4486), .S(n3_adj_4581));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4506), .S(n3_adj_4582));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4547), .S(n3_adj_4583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4548), .S(n3_adj_4584));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4552), .S(n3_adj_4585));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4553), .S(n3_adj_4586));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4573), .S(n3_adj_4587));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4588), .S(n3_adj_4589));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4590), .S(n3_adj_4591));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4592), .S(n3_adj_4593));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4594), .S(n3_adj_4595));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4596), .S(n3_adj_4597));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4598), .S(n3_adj_4599));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4600), .S(n3_adj_4601));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4602), .S(n3_adj_4603));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4604), .S(n3_adj_4605));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1189 (.I0(n29034), .I1(\data_out_frame[5] [6]), 
            .I2(n46086), .I3(\data_out_frame[5] [5]), .O(n18_adj_4606));
    defparam i7_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4607), .S(n3_adj_4608));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4609), .S(n3_adj_4610));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4611), .S(n3_adj_4612));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4613), .S(n3_adj_4614));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4615), .S(n3_adj_4616));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4617), .S(n3_adj_4618));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4619), .S(n3_adj_4620));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4621), .S(n3_adj_4622));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4623), .S(n3_adj_4624));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4625), .S(n3_adj_4626));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1190 (.I0(\data_out_frame[19] [6]), .I1(n45777), 
            .I2(\data_out_frame[20][0] ), .I3(\data_out_frame[22] [2]), 
            .O(n48133));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_993));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_43_22 (.CI(n40509), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n40510));
    SB_LUT4 i5_2_lut (.I0(n45712), .I1(n29293), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4627));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1191 (.I0(\data_out_frame[11] [5]), .I1(n18_adj_4606), 
            .I2(n45737), .I3(n46263), .O(n20_adj_4628));
    defparam i9_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1192 (.I0(n46178), .I1(n20_adj_4628), .I2(n16_adj_4627), 
            .I3(n46071), .O(n28113));
    defparam i10_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_out_frame[14] [1]), .I1(n45869), 
            .I2(GND_net), .I3(GND_net), .O(n28941));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1194 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n46178));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_21_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n40508), .O(n2_adj_4588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1195 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(n45901), .I3(n6_adj_4629), .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4630));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1197 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[4] [2]), .I3(n6_adj_4630), .O(n45784));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1198 (.I0(\data_out_frame[5] [6]), .I1(n45784), 
            .I2(\data_out_frame[6] [3]), .I3(\data_out_frame[6] [2]), .O(n12_adj_4631));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1199 (.I0(\data_out_frame[6] [1]), .I1(n12_adj_4631), 
            .I2(n1519), .I3(\data_out_frame[10] [4]), .O(n45824));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29502));
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_out_frame[14] [7]), .I1(n45824), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4496));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1202 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[16] [7]), 
            .I2(n45752), .I3(n6_adj_4632), .O(n47800));
    defparam i4_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1203 (.I0(n45846), .I1(\data_out_frame[19] [1]), 
            .I2(\data_out_frame[21][3] ), .I3(n46151), .O(n10_adj_4633));
    defparam i4_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1204 (.I0(n47800), .I1(n10_adj_4633), .I2(\data_out_frame[19] [2]), 
            .I3(GND_net), .O(n43816));
    defparam i5_3_lut_adj_1204.LUT_INIT = 16'h6969;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(85[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[19] [2]), .I1(n45976), 
            .I2(GND_net), .I3(GND_net), .O(n46213));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1206 (.I0(n28510), .I1(n46169), .I2(\data_out_frame[6] [0]), 
            .I3(n1247), .O(n12_adj_4634));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(n1668), .I1(n12_adj_4634), .I2(n46074), 
            .I3(\data_out_frame[13] [0]), .O(n42909));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28519));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46017));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1210 (.I0(\data_out_frame[17] [2]), .I1(n46017), 
            .I2(\data_out_frame[21][4] ), .I3(n28519), .O(n12_adj_4635));
    defparam i5_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_CARRY add_43_21 (.CI(n40508), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n40509));
    SB_LUT4 i4_4_lut_adj_1211 (.I0(Kp_23__N_993), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [1]), .I3(n6_adj_4636), .O(Kp_23__N_988));   // verilog/coms.v(73[16:34])
    defparam i4_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_20_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n40507), .O(n2_adj_4590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n40507), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n40508));
    SB_LUT4 i6_4_lut_adj_1212 (.I0(n42909), .I1(n12_adj_4635), .I2(n46213), 
            .I3(\data_out_frame[19] [3]), .O(n47627));
    defparam i6_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_19_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n40506), .O(n2_adj_4592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1213 (.I0(n43121), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[21][1] ), .I3(n6_adj_4637), .O(n46231));
    defparam i4_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[9] [4]), .I1(n45770), 
            .I2(GND_net), .I3(GND_net), .O(n46119));
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1215 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(n46172), .I3(n29044), .O(n10_adj_4638));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1216 (.I0(\data_out_frame[10] [0]), .I1(n10_adj_4638), 
            .I2(\data_out_frame[10] [1]), .I3(GND_net), .O(n45709));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_adj_1216.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1217 (.I0(\data_in_frame[7] [2]), .I1(n27216), 
            .I2(n45872), .I3(n6_adj_4639), .O(n29226));
    defparam i4_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1218 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n45893));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n46169));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1220 (.I0(\data_out_frame[10] [5]), .I1(n46169), 
            .I2(n45893), .I3(\data_out_frame[10] [1]), .O(n1537));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_CARRY add_43_19 (.CI(n40506), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n40507));
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_out_frame[9] [1]), .I1(n45685), 
            .I2(GND_net), .I3(GND_net), .O(n46157));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1222 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n46234));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1223 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n45678));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45761));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1225 (.I0(\data_out_frame[5] [4]), .I1(n45925), 
            .I2(n28500), .I3(n1191), .O(n1168));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_18_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n40505), .O(n2_adj_4594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37232 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n52876));
    defparam byte_transmit_counter_0__bdd_4_lut_37232.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1226 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n28997));
    defparam i2_3_lut_adj_1226.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1227 (.I0(n28997), .I1(n4_adj_4543), .I2(GND_net), 
            .I3(GND_net), .O(n46175));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_adj_1227.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n45901));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1229 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45729));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1229.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n45837));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28500));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n45790));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(n45790), .I1(n45896), .I2(n29293), 
            .I3(GND_net), .O(n28719));
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1234 (.I0(n45901), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(\data_out_frame[4] [5]), .O(n18_adj_4640));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_CARRY add_43_18 (.CI(n40505), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n40506));
    SB_LUT4 add_43_17_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n40504), .O(n2_adj_4596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i9_4_lut_adj_1235 (.I0(\data_out_frame[4] [7]), .I1(n18_adj_4640), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[7] [1]), .O(n20_adj_4641));   // verilog/coms.v(75[16:43])
    defparam i9_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_CARRY add_43_17 (.CI(n40504), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n40505));
    SB_LUT4 i10_4_lut_adj_1236 (.I0(n46175), .I1(n20_adj_4641), .I2(n16_adj_4642), 
            .I3(\data_out_frame[4] [0]), .O(n47801));   // verilog/coms.v(75[16:43])
    defparam i10_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1237 (.I0(n46074), .I1(n29458), .I2(n45761), 
            .I3(n18_adj_4643), .O(n30_adj_4644));   // verilog/coms.v(72[16:27])
    defparam i13_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1238 (.I0(n45790), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [4]), .I3(n29044), .O(n28_adj_4645));   // verilog/coms.v(72[16:27])
    defparam i11_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_16_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n40503), .O(n2_adj_4598)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12_4_lut_adj_1239 (.I0(\data_out_frame[7] [4]), .I1(n47801), 
            .I2(n45888), .I3(n46234), .O(n29_adj_4646));   // verilog/coms.v(72[16:27])
    defparam i12_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1240 (.I0(n46157), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[9] [6]), .I3(n46082), .O(n27_adj_4647));   // verilog/coms.v(72[16:27])
    defparam i10_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1241 (.I0(n27_adj_4647), .I1(n29_adj_4646), .I2(n28_adj_4645), 
            .I3(n30_adj_4644), .O(n43887));   // verilog/coms.v(72[16:27])
    defparam i16_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(n43887), .I1(n1537), .I2(GND_net), 
            .I3(GND_net), .O(n43979));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(n43887), .I1(n28719), .I2(GND_net), 
            .I3(GND_net), .O(n43805));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n45925));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_CARRY add_43_16 (.CI(n40503), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n40504));
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(71[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1245 (.I0(n46082), .I1(n1537), .I2(\data_out_frame[7] [6]), 
            .I3(\data_out_frame[11] [7]), .O(n14_adj_4648));
    defparam i6_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1246 (.I0(\data_out_frame[10] [0]), .I1(n45925), 
            .I2(n43805), .I3(n43979), .O(n13_adj_4649));
    defparam i5_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1247 (.I0(\data_out_frame[12] [1]), .I1(n13_adj_4649), 
            .I2(n14_adj_4648), .I3(GND_net), .O(n9_adj_4650));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n45896));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_15_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n40502), .O(n2_adj_4600)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n46025));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_CARRY add_43_15 (.CI(n40502), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n40503));
    SB_LUT4 add_43_14_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n40501), .O(n2_adj_4602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n40501), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n40502));
    SB_LUT4 n52876_bdd_4_lut (.I0(n52876), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n52879));
    defparam n52876_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1250 (.I0(n9_adj_4650), .I1(n46237), .I2(\data_out_frame[5] [4]), 
            .I3(GND_net), .O(n12_adj_4651));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1251 (.I0(n45743), .I1(n12_adj_4651), .I2(\data_out_frame[14] [2]), 
            .I3(n46172), .O(n45869));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_out_frame[14] [3]), .I1(n45970), 
            .I2(GND_net), .I3(GND_net), .O(n43025));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n46082));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n45699));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28542));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1256 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n45737));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_13_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n40500), .O(n2_adj_4604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46104));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[13] [3]), .I1(n28861), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4652));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1259 (.I0(n29044), .I1(n46104), .I2(n45737), 
            .I3(n28542), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1260 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4653));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37282 (.I0(byte_transmit_counter[3]), 
            .I1(n52753), .I2(n51116), .I3(byte_transmit_counter[4]), .O(n52870));
    defparam byte_transmit_counter_3__bdd_4_lut_37282.LUT_INIT = 16'he4aa;
    SB_LUT4 n52870_bdd_4_lut (.I0(n52870), .I1(n52807), .I2(n7_adj_4654), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n52870_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37208 (.I0(byte_transmit_counter[3]), 
            .I1(n52759), .I2(n51117), .I3(byte_transmit_counter[4]), .O(n52864));
    defparam byte_transmit_counter_3__bdd_4_lut_37208.LUT_INIT = 16'he4aa;
    SB_LUT4 n52864_bdd_4_lut (.I0(n52864), .I1(n52861), .I2(n7_adj_4655), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n52864_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n50163), .I2(n50164), .I3(byte_transmit_counter[2]), .O(n52858));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n52858_bdd_4_lut (.I0(n52858), .I1(n50272), .I2(n50271), .I3(byte_transmit_counter[2]), 
            .O(n52861));
    defparam n52858_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37198 (.I0(byte_transmit_counter[1]), 
            .I1(n50196), .I2(n50197), .I3(byte_transmit_counter[2]), .O(n52852));
    defparam byte_transmit_counter_1__bdd_4_lut_37198.LUT_INIT = 16'he4aa;
    SB_LUT4 n52852_bdd_4_lut (.I0(n52852), .I1(n50251), .I2(n50250), .I3(byte_transmit_counter[2]), 
            .O(n14_adj_4656));
    defparam n52852_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37193 (.I0(byte_transmit_counter[1]), 
            .I1(n50226), .I2(n50227), .I3(byte_transmit_counter[2]), .O(n52846));
    defparam byte_transmit_counter_1__bdd_4_lut_37193.LUT_INIT = 16'he4aa;
    SB_LUT4 n52846_bdd_4_lut (.I0(n52846), .I1(n50245), .I2(n50244), .I3(byte_transmit_counter[2]), 
            .O(n14_adj_4657));
    defparam n52846_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37188 (.I0(byte_transmit_counter[1]), 
            .I1(n50262), .I2(n50263), .I3(byte_transmit_counter[2]), .O(n52840));
    defparam byte_transmit_counter_1__bdd_4_lut_37188.LUT_INIT = 16'he4aa;
    SB_LUT4 n52840_bdd_4_lut (.I0(n52840), .I1(n50236), .I2(n50235), .I3(byte_transmit_counter[2]), 
            .O(n52843));
    defparam n52840_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37183 (.I0(byte_transmit_counter[1]), 
            .I1(n50274), .I2(n50275), .I3(byte_transmit_counter[2]), .O(n52834));
    defparam byte_transmit_counter_1__bdd_4_lut_37183.LUT_INIT = 16'he4aa;
    SB_LUT4 n52834_bdd_4_lut (.I0(n52834), .I1(n50290), .I2(n50289), .I3(byte_transmit_counter[2]), 
            .O(n52837));
    defparam n52834_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1261 (.I0(\data_out_frame[10] [1]), .I1(n28542), 
            .I2(n45699), .I3(\data_out_frame[8] [1]), .O(n14_adj_4658));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1262 (.I0(\data_out_frame[12] [3]), .I1(n14_adj_4658), 
            .I2(n10_adj_4653), .I3(n46082), .O(n45814));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1263 (.I0(\data_out_frame[14] [5]), .I1(n45814), 
            .I2(\data_out_frame[12] [4]), .I3(n1516), .O(n29091));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[16] [4]), .I1(n43854), 
            .I2(GND_net), .I3(GND_net), .O(n43940));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1265 (.I0(\data_in_frame[11] [1]), .I1(n4_adj_4652), 
            .I2(n8_adj_4659), .I3(n46011), .O(n48270));
    defparam i2_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1266 (.I0(n45976), .I1(n46276), .I2(n43940), 
            .I3(GND_net), .O(n47669));
    defparam i2_3_lut_adj_1266.LUT_INIT = 16'h6969;
    SB_LUT4 i22206_2_lut_3_lut (.I0(n63_adj_4412), .I1(n63_adj_4415), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n1[1]));   // verilog/coms.v(157[6] 159[9])
    defparam i22206_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[21][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n45755));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1268 (.I0(n43025), .I1(n46148), .I2(n46017), 
            .I3(n29380), .O(n47182));
    defparam i3_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1269 (.I0(\data_out_frame[19] [1]), .I1(n45755), 
            .I2(n47182), .I3(n47669), .O(n28578));
    defparam i3_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_CARRY add_43_13 (.CI(n40500), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n40501));
    SB_LUT4 add_43_12_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n40499), .O(n2_adj_4607)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(n29195), .I1(n46030), .I2(n29261), 
            .I3(n48270), .O(n43862));
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1271 (.I0(n63_adj_4412), .I1(n63_adj_4415), 
            .I2(n63_adj_3), .I3(GND_net), .O(n25438));   // verilog/coms.v(157[6] 159[9])
    defparam i2_2_lut_3_lut_adj_1271.LUT_INIT = 16'h8080;
    SB_LUT4 i21984_2_lut_3_lut_4_lut (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(n45642), .O(n35660));
    defparam i21984_2_lut_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(\data_out_frame[23] [3]), .I1(n28578), 
            .I2(GND_net), .I3(GND_net), .O(n45964));
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1273 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[23] [5]), 
            .I2(\data_out_frame[25] [6]), .I3(n45964), .O(n10_adj_4660));
    defparam i4_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1274 (.I0(n46231), .I1(n10_adj_4660), .I2(n47627), 
            .I3(GND_net), .O(n45745));
    defparam i5_3_lut_adj_1274.LUT_INIT = 16'h6969;
    SB_LUT4 i26716_2_lut_3_lut_4_lut (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [28]), 
            .I3(n45642), .O(n42278));
    defparam i26716_2_lut_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_3_lut_4_lut (.I0(n25438), .I1(n3807), .I2(n3_adj_4661), 
            .I3(\FRAME_MATCHER.state[3] ), .O(n44896));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i7_4_lut_adj_1275 (.I0(n46163), .I1(n45817), .I2(\data_in_frame[15] [6]), 
            .I3(\data_in_frame[16] [0]), .O(n18_adj_4662));   // verilog/coms.v(70[16:27])
    defparam i7_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n25438), .I1(n3807), .I2(n771), 
            .I3(n42259), .O(n45651));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i1_2_lut_4_lut_adj_1276 (.I0(\data_in_frame[1] [2]), .I1(n10_adj_4433), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[5] [5]), .O(n45910));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [22]), 
            .I3(n45642), .O(n36461));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_4_lut_4_lut (.I0(n25438), .I1(n3807), .I2(n38), .I3(n46495), 
            .O(n11_adj_4663));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1277 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [20]), 
            .I3(n45642), .O(n8_adj_4563));
    defparam i1_2_lut_3_lut_4_lut_adj_1277.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1278 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [18]), 
            .I3(n45642), .O(n8_adj_4565));
    defparam i1_2_lut_3_lut_4_lut_adj_1278.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1279 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [17]), 
            .I3(n45642), .O(n8_adj_4567));
    defparam i1_2_lut_3_lut_4_lut_adj_1279.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_4_lut_adj_1280 (.I0(\data_in_frame[1] [2]), .I1(n10_adj_4433), 
            .I2(\data_in_frame[3] [3]), .I3(n45875), .O(n42921));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_CARRY add_43_12 (.CI(n40499), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n40500));
    SB_LUT4 i1_2_lut_4_lut_adj_1281 (.I0(n28977), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_988), .I3(\data_in_frame[7] [5]), .O(n6_adj_4491));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1282 (.I0(n28977), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_988), .I3(n45764), .O(n6_adj_4664));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i26715_2_lut_3_lut_4_lut (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [16]), 
            .I3(n45642), .O(n42276));
    defparam i26715_2_lut_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1283 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [15]), 
            .I3(n45642), .O(n8_adj_4568));
    defparam i1_2_lut_3_lut_4_lut_adj_1283.LUT_INIT = 16'hf080;
    SB_LUT4 i5_2_lut_adj_1284 (.I0(\data_in_frame[13] [5]), .I1(n29226), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4665));   // verilog/coms.v(70[16:27])
    defparam i5_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1285 (.I0(n46025), .I1(n18_adj_4662), .I2(\data_in_frame[18] [2]), 
            .I3(n29105), .O(n20_adj_4666));   // verilog/coms.v(70[16:27])
    defparam i9_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [12]), 
            .I3(n45642), .O(n44902));
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1287 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [11]), 
            .I3(n45642), .O(n8_adj_4569));
    defparam i1_2_lut_3_lut_4_lut_adj_1287.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1288 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [24]), 
            .I3(n45642), .O(n8_adj_4561));
    defparam i1_2_lut_3_lut_4_lut_adj_1288.LUT_INIT = 16'hf080;
    SB_LUT4 add_43_11_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n40498), .O(n2_adj_4609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1289 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [5]), 
            .I3(n45642), .O(n44968));
    defparam i1_2_lut_3_lut_4_lut_adj_1289.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1290 (.I0(n25438), .I1(n3807), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(n45642), .O(n44910));
    defparam i1_2_lut_3_lut_4_lut_adj_1290.LUT_INIT = 16'hf080;
    SB_LUT4 i3_3_lut_4_lut (.I0(n28750), .I1(n6_adj_4479), .I2(n46249), 
            .I3(n28977), .O(n45872));   // verilog/coms.v(74[16:43])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_43_11 (.CI(n40498), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n40499));
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37178 (.I0(byte_transmit_counter[1]), 
            .I1(n50223), .I2(n50224), .I3(byte_transmit_counter[2]), .O(n52822));
    defparam byte_transmit_counter_1__bdd_4_lut_37178.LUT_INIT = 16'he4aa;
    SB_LUT4 n52822_bdd_4_lut (.I0(n52822), .I1(n50302), .I2(n50301), .I3(byte_transmit_counter[2]), 
            .O(n52825));
    defparam n52822_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_adj_1291 (.I0(n28750), .I1(n6_adj_4479), .I2(n29137), 
            .I3(GND_net), .O(n10_adj_4475));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_adj_1291.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_10_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n40497), .O(n2_adj_4611)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n40497), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n40498));
    SB_LUT4 add_43_9_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n40496), .O(n2_adj_4613)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10_4_lut_adj_1292 (.I0(\data_in_frame[16] [1]), .I1(n20_adj_4666), 
            .I2(n16_adj_4665), .I3(\data_in_frame[13] [4]), .O(n46133));   // verilog/coms.v(70[16:27])
    defparam i10_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_CARRY add_43_9 (.CI(n40496), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n40497));
    SB_LUT4 i16754_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n30443));
    defparam i16754_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_8_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n40495), .O(n2_adj_4615)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37169 (.I0(byte_transmit_counter[1]), 
            .I1(n50298), .I2(n50299), .I3(byte_transmit_counter[2]), .O(n52816));
    defparam byte_transmit_counter_1__bdd_4_lut_37169.LUT_INIT = 16'he4aa;
    SB_LUT4 n52816_bdd_4_lut (.I0(n52816), .I1(n50221), .I2(n50220), .I3(byte_transmit_counter[2]), 
            .O(n52819));
    defparam n52816_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37164 (.I0(byte_transmit_counter[1]), 
            .I1(n50304), .I2(n50305), .I3(byte_transmit_counter[2]), .O(n52804));
    defparam byte_transmit_counter_1__bdd_4_lut_37164.LUT_INIT = 16'he4aa;
    SB_LUT4 n52804_bdd_4_lut (.I0(n52804), .I1(n50284), .I2(n50283), .I3(byte_transmit_counter[2]), 
            .O(n52807));
    defparam n52804_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37203 (.I0(byte_transmit_counter[3]), 
            .I1(n51822), .I2(n51122), .I3(byte_transmit_counter[4]), .O(n52798));
    defparam byte_transmit_counter_3__bdd_4_lut_37203.LUT_INIT = 16'he4aa;
    SB_LUT4 n52798_bdd_4_lut (.I0(n52798), .I1(n14_adj_4656), .I2(n7_adj_4668), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n52798_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37213 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[1]), .O(n52792));
    defparam byte_transmit_counter_0__bdd_4_lut_37213.LUT_INIT = 16'he4aa;
    SB_LUT4 n52792_bdd_4_lut (.I0(n52792), .I1(\data_out_frame[21][0] ), 
            .I2(\data_out_frame[20][0] ), .I3(byte_transmit_counter[1]), 
            .O(n52795));
    defparam n52792_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_8 (.CI(n40495), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n40496));
    SB_LUT4 add_43_7_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n40494), .O(n2_adj_4617)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n40494), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n40495));
    SB_LUT4 i16755_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n30444));
    defparam i16755_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_6_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n40493), .O(n2_adj_4619)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16756_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n30445));
    defparam i16756_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16757_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n30446));
    defparam i16757_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21978_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2025));
    defparam i21978_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1293 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n54), .I3(\FRAME_MATCHER.state[3] ), .O(n63));   // verilog/coms.v(201[5:24])
    defparam i3_4_lut_adj_1293.LUT_INIT = 16'hfeff;
    SB_LUT4 i16758_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n30447));
    defparam i16758_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16759_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n30448));
    defparam i16759_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1294 (.I0(n29645), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n45), .O(n39711));
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'haa2a;
    SB_LUT4 i16760_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n30449));
    defparam i16760_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16761_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n30450));
    defparam i16761_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_6 (.CI(n40493), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n40494));
    SB_LUT4 i16746_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n30435));
    defparam i16746_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16747_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n30436));
    defparam i16747_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_37150 (.I0(byte_transmit_counter[3]), 
            .I1(n52741), .I2(n51118), .I3(byte_transmit_counter[4]), .O(n52786));
    defparam byte_transmit_counter_3__bdd_4_lut_37150.LUT_INIT = 16'he4aa;
    SB_LUT4 i16748_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n30437));
    defparam i16748_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16749_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n30438));
    defparam i16749_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16750_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n30439));
    defparam i16750_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30774_2_lut (.I0(n46), .I1(n4452), .I2(GND_net), .I3(GND_net), 
            .O(n46338));
    defparam i30774_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16751_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n30440));
    defparam i16751_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_685_Select_1_i5_4_lut (.I0(n63_adj_3), .I1(n42261), .I2(n3303), 
            .I3(n1[1]), .O(n5_adj_4672));
    defparam select_685_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i16752_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n30441));
    defparam i16752_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_5_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n40492), .O(n2_adj_4621)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n40492), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n40493));
    SB_LUT4 i2_4_lut_adj_1295 (.I0(n1[1]), .I1(n5_adj_4672), .I2(n46338), 
            .I3(n63_adj_3), .O(n6_adj_4673));
    defparam i2_4_lut_adj_1295.LUT_INIT = 16'hcecf;
    SB_LUT4 i3_4_lut_adj_1296 (.I0(n63), .I1(n6_adj_4673), .I2(\FRAME_MATCHER.state_31__N_2692 [1]), 
            .I3(n42259), .O(n52972));
    defparam i3_4_lut_adj_1296.LUT_INIT = 16'hddfd;
    SB_LUT4 i16753_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n30442));
    defparam i16753_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_300_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4670));   // verilog/coms.v(154[7:23])
    defparam equal_300_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_291_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4674));   // verilog/coms.v(154[7:23])
    defparam equal_291_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i16738_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n30427));
    defparam i16738_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16739_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n30428));
    defparam i16739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1297 (.I0(\FRAME_MATCHER.state[3] ), .I1(n94), 
            .I2(n45642), .I3(GND_net), .O(n94_adj_4675));
    defparam i1_3_lut_adj_1297.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_1298 (.I0(n28494), .I1(n94_adj_4675), .I2(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .I3(n28386), .O(n10_adj_4572));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1298.LUT_INIT = 16'hccdc;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44892));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h8888;
    SB_LUT4 i16740_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n30429));
    defparam i16740_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n7_adj_4676), 
            .I2(GND_net), .I3(GND_net), .O(n44966));
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h8888;
    SB_LUT4 n52786_bdd_4_lut (.I0(n52786), .I1(n14_adj_4657), .I2(n7_adj_4677), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n52786_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n7_adj_4676), 
            .I2(GND_net), .I3(GND_net), .O(n44964));
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1302 (.I0(n38), .I1(n45651), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n25525), .O(n7_adj_4676));
    defparam i1_4_lut_adj_1302.LUT_INIT = 16'hdccc;
    SB_LUT4 i16741_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n30430));
    defparam i16741_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16742_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n30431));
    defparam i16742_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n7_adj_4676), 
            .I2(GND_net), .I3(GND_net), .O(n44962));
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h8888;
    SB_LUT4 i34510_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n50143), .I3(n20_adj_4432), .O(n50144));
    defparam i34510_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 add_43_4_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n40491), .O(n2_adj_4623)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n40491), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n40492));
    SB_LUT4 i34513_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n50146), .I3(n20_adj_4438), .O(n50147));
    defparam i34513_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i16743_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n30432));
    defparam i16743_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44958));
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h8888;
    SB_LUT4 i77_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n58));   // verilog/coms.v(112[11:16])
    defparam i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1305 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28389));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'hbbbb;
    SB_LUT4 i16744_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n30433));
    defparam i16744_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16745_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n30434));
    defparam i16745_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34516_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n50149), .I3(n20_adj_4447), .O(n50150));
    defparam i34516_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i22055_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i22055_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50180), .I3(n50178), .O(n7_adj_4677));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50174), .I3(n50172), .O(n7_adj_4668));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i4_4_lut_adj_1306 (.I0(\data_in_frame[7] [3]), .I1(n29223), 
            .I2(\data_in_frame[5] [1]), .I3(n6_adj_4664), .O(n43430));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44956));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [4]), 
            .I3(GND_net), .O(n45050));
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50168), .I3(n50166), .O(n7_adj_4655));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1309 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [5]), 
            .I3(GND_net), .O(n45006));
    defparam i1_2_lut_3_lut_adj_1309.LUT_INIT = 16'he0e0;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
           .D(n44944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n30166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n30165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n30164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n30163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n30162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n30161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n30160));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1310 (.I0(\FRAME_MATCHER.state [0]), 
            .I1(\FRAME_MATCHER.state_c [1]), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n67), .O(n4_c));
    defparam i1_2_lut_3_lut_4_lut_adj_1310.LUT_INIT = 16'h5554;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44884));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h8888;
    SB_LUT4 i36477_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n67), .O(n36742));
    defparam i36477_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1312 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [6]), 
            .I3(GND_net), .O(n45054));
    defparam i1_2_lut_3_lut_adj_1312.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [7]), 
            .I3(GND_net), .O(n45058));
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_3_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n40490), .O(n2_adj_4625)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1314 (.I0(n45491), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(\FRAME_MATCHER.state_c [15]), .I3(n45635), .O(n28494));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1314.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1315 (.I0(n45491), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(\FRAME_MATCHER.state_c [15]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n54));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1315.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1316 (.I0(\data_in_frame[18] [7]), .I1(n45999), 
            .I2(\data_in_frame[18] [6]), .I3(\data_in_frame[16] [4]), .O(n45996));
    defparam i3_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1317 (.I0(n43811), .I1(n46279), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4679));
    defparam i4_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1318 (.I0(n54), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n28426));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1318.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1319 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [8]), 
            .I3(GND_net), .O(n45062));
    defparam i1_2_lut_3_lut_adj_1319.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50159), .I3(n50157), .O(n7_adj_4654));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1320 (.I0(\data_out_frame[14] [1]), .I1(n45869), 
            .I2(n28113), .I3(\data_out_frame[16] [3]), .O(n28910));
    defparam i1_2_lut_3_lut_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1321 (.I0(n46139), .I1(\data_in_frame[9] [7]), 
            .I2(n45916), .I3(\data_in_frame[9] [6]), .O(n24_adj_4680));
    defparam i10_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1322 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[11] [6]), 
            .I2(n43836), .I3(n29505), .O(n22));
    defparam i8_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1323 (.I0(n46228), .I1(n24_adj_4680), .I2(n18_adj_4679), 
            .I3(n28981), .O(n26_adj_4681));
    defparam i12_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1324 (.I0(n42892), .I1(n26_adj_4681), .I2(n22), 
            .I3(n43430), .O(n45750));
    defparam i13_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1325 (.I0(n43899), .I1(n45930), .I2(n43915), 
            .I3(GND_net), .O(n27975));
    defparam i2_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1326 (.I0(n43606), .I1(n43899), .I2(n46203), 
            .I3(GND_net), .O(n8_adj_4682));
    defparam i3_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1327 (.I0(\data_in_frame[19] [0]), .I1(n45750), 
            .I2(n8_adj_4682), .I3(n45996), .O(n45904));
    defparam i1_4_lut_adj_1327.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1328 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4683));
    defparam i2_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 i21963_2_lut_2_lut_3_lut (.I0(n36474), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n35635));
    defparam i21963_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [9]), 
            .I3(GND_net), .O(n45066));
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1330 (.I0(\data_out_frame[14] [1]), .I1(n45869), 
            .I2(n28113), .I3(\data_out_frame[17] [7]), .O(n46206));
    defparam i1_2_lut_3_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [10]), 
            .I3(GND_net), .O(n45070));
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1332 (.I0(\data_out_frame[16] [4]), .I1(n43854), 
            .I2(n46151), .I3(n46276), .O(n42898));
    defparam i1_2_lut_3_lut_4_lut_adj_1332.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1333 (.I0(n46042), .I1(n43800), .I2(n29261), 
            .I3(\data_in_frame[17] [7]), .O(n14_adj_4684));
    defparam i6_4_lut_adj_1333.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1334 (.I0(\data_in_frame[15] [6]), .I1(n14_adj_4684), 
            .I2(n10_adj_4683), .I3(n43862), .O(n43222));
    defparam i7_4_lut_adj_1334.LUT_INIT = 16'h9669;
    SB_LUT4 i1_rep_74_2_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[19] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n53051));
    defparam i1_rep_74_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1335 (.I0(\data_in_frame[18] [5]), .I1(n10_adj_4436), 
            .I2(\data_in_frame[19] [0]), .I3(GND_net), .O(n12_adj_4685));
    defparam i5_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1336 (.I0(n43797), .I1(\data_in_frame[20] [0]), 
            .I2(n43222), .I3(n53051), .O(n10_adj_4686));
    defparam i4_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1337 (.I0(n43876), .I1(n12_adj_4685), .I2(n46219), 
            .I3(\data_in_frame[20] [7]), .O(n47755));
    defparam i6_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(n29255), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4687));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1339 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n6_adj_4688));
    defparam i2_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1340 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [2]), .I3(GND_net), .O(n7_adj_4689));
    defparam i2_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1341 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[6] [3]), .O(n1247));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i21977_2_lut_3_lut (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [11]), 
            .I3(GND_net), .O(n35650));
    defparam i21977_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [12]), 
            .I3(GND_net), .O(n45010));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44954));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1344 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[5] [2]), .O(n46172));
    defparam i1_2_lut_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [13]), 
            .I3(GND_net), .O(n45074));
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1346 (.I0(n45491), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n45670), .O(n45));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1346.LUT_INIT = 16'hffef;
    SB_LUT4 i3_4_lut_adj_1347 (.I0(\data_in_frame[20] [6]), .I1(n45913), 
            .I2(n43876), .I3(Kp_23__N_1803), .O(n47169));
    defparam i3_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50156), .I3(n50154), .O(n7_adj_4558));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n30742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n30741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n30740));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n30739));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n30738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n30737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n30736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n30735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n30734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n30733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n30732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n30731));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44952));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50189), .I3(n50187), .O(n7));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(tx_transmit_N_3513), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3616[0]), .I3(n28383), .O(n7_adj_4690));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'h00fe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1350 (.I0(n28750), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(\data_in_frame[0] [2]), .O(Kp_23__N_1020));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i22333_2_lut_3_lut_4_lut (.I0(n63_adj_3), .I1(n42507), .I2(\FRAME_MATCHER.i [31]), 
            .I3(n1[1]), .O(\FRAME_MATCHER.state_31__N_2692 [1]));   // verilog/coms.v(157[6] 159[9])
    defparam i22333_2_lut_3_lut_4_lut.LUT_INIT = 16'hff5d;
    SB_LUT4 equal_2181_i19_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4190));
    defparam equal_2181_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44950));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1352 (.I0(\data_out_frame[11] [5]), .I1(n29293), 
            .I2(\data_out_frame[9] [4]), .I3(n45770), .O(n46039));
    defparam i1_2_lut_3_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i85_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n43663), 
            .I2(n160), .I3(n45614), .O(n67));
    defparam i85_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1353 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[6] [3]), .O(n46071));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(n28276), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25438), .I3(GND_net), .O(n25525));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44948));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1356 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n45936), .I3(\data_in_frame[10] [0]), .O(n42892));
    defparam i1_2_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(n25525), .I1(n42261), .I2(GND_net), 
            .I3(GND_net), .O(n117));
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_adj_1358 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n25525), 
            .I2(n42261), .I3(n45651), .O(n44960));
    defparam i1_3_lut_4_lut_adj_1358.LUT_INIT = 16'haa08;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [14]), 
            .I3(GND_net), .O(n45012));
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1360 (.I0(Kp_23__N_1195), .I1(\data_in_frame[8] [6]), 
            .I2(n8_adj_4429), .I3(n46269), .O(n29105));
    defparam i1_2_lut_3_lut_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i21982_2_lut_3_lut (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [15]), 
            .I3(GND_net), .O(n35656));
    defparam i21982_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(Kp_23__N_1195), .I1(\data_in_frame[8] [6]), 
            .I2(n8_adj_4429), .I3(n28892), .O(n10_adj_4457));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1361 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44946));
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50204), .I3(n50202), .O(n7_adj_4448));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [16]), 
            .I3(GND_net), .O(n45078));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n7227));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [17]), 
            .I3(GND_net), .O(n7_adj_4566));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n50195), .I3(n50193), .O(n7_adj_4440));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i34521_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50155));
    defparam i34521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34522_4_lut (.I0(n50155), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n50156));
    defparam i34522_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i34520_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n50154));
    defparam i34520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35594_2_lut (.I0(n52957), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n51114));
    defparam i35594_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i36125_3_lut (.I0(n52879), .I1(n52795), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n51760));
    defparam i36125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36599_3_lut_4_lut (.I0(n63), .I1(tx_active), .I2(r_SM_Main_2__N_3616[0]), 
            .I3(n28383), .O(n29645));
    defparam i36599_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 equal_285_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4667));   // verilog/coms.v(154[7:23])
    defparam equal_285_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(n46139), .I1(n46249), .I2(n28827), 
            .I3(GND_net), .O(n45936));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [18]), 
            .I3(GND_net), .O(n7_adj_4564));
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'he0e0;
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n30730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n30729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n30728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n30727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n30726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n30725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n30724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n30723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n30722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n30721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n30719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n30718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n30717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n30716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n30715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n30714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n30713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n30712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n30711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n30710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n30709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n30708));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_3 (.CI(n40490), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n40491));
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44942));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [19]), 
            .I3(GND_net), .O(n45082));
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1369 (.I0(n43017), .I1(n43862), .I2(n46219), 
            .I3(GND_net), .O(n6_adj_4691));
    defparam i2_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_2_lut (.I0(n3059), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [20]), 
            .I3(GND_net), .O(n7_adj_4562));
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n40490));
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n30707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n30706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n30705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n30704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n30703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n30702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n30701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n30700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n30699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n30698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n30697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n30696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n30695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n30694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n30693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n30692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n30691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n30690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n30689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n30688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n30687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n30686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n30685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n30684));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n30683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n30682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n30681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n30680));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n30679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n30678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n30677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n30676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n30675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n30674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n30673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n30671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n30670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n30669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n30668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n30667));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n30666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n30665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n30664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n30663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n30662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n30661));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n30660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n30659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n30658));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n30657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n30656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n30655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n30654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n30653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n30652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n30651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n30650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n30649));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n30648));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n30647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n30646));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n30645));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n30644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n30643));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n30642));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n30641));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n30640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n30639));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n30638));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1371 (.I0(n43017), .I1(n45885), .I2(n29255), 
            .I3(\data_in_frame[21] [1]), .O(n46949));
    defparam i2_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [21]), 
            .I3(GND_net), .O(n45086));
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [22]), 
            .I3(GND_net), .O(n35658));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [23]), 
            .I3(GND_net), .O(n45090));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n30637));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n30636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n30635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n30634));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n30633));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n30632));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n30631));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n30630));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n30629));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n30628));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1375 (.I0(\data_out_frame[14] [3]), .I1(n45970), 
            .I2(n45869), .I3(GND_net), .O(n43854));
    defparam i1_2_lut_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n29044));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [24]), 
            .I3(GND_net), .O(n7_adj_4560));
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n30627));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n30626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n30625));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n30624));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n30623));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n30622));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n30621));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n30620));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n30619));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n30618));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n30617));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n30616));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n30615));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n30614));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n30613));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n30612));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n30611));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_286_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4692));   // verilog/coms.v(154[7:23])
    defparam equal_286_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n30610));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n30609));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n30608));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n30607));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n30606));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n30605));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n30604));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n30603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n30602));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n30601));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n30600));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n30599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n30598));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n30597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n30596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n30595));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n30594));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n30593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n30592));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n30591));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n30590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n30589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n30588));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n30587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n30586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n30585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n30584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n30583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n30582));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n30581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n30580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n30579));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n30578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n30577));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n30576));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n30575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n30574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n30573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n30572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n30571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n30570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n30569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n30568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n30567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n30566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n30565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n30564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n30563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n30562));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n30561));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n30560));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n30559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n30558));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n30557));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n30556));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n30555));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n30554));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n30553));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n30552));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n30551));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n30550));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n30549));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n30548));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n30547));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n30546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n30545));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n30544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n30543));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n30542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n30541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n30540));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n30539));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n30538));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n30537));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n30536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n30535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n30534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n30533));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(GND_net), .O(n7_adj_4559));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n30532));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n30531));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [26]), 
            .I3(GND_net), .O(n45094));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n30530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n30529));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(GND_net), .O(n45098));
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20][0] ), .C(CLK_c), 
           .D(n30528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20][1] ), .C(CLK_c), 
           .D(n30527));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1381 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [28]), 
            .I3(GND_net), .O(n45040));
    defparam i1_2_lut_3_lut_adj_1381.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n30526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n30525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20]_c [4]), .C(CLK_c), 
           .D(n30524));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [29]), 
            .I3(GND_net), .O(n45102));
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n30523));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(n94), .I1(n3_adj_4661), .I2(\FRAME_MATCHER.state_c [30]), 
            .I3(GND_net), .O(n7_adj_4556));
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n30522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n30521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21][0] ), .C(CLK_c), 
           .D(n30520));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_3_lut_4_lut_adj_1384 (.I0(n29105), .I1(n43836), .I2(n28776), 
            .I3(\data_in_frame[9] [1]), .O(n8_adj_4659));
    defparam i3_3_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21][1] ), .C(CLK_c), 
           .D(n30519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21][2] ), .C(CLK_c), 
           .D(n30518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21][3] ), .C(CLK_c), 
           .D(n30517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21][4] ), .C(CLK_c), 
           .D(n30516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(CLK_c), 
           .D(n30515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(CLK_c), 
           .D(n30514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(CLK_c), 
           .D(n30513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(CLK_c), 
           .D(n30512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(CLK_c), 
           .D(n30511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(CLK_c), 
           .D(n30510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(CLK_c), 
           .D(n30509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(CLK_c), 
           .D(n30508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n30507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n30505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n30504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n30503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n30502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n30500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n30499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n30498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n30497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n30496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n30495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n30494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n30493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n30492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n30491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n30490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n30489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n30488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n30487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n30486));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n30485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n30484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n30483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n30482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i218 (.Q(\data_out_frame[27][1] ), .C(CLK_c), 
           .D(n30481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n30480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n30479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n30478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n30477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n30476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n30475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n30474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n30473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n30472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n30471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n30470));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n30469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n30468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n30467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n30466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n30465));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n30464));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n30463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n30462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n30461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n30460));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n30459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n30458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n30457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n30456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n30455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n30454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n30453));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n30452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n30451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n30450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n30449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n30448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n30447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n30446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n30445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n30444));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n30443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n30442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n30441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n30440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n30439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n30438));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(n29293), .I1(\data_out_frame[9] [4]), 
            .I2(n45770), .I3(GND_net), .O(n45743));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n30437));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[12] [0]), .I3(GND_net), .O(n46237));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n30436));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n30435));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n18_adj_4643));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n30434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n30433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n30432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n30431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n30430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n30429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n30428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n30427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n30426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n30425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n30424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n30423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n30422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n30421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n30420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n30419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n30418));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1388 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[5] [1]), .O(n29293));
    defparam i1_2_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n30417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n30416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n30415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n30414));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n45888));
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n30413));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n28510));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n30412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n30411));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n30410));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(n45678), .I3(\data_out_frame[8] [2]), .O(n46074));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1392 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(n45729), .O(n45685));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1393 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[5] [1]), .I3(\data_in_frame[5] [0]), .O(n6_adj_4639));
    defparam i1_2_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37145 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n52780));
    defparam byte_transmit_counter_0__bdd_4_lut_37145.LUT_INIT = 16'he4aa;
    SB_LUT4 n52780_bdd_4_lut (.I0(n52780), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n52783));
    defparam n52780_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37136 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n52774));
    defparam byte_transmit_counter_0__bdd_4_lut_37136.LUT_INIT = 16'he4aa;
    SB_LUT4 n52774_bdd_4_lut (.I0(n52774), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n52777));
    defparam n52774_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n30409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n30408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n30407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n30406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n30405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n30404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n30403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n30402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n30401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n30400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n30399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n30398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n30397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n30396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n30395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n30394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n30393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n30392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n30391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n30390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n30389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n30388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n30387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n30386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n30385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n30384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n30383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n30382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n30381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n30380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n30379));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n30378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n30377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n30376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n30375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n30374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n30373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n30372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n30371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n30370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n30369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n30368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n30367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n30366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n30365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n30364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n30363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n30362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n30361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n30360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n30359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n30358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n30357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n30356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n30355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n30354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n30353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n30352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n30351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n30350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n30349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n30348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n30347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n30346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n30345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n30344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n30343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n30342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n30341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n30340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n30339));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n30338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n30337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n30336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n30335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n30334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n30333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n30332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n30331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n30330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n30329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n30328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n30327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n30326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n30325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n30324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n30323));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_4_lut (.I0(n45709), .I1(\data_out_frame[12] [1]), .I2(n13_adj_4649), 
            .I3(n14_adj_4648), .O(n45970));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n30322));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1394 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[4] [6]), .O(n45770));
    defparam i1_2_lut_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n30321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n30320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n30319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n30318));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n30317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n30316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n30124));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[14] [3]), 
            .I2(n45970), .I3(GND_net), .O(n46151));
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1396 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n6_adj_4636));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1396.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n30315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n30314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n30313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n30312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n30311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n30310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n30309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n30308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n30307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n30306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n30305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n30304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n30303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n30302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n30301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n30300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n30299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n30298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n30297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n30296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n30295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n30294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n30293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n30292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n30291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n30290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n30289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n30288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n30287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n30286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n30285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n30284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n30283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n30282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n30281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n30280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n30279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n30278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n30277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n30276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n30275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n30274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n30273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n30272));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[14] [7]), 
            .I2(n45824), .I3(GND_net), .O(n6_adj_4632));
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(n29091), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n45752));
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n29034));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n46246));
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [5]), .O(n45712));
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n46127));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1403 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[15] [1]), 
            .O(n45841));
    defparam i1_2_lut_3_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i16730_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n30419));
    defparam i16730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16731_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n30420));
    defparam i16731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35725_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), 
            .I2(tx_transmit_N_3513), .I3(\FRAME_MATCHER.state [0]), .O(n51044));   // verilog/coms.v(145[4] 299[11])
    defparam i35725_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(n43663), .I1(n160), .I2(n45614), 
            .I3(GND_net), .O(n32424));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'hfefe;
    SB_LUT4 i22866_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n67), .I3(GND_net), .O(n36547));
    defparam i22866_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i16732_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n30421));
    defparam i16732_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_rep_64_2_lut (.I0(n43017), .I1(n29255), .I2(GND_net), .I3(GND_net), 
            .O(n53041));
    defparam i1_rep_64_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16733_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n30422));
    defparam i16733_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1405 (.I0(n54), .I1(n45635), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(n54_c), .O(n29618));
    defparam i2_3_lut_4_lut_adj_1405.LUT_INIT = 16'h0010;
    SB_LUT4 i16734_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n30423));
    defparam i16734_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16735_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n30424));
    defparam i16735_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut (.I0(n28113), .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[9] [4]), 
            .I3(\data_out_frame[9] [3]), .O(n14_adj_4545));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1406 (.I0(\data_out_frame[16] [4]), .I1(n43854), 
            .I2(n43121), .I3(\data_out_frame[23] [1]), .O(n45939));
    defparam i2_3_lut_4_lut_adj_1406.LUT_INIT = 16'h9669;
    SB_LUT4 i16736_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n30425));
    defparam i16736_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n67), .O(n29783));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2_3_lut_4_lut_adj_1407 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [4]), 
            .I2(n27987), .I3(n47174), .O(n46005));
    defparam i2_3_lut_4_lut_adj_1407.LUT_INIT = 16'h9669;
    SB_LUT4 i5_2_lut_4_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[6] [3]), .O(n16_adj_4642));   // verilog/coms.v(75[16:43])
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1408 (.I0(n45904), .I1(n43017), .I2(n29255), 
            .I3(GND_net), .O(n6_adj_4694));
    defparam i2_3_lut_adj_1408.LUT_INIT = 16'h6969;
    SB_LUT4 i5_3_lut_4_lut_adj_1409 (.I0(n29458), .I1(\data_out_frame[11] [4]), 
            .I2(n10_adj_4537), .I3(n46039), .O(n42930));
    defparam i5_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i16737_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n30426));
    defparam i16737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(n25438), .I1(n42259), .I2(n771), 
            .I3(n117), .O(n45642));
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'hff02;
    SB_LUT4 i1_2_lut_4_lut_adj_1411 (.I0(n28941), .I1(n28113), .I2(\data_out_frame[17] [7]), 
            .I3(n43025), .O(n8_adj_4533));
    defparam i1_2_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1412 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[15] [6]), .I3(n43007), .O(n8_adj_4527));
    defparam i2_2_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1413 (.I0(\data_in_frame[19] [6]), .I1(n53041), 
            .I2(\data_in_frame[21] [7]), .I3(\data_in_frame[19] [5]), .O(n47172));
    defparam i3_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 equal_298_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4693));   // verilog/coms.v(154[7:23])
    defparam equal_298_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1414 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n29147));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 equal_297_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4695));   // verilog/coms.v(154[7:23])
    defparam equal_297_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n45801));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n30271));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1416 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(n45961), .O(n28595));
    defparam i1_2_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i16722_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n30411));
    defparam i16722_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16723_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n30412));
    defparam i16723_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16724_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n30413));
    defparam i16724_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16725_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n30414));
    defparam i16725_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16726_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n30415));
    defparam i16726_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34455_4_lut (.I0(n47755), .I1(n10_adj_4686), .I2(n46219), 
            .I3(GND_net), .O(n50031));
    defparam i34455_4_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i16727_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n30416));
    defparam i16727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n30270));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16728_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n30417));
    defparam i16728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_3_lut_4_lut_adj_1417 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[14] [3]), .I3(n47669), .O(n11_adj_4518));
    defparam i4_3_lut_4_lut_adj_1417.LUT_INIT = 16'h9669;
    SB_LUT4 i16729_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n30418));
    defparam i16729_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22995_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4177));
    defparam i22995_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n6496));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 select_657_Select_1_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4626));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_2_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4624));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_3_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4622));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i4_2_lut_4_lut (.I0(n46231), .I1(n10_adj_4660), .I2(n47627), 
            .I3(\data_out_frame[19] [6]), .O(n43_adj_4515));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1418 (.I0(\data_in_frame[20] [5]), .I1(n45987), 
            .I2(\data_in_frame[18] [4]), .I3(Kp_23__N_1803), .O(n47094));
    defparam i3_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 select_657_Select_4_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4620));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[13] [1]), .I1(n27979), 
            .I2(\data_out_frame[15] [4]), .I3(\data_out_frame[15] [3]), 
            .O(n45862));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 select_657_Select_5_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4618));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_6_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4616));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_7_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4614));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_8_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4612));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_9_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4610));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_10_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4608));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_11_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4605));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_12_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4603));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_3_lut_adj_1420 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n29137));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1420.LUT_INIT = 16'h9696;
    SB_LUT4 select_657_Select_13_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4601));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_14_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4599));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_15_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4597));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i22846_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n36526));
    defparam i22846_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_657_Select_16_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4595));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_17_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4593));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i34449_4_lut (.I0(\data_in_frame[21] [0]), .I1(n47172), .I2(n6_adj_4694), 
            .I3(n45885), .O(n50025));
    defparam i34449_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_657_Select_18_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4591));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_19_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4589));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_20_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4587));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i4_4_lut_adj_1421 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[19] [3]), 
            .I2(n47973), .I3(n6_adj_4687), .O(n46996));
    defparam i4_4_lut_adj_1421.LUT_INIT = 16'h9669;
    SB_LUT4 select_657_Select_21_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4586));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_22_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4585));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_23_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4584));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_24_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4583));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_25_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4582));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 equal_288_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4697));
    defparam equal_288_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2859_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8));
    defparam i2859_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 select_657_Select_26_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4581));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_27_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4580));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_28_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4579));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_29_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4578));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_30_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4577));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_31_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4576));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 select_657_Select_0_i3_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), 
            .I1(n36474), .I2(n28426), .I3(\FRAME_MATCHER.i [0]), .O(n3));   // verilog/coms.v(112[11:16])
    defparam select_657_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n45936), .I3(GND_net), .O(n42655));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n46064), .I3(GND_net), .O(n6_adj_4458));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 i16714_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n30403));
    defparam i16714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16715_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n30404));
    defparam i16715_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16716_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n30405));
    defparam i16716_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16717_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n30406));
    defparam i16717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_adj_1424 (.I0(n63_adj_3), .I1(n771), .I2(n7_adj_4690), 
            .I3(n42259), .O(n5_adj_4));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut_adj_1424.LUT_INIT = 16'ha0a2;
    SB_LUT4 i16718_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n30407));
    defparam i16718_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16719_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n30408));
    defparam i16719_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1425 (.I0(n43797), .I1(n49), .I2(n6_adj_4688), 
            .I3(n43795), .O(n26_adj_4699));
    defparam i8_4_lut_adj_1425.LUT_INIT = 16'hedde;
    SB_LUT4 i16720_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n30409));
    defparam i16720_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1426 (.I0(n29188), .I1(n28870), .I2(n45910), 
            .I3(n45991), .O(n42954));
    defparam i1_2_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i16721_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n30410));
    defparam i16721_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1427 (.I0(tx_transmit_N_3513), .I1(n2025), 
            .I2(n25438), .I3(n28383), .O(n94));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut_adj_1427.LUT_INIT = 16'h00e0;
    SB_LUT4 i14_4_lut_adj_1428 (.I0(n50025), .I1(n47094), .I2(n50031), 
            .I3(n9), .O(n32));
    defparam i14_4_lut_adj_1428.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(n1[1]), .I1(n63_adj_3), .I2(n45649), 
            .I3(GND_net), .O(n44890));   // verilog/coms.v(142[4] 144[7])
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'hb0b0;
    SB_LUT4 i2_2_lut_3_lut_adj_1430 (.I0(\data_out_frame[15] [5]), .I1(n29389), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n45696));
    defparam i2_2_lut_3_lut_adj_1430.LUT_INIT = 16'h9696;
    SB_LUT4 i16706_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n30395));
    defparam i16706_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16707_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n30396));
    defparam i16707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_4_lut_adj_1431 (.I0(n160), .I1(n21_adj_4551), .I2(n19_adj_4550), 
            .I3(n20_adj_4549), .O(n8_adj_4571));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 i16708_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n30397));
    defparam i16708_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1432 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [2]), 
            .I2(n43889), .I3(\data_in_frame[21] [4]), .O(n47851));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1432.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1433 (.I0(n29188), .I1(n28870), .I2(n45910), 
            .I3(GND_net), .O(n45827));
    defparam i1_2_lut_3_lut_adj_1433.LUT_INIT = 16'h9696;
    SB_LUT4 i16709_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n30398));
    defparam i16709_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16710_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n30399));
    defparam i16710_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16711_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n30400));
    defparam i16711_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16712_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n30401));
    defparam i16712_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16713_3_lut_4_lut (.I0(n36526), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n30402));
    defparam i16713_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1434 (.I0(n45491), .I1(n28389), .I2(n58), 
            .I3(n45670), .O(n28383));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1434.LUT_INIT = 16'hffef;
    SB_LUT4 i16698_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n30387));
    defparam i16698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16699_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n30388));
    defparam i16699_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16700_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n30389));
    defparam i16700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16701_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n30390));
    defparam i16701_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16702_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n30391));
    defparam i16702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16703_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n30392));
    defparam i16703_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16704_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n30393));
    defparam i16704_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16705_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n30394));
    defparam i16705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16690_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n30379));
    defparam i16690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16691_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n30380));
    defparam i16691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16692_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n30381));
    defparam i16692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16693_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n30382));
    defparam i16693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16694_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n30383));
    defparam i16694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16695_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n30384));
    defparam i16695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16696_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n30385));
    defparam i16696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16697_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n30386));
    defparam i16697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18451_3_lut (.I0(\data_out_frame[20]_c [4]), .I1(\displacement[4] ), 
            .I2(n25701), .I3(GND_net), .O(n30524));
    defparam i18451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(n29091), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n45846));
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1436 (.I0(n29091), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n46276));
    defparam i1_2_lut_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1437 (.I0(\data_in_frame[4] [5]), .I1(n28750), 
            .I2(n29137), .I3(GND_net), .O(n29188));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1437.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1438 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n28870));
    defparam i1_2_lut_3_lut_adj_1438.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[19] [6]), 
            .I2(n45777), .I3(\data_out_frame[22] [0]), .O(n46061));
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1440 (.I0(\data_in_frame[4] [5]), .I1(Kp_23__N_1020), 
            .I2(n45916), .I3(n46249), .O(n29210));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1441 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(\data_out_frame[20] [5]), 
            .O(n46095));
    defparam i2_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i16682_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n30371));
    defparam i16682_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1442 (.I0(n45947), .I1(n47698), .I2(n43858), 
            .I3(\data_out_frame[22] [3]), .O(n14_adj_4492));
    defparam i5_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i16683_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n30372));
    defparam i16683_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16684_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n30373));
    defparam i16684_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16685_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n30374));
    defparam i16685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1443 (.I0(\data_out_frame[24] [5]), .I1(n43906), 
            .I2(n10_adj_4489), .I3(n28003), .O(n48289));
    defparam i5_3_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(n45721), .I1(n46095), .I2(n43803), 
            .I3(\data_out_frame[20][0] ), .O(n47041));
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i16686_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n30375));
    defparam i16686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16687_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n30376));
    defparam i16687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16688_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n30377));
    defparam i16688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16689_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n30378));
    defparam i16689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(n45824), .I3(n43910), .O(n46263));
    defparam i1_3_lut_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1446 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(n46253), .I3(\data_out_frame[6] [6]), .O(n4_adj_4543));   // verilog/coms.v(76[16:27])
    defparam i1_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n46112));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1448 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[4] [6]), .O(n29458));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1449 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[4] [5]), .I3(\data_out_frame[6] [7]), .O(n46253));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i16674_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n30363));
    defparam i16674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[1] [6]), .O(n46184));   // verilog/coms.v(96[12:25])
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n46266));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i16675_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n30364));
    defparam i16675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1452 (.I0(n7_adj_4689), .I1(n47973), .I2(n43899), 
            .I3(n45930), .O(n47333));
    defparam i4_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i16676_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n30365));
    defparam i16676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16762_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n30451));
    defparam i16762_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16763_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n30452));
    defparam i16763_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16677_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n30366));
    defparam i16677_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16678_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n30367));
    defparam i16678_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16679_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n30368));
    defparam i16679_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16680_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n30369));
    defparam i16680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16764_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n30453));
    defparam i16764_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16681_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n30370));
    defparam i16681_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(n29458), .I3(GND_net), .O(n6_adj_4535));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1454 (.I0(n45987), .I1(n46133), .I2(\data_in_frame[20] [4]), 
            .I3(GND_net), .O(n47097));
    defparam i2_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i16765_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n30454));
    defparam i16765_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1455 (.I0(\data_out_frame[23] [5]), .I1(n43816), 
            .I2(n47627), .I3(\data_out_frame[25] [7]), .O(n6_adj_4481));
    defparam i1_2_lut_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1456 (.I0(n45709), .I1(n45814), .I2(\data_out_frame[14] [4]), 
            .I3(n45846), .O(n29380));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1457 (.I0(n45709), .I1(n45814), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[16] [6]), .O(n45976));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i16766_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n30455));
    defparam i16766_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16666_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n30355));
    defparam i16666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16767_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n30456));
    defparam i16767_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16667_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n30356));
    defparam i16667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16668_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n30357));
    defparam i16668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16669_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n30358));
    defparam i16669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16670_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n30359));
    defparam i16670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16768_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n30457));
    defparam i16768_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1458 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n6_adj_4479));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1458.LUT_INIT = 16'h9696;
    SB_LUT4 i16671_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n30360));
    defparam i16671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16672_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n30361));
    defparam i16672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16673_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n30362));
    defparam i16673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(n43940), .I1(n46151), .I2(\data_out_frame[19] [0]), 
            .I3(n45846), .O(n43121));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_4_lut_adj_1460 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[1] [6]), .I3(n45795), .O(n8_adj_4478));   // verilog/coms.v(78[16:27])
    defparam i3_3_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[1] [3]), 
            .I2(n45952), .I3(n28595), .O(n28827));
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1462 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[3] [6]), .O(n45795));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1463 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(n29137), .I3(GND_net), .O(n45758));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1464 (.I0(\data_in_frame[4] [5]), .I1(n28750), 
            .I2(n10_adj_4472), .I3(n45758), .O(n8_adj_4429));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1465 (.I0(n9_adj_4471), .I1(n7_adj_4470), 
            .I2(n8_adj_4468), .I3(n9), .O(n61));
    defparam i1_2_lut_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1466 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(n46107), .I3(GND_net), .O(n46260));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1467 (.I0(\data_in_frame[9] [1]), .I1(n28776), 
            .I2(n8_adj_4429), .I3(GND_net), .O(n45817));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1467.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1468 (.I0(\data_in_frame[9] [2]), .I1(n43430), 
            .I2(n29226), .I3(GND_net), .O(n10_adj_4465));
    defparam i2_2_lut_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(\data_out_frame[18] [5]), .I1(n28910), 
            .I2(\data_out_frame[20] [6]), .I3(n43940), .O(n48169));
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i62_3_lut (.I0(n46), .I1(n4452), .I2(n25438), .I3(GND_net), 
            .O(n3_adj_4661));   // verilog/coms.v(115[11:12])
    defparam i62_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i30925_4_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n42507), .I2(n28276), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n46495));
    defparam i30925_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[18] [5]), .I1(n28910), 
            .I2(n43816), .I3(GND_net), .O(n6_adj_4637));
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i16475_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45626), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n30164));
    defparam i16475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1471 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n35635), .O(n45654));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1471.LUT_INIT = 16'hefff;
    SB_LUT4 i16658_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n30347));
    defparam i16658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(\FRAME_MATCHER.state_c [31]), .I1(n11_adj_4663), 
            .I2(GND_net), .I3(GND_net), .O(n44886));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\FRAME_MATCHER.state_c [31]), .I1(n3_adj_4661), 
            .I2(GND_net), .I3(GND_net), .O(n45580));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h8888;
    SB_LUT4 i16659_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n30348));
    defparam i16659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16660_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30349));
    defparam i16660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16661_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n30350));
    defparam i16661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16662_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30351));
    defparam i16662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16663_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30352));
    defparam i16663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1474 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n35635), .O(n45626));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1474.LUT_INIT = 16'hfeff;
    SB_LUT4 i16664_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30353));
    defparam i16664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16665_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30354));
    defparam i16665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1475 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[13] [2]), 
            .O(n14_adj_4525));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1476 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(n46178), .I3(GND_net), .O(n6_adj_4629));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n26683));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1478 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_988), .I3(GND_net), .O(n27216));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1478.LUT_INIT = 16'h9696;
    SB_LUT4 i16650_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n30339));
    defparam i16650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16651_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n30340));
    defparam i16651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16652_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n30341));
    defparam i16652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16653_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n30342));
    defparam i16653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16654_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n30343));
    defparam i16654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37131 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n52762));
    defparam byte_transmit_counter_0__bdd_4_lut_37131.LUT_INIT = 16'he4aa;
    SB_LUT4 i16655_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n30344));
    defparam i16655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16656_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n30345));
    defparam i16656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16657_3_lut_4_lut (.I0(n8_adj_4697), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n30346));
    defparam i16657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16642_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n30331));
    defparam i16642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16643_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n30332));
    defparam i16643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16644_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n30333));
    defparam i16644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16645_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n30334));
    defparam i16645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1479 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n43846), .I3(\data_out_frame[18] [3]), .O(n46187));
    defparam i1_2_lut_4_lut_adj_1479.LUT_INIT = 16'h9669;
    SB_LUT4 i16646_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n30335));
    defparam i16646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16647_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n30336));
    defparam i16647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16648_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n30337));
    defparam i16648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16649_3_lut_4_lut (.I0(n36526), .I1(n45654), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n30338));
    defparam i16649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16634_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n30323));
    defparam i16634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16635_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n30324));
    defparam i16635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16636_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n30325));
    defparam i16636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16637_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n30326));
    defparam i16637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16638_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n30327));
    defparam i16638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16639_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n30328));
    defparam i16639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16640_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n30329));
    defparam i16640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16641_3_lut_4_lut (.I0(n8_adj_4692), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n30330));
    defparam i16641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1480 (.I0(n45491), .I1(n45670), .I2(n58), 
            .I3(n28389), .O(n36474));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1481 (.I0(\data_in_frame[8] [4]), .I1(n28776), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n12_adj_4463));
    defparam i1_2_lut_3_lut_adj_1481.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1482 (.I0(n42921), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n46064));
    defparam i1_2_lut_3_lut_adj_1482.LUT_INIT = 16'h9696;
    SB_LUT4 i16626_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n30315));
    defparam i16626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1483 (.I0(n28870), .I1(n45910), .I2(n46077), 
            .I3(GND_net), .O(n6_adj_4454));   // verilog/coms.v(96[12:25])
    defparam i1_2_lut_3_lut_adj_1483.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1484 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [6]), .I3(GND_net), .O(n46166));
    defparam i1_2_lut_3_lut_adj_1484.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1485 (.I0(\data_in_frame[21] [2]), .I1(n45904), 
            .I2(\data_in_frame[19] [1]), .I3(n27975), .O(n47108));
    defparam i3_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1486 (.I0(n43795), .I1(n43606), .I2(\data_in_frame[17] [0]), 
            .I3(GND_net), .O(n43889));
    defparam i1_2_lut_3_lut_adj_1486.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1487 (.I0(n28809), .I1(n28892), .I2(\data_in_frame[10] [4]), 
            .I3(\data_in_frame[14] [6]), .O(n46203));
    defparam i2_3_lut_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i16627_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n30316));
    defparam i16627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(n42988), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[16] [7]), .I3(\data_in_frame[12] [5]), .O(n45999));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1489 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[10] [6]), 
            .I2(n10_adj_4442), .I3(n46273), .O(n43797));
    defparam i5_3_lut_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i16628_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n30317));
    defparam i16628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1490 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[8] [6]), 
            .I2(\data_in_frame[15] [2]), .I3(GND_net), .O(n6_adj_4441));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1490.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(\data_in_frame[16] [3]), .I1(n48165), 
            .I2(n46107), .I3(\data_in_frame[16] [4]), .O(n43876));
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h9669;
    SB_LUT4 i26704_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n45), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n42261));
    defparam i26704_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_3_lut_4_lut_adj_1492 (.I0(n8_adj_4692), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n28400), .I3(\FRAME_MATCHER.i [3]), .O(n28276));
    defparam i1_3_lut_4_lut_adj_1492.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_1493 (.I0(\data_in_frame[20] [3]), .I1(n46133), 
            .I2(n43862), .I3(\data_in_frame[18] [1]), .O(n47090));
    defparam i3_4_lut_adj_1493.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1494 (.I0(\data_in_frame[18] [1]), .I1(n47169), 
            .I2(\data_in_frame[20] [2]), .I3(n43222), .O(n24_adj_4459));
    defparam i6_4_lut_adj_1494.LUT_INIT = 16'hedde;
    SB_LUT4 i22542_3_lut_3_lut (.I0(n28494), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36220));
    defparam i22542_3_lut_3_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n45), .I3(GND_net), .O(n46));
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'hfdfd;
    SB_LUT4 n52762_bdd_4_lut (.I0(n52762), .I1(\data_out_frame[21][3] ), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n52765));
    defparam n52762_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i26702_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n45), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(GND_net), .O(n42259));
    defparam i26702_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1496 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n28494), .I3(n62), .O(n47127));
    defparam i2_3_lut_4_lut_adj_1496.LUT_INIT = 16'hfff7;
    SB_LUT4 i16629_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n30318));
    defparam i16629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16630_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n30319));
    defparam i16630_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16631_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n30320));
    defparam i16631_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37155 (.I0(byte_transmit_counter[1]), 
            .I1(n50268), .I2(n50269), .I3(byte_transmit_counter[2]), .O(n52756));
    defparam byte_transmit_counter_1__bdd_4_lut_37155.LUT_INIT = 16'he4aa;
    SB_LUT4 i16632_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n30321));
    defparam i16632_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16633_3_lut_4_lut (.I0(n8_adj_4667), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n30322));
    defparam i16633_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n52756_bdd_4_lut (.I0(n52756), .I1(n50257), .I2(n50256), .I3(byte_transmit_counter[2]), 
            .O(n52759));
    defparam n52756_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16618_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n30307));
    defparam i16618_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37117 (.I0(byte_transmit_counter[1]), 
            .I1(n50280), .I2(n50281), .I3(byte_transmit_counter[2]), .O(n52750));
    defparam byte_transmit_counter_1__bdd_4_lut_37117.LUT_INIT = 16'he4aa;
    SB_LUT4 n52750_bdd_4_lut (.I0(n52750), .I1(n50278), .I2(n50277), .I3(byte_transmit_counter[2]), 
            .O(n52753));
    defparam n52750_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16619_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n30308));
    defparam i16619_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16620_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n30309));
    defparam i16620_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16621_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n30310));
    defparam i16621_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16622_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n30311));
    defparam i16622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16623_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n30312));
    defparam i16623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16624_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n30313));
    defparam i16624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16625_3_lut_4_lut (.I0(n8_adj_4670), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n30314));
    defparam i16625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i37090_2_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n32424), .O(n46478));
    defparam i37090_2_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16610_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n30299));
    defparam i16610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16611_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n30300));
    defparam i16611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16612_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n30301));
    defparam i16612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16613_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n30302));
    defparam i16613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16614_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n30303));
    defparam i16614_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_37122 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n52744));
    defparam byte_transmit_counter_0__bdd_4_lut_37122.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_adj_1497 (.I0(\FRAME_MATCHER.state_31__N_2724 [3]), .I1(n32424), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4700));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_adj_1497.LUT_INIT = 16'h2222;
    SB_LUT4 i16615_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n30304));
    defparam i16615_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16616_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n30305));
    defparam i16616_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16617_3_lut_4_lut (.I0(n8_adj_4674), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n30306));
    defparam i16617_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16602_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n30291));
    defparam i16602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1498 (.I0(n7_adj_4700), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(n46329), .I3(\FRAME_MATCHER.state[3] ), .O(n25701));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1498.LUT_INIT = 16'h0008;
    SB_LUT4 i37082_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n29930));
    defparam i37082_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i16603_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n30292));
    defparam i16603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16604_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n30293));
    defparam i16604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16605_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n30294));
    defparam i16605_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n52744_bdd_4_lut (.I0(n52744), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n52747));
    defparam n52744_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16606_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n30295));
    defparam i16606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16607_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n30296));
    defparam i16607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16608_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n30297));
    defparam i16608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16609_3_lut_4_lut (.I0(n8_adj_4693), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n30298));
    defparam i16609_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16594_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n30283));
    defparam i16594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16595_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n30284));
    defparam i16595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16596_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n30285));
    defparam i16596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16597_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n30286));
    defparam i16597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16598_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n30287));
    defparam i16598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16599_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n30288));
    defparam i16599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(n45693), .I2(\data_in_frame[1] [4]), 
            .I3(n29137), .O(n20));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0090;
    SB_LUT4 i16600_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n30289));
    defparam i16600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_37112 (.I0(byte_transmit_counter[1]), 
            .I1(n50241), .I2(n50242), .I3(byte_transmit_counter[2]), .O(n52738));
    defparam byte_transmit_counter_1__bdd_4_lut_37112.LUT_INIT = 16'he4aa;
    SB_LUT4 n52738_bdd_4_lut (.I0(n52738), .I1(n50239), .I2(n50238), .I3(byte_transmit_counter[2]), 
            .O(n52741));
    defparam n52738_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16601_3_lut_4_lut (.I0(n8_adj_4695), .I1(n45616), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n30290));
    defparam i16601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_3_lut_4_lut_adj_1499 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(Kp_23__N_969), .I3(\data_in_frame[2] [1]), .O(n17));
    defparam i4_3_lut_4_lut_adj_1499.LUT_INIT = 16'h0990;
    SB_LUT4 i34451_4_lut (.I0(n46949), .I1(\data_in_frame[19] [7]), .I2(n6_adj_4691), 
            .I3(\data_in_frame[20] [1]), .O(n50027));
    defparam i34451_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16_4_lut_adj_1500 (.I0(n47851), .I1(n32), .I2(n26_adj_4699), 
            .I3(n46996), .O(n34));
    defparam i16_4_lut_adj_1500.LUT_INIT = 16'hfeff;
    uart_tx tx (.CLK_c(CLK_c), .\r_SM_Main_2__N_3616[0] (r_SM_Main_2__N_3616[0]), 
            .r_SM_Main({r_SM_Main}), .n20694(n20694), .GND_net(GND_net), 
            .r_Bit_Index({Open_36, Open_37, \r_Bit_Index[0] }), .tx_o(tx_o), 
            .tx_data({tx_data}), .n29684(n29684), .n45512(n45512), .\r_SM_Main_2__N_3613[1] (\r_SM_Main_2__N_3613[1] ), 
            .n53023(n53023), .n30173(n30173), .tx_active(tx_active), .n4(n4), 
            .n30186(n30186), .VCC_net(VCC_net), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.CLK_c(CLK_c), .n29701(n29701), .n4(n4_adj_5), .GND_net(GND_net), 
            .n4_adj_1(n4_adj_6), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_7 ), 
            .n28484(n28484), .n35741(n35741), .r_SM_Main({r_SM_Main_adj_12}), 
            .r_Rx_Data(r_Rx_Data), .\r_SM_Main_2__N_3542[2] (\r_SM_Main_2__N_3542[2] ), 
            .RX_N_10(RX_N_10), .n28489(n28489), .n4_adj_2(n4_adj_11), 
            .n30197(n30197), .rx_data({rx_data}), .n45507(n45507), .n30156(n30156), 
            .n30155(n30155), .n30154(n30154), .n30153(n30153), .n30152(n30152), 
            .n30151(n30151), .n30150(n30150), .n45602(n45602), .n29660(n29660), 
            .n30189(n30189), .n45162(n45162), .rx_data_ready(rx_data_ready), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (CLK_c, \r_SM_Main_2__N_3616[0] , r_SM_Main, n20694, 
            GND_net, r_Bit_Index, tx_o, tx_data, n29684, n45512, 
            \r_SM_Main_2__N_3613[1] , n53023, n30173, tx_active, n4, 
            n30186, VCC_net, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    input \r_SM_Main_2__N_3616[0] ;
    output [2:0]r_SM_Main;
    output n20694;
    input GND_net;
    output [2:0]r_Bit_Index;
    output tx_o;
    input [7:0]tx_data;
    output n29684;
    output n45512;
    output \r_SM_Main_2__N_3613[1] ;
    input n53023;
    input n30173;
    output tx_active;
    output n4;
    input n30186;
    input VCC_net;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n30054;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n50229, n50230, n50233, n50232, n3, n25529, n20844;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index_c;   // verilog/uart_tx.v(33[16:27])
    
    wire n29963, n3_adj_4407, n20843, n46344, o_Tx_Serial_N_3644, 
        n52828, n46999, n10, n41871, n41870, n41869, n41868, n41867, 
        n41866, n41865, n41864;
    
    SB_DFFESR r_Clock_Count_2200__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2200__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i7147_2_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n20694));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7147_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34595_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n50229));
    defparam i34595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34596_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n50230));
    defparam i34596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34599_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n50233));
    defparam i34599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34598_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n50232));
    defparam i34598_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n25529), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n20844), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(CLK_c), .E(n29684), 
            .D(n307[1]), .R(n29963));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(CLK_c), .E(n29684), 
            .D(n307[2]), .R(n29963));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4407), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n25529), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n25529), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n25529), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n25529), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n25529), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n25529), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n25529), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2362_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2362_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2355_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2355_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45512));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7292_3_lut (.I0(n20843), .I1(\r_SM_Main_2__N_3613[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n20844));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7292_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i30780_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n46344));
    defparam i30780_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3644), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index_c[1]), .I1(n50232), 
            .I2(n50233), .I3(r_Bit_Index_c[2]), .O(n52828));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n52828_bdd_4_lut (.I0(n52828), .I1(n50230), .I2(n50229), .I3(r_Bit_Index_c[2]), 
            .O(o_Tx_Serial_N_3644));
    defparam n52828_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut (.I0(n45512), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(n46344), .O(n29963));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFFESR r_Clock_Count_2200__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n30054));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i7291_3_lut_4_lut (.I0(n45512), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3616[0] ), .O(n20843));
    defparam i7291_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 i11614_2_lut_3_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4407));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i11614_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n53023));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n30173));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n46999));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n46999), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3613[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i36395_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n30054));
    defparam i36395_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n30186));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_2200_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n41871), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2200_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n41870), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_9 (.CI(n41870), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n41871));
    SB_LUT4 r_Clock_Count_2200_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n41869), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_8 (.CI(n41869), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n41870));
    SB_LUT4 r_Clock_Count_2200_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n41868), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_7 (.CI(n41868), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n41869));
    SB_LUT4 r_Clock_Count_2200_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n41867), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_6 (.CI(n41867), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n41868));
    SB_LUT4 r_Clock_Count_2200_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n41866), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_5 (.CI(n41866), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n41867));
    SB_LUT4 r_Clock_Count_2200_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n41865), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_4 (.CI(n41865), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n41866));
    SB_LUT4 r_Clock_Count_2200_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n41864), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_3 (.CI(n41864), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n41865));
    SB_LUT4 r_Clock_Count_2200_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2200_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2200_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n41864));
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3616[0] ), .O(n25529));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_4_lut_adj_866 (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n29684));
    defparam i1_3_lut_4_lut_adj_866.LUT_INIT = 16'h0203;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (CLK_c, n29701, n4, GND_net, n4_adj_1, \r_Bit_Index[0] , 
            n28484, n35741, r_SM_Main, r_Rx_Data, \r_SM_Main_2__N_3542[2] , 
            RX_N_10, n28489, n4_adj_2, n30197, rx_data, n45507, 
            n30156, n30155, n30154, n30153, n30152, n30151, n30150, 
            n45602, n29660, n30189, n45162, rx_data_ready, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n29701;
    output n4;
    input GND_net;
    output n4_adj_1;
    output \r_Bit_Index[0] ;
    output n28484;
    output n35741;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    output \r_SM_Main_2__N_3542[2] ;
    input RX_N_10;
    output n28489;
    output n4_adj_2;
    input n30197;
    output [7:0]rx_data;
    output n45507;
    input n30156;
    input n30155;
    input n30154;
    input n30153;
    input n30152;
    input n30151;
    input n30150;
    input n45602;
    output n29660;
    input n30189;
    input n45162;
    output rx_data_ready;
    input VCC_net;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n37;
    
    wire n29789;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n30052;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n29972, n28243;
    wire [2:0]r_SM_Main_2__N_3548;
    
    wire n51101, n36644, n52897, r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n52894, n9, n28272, n6, n51126, n51124, n6_adj_4406, 
        n41863, n41862, n41861, n41860, n41859, n41858, n41857;
    
    SB_DFFESR r_Clock_Count_2198__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n29789), 
            .D(n37[7]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n29789), 
            .D(n37[6]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n29789), 
            .D(n37[5]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n29789), 
            .D(n37[4]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n29789), 
            .D(n37[3]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n29789), 
            .D(n37[2]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2198__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n29789), 
            .D(n37[1]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n29701), 
            .D(n326[1]), .R(n29972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_331_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_331_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_330_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_330_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n29701), 
            .D(n326[2]), .R(n29972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(n28243), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28484));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i22065_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35741));
    defparam i22065_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35688_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n51101));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i35688_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n51101), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n36644));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFESR r_Clock_Count_2198__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n29789), 
            .D(n37[0]), .R(n30052));   // verilog/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n52897), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n36644), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n28243));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_861 (.I0(n28243), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28489));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_861.LUT_INIT = 16'heeee;
    SB_LUT4 equal_333_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_333_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n30197));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2340_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2340_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n45507));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i22910_2_lut (.I0(n45507), .I1(\r_SM_Main_2__N_3542[2] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3545[0]));
    defparam i22910_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2333_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2333_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n52894_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_3548[0]), 
            .I3(n52894), .O(n52897));   // verilog/uart_rx.v(70[21:38])
    defparam n52894_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i3_4_lut_adj_862 (.I0(n9), .I1(r_Clock_Count[3]), .I2(n28272), 
            .I3(r_Clock_Count[1]), .O(r_SM_Main_2__N_3548[0]));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22857_4_lut (.I0(r_Clock_Count[0]), .I1(n28272), .I2(n6), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3542[2] ));
    defparam i22857_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3_2_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_863 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_Clock_Count[5]), .O(n28272));   // verilog/uart_rx.v(68[17:52])
    defparam i3_4_lut_adj_863.LUT_INIT = 16'hfffe;
    SB_LUT4 i35511_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n28272), 
            .I3(r_Clock_Count[3]), .O(n51126));
    defparam i35511_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i35701_3_lut (.I0(n51126), .I1(r_SM_Main[0]), .I2(n9), .I3(GND_net), 
            .O(n51124));
    defparam i35701_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n51124), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[1]), .O(n30052));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut_adj_864 (.I0(r_SM_Main_2__N_3548[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4406));
    defparam i2_2_lut_adj_864.LUT_INIT = 16'h4444;
    SB_LUT4 i36381_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4406), 
            .I3(r_Rx_Data), .O(n29789));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36381_4_lut.LUT_INIT = 16'h4555;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n30156));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n30155));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n30154));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n30153));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n30152));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n30151));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n30150));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n45602));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i13_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[0]), .O(n29660));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3542[2] ), 
            .I1(r_SM_Main[1]), .I2(n45507), .I3(r_SM_Main[0]), .O(n52894));
    defparam r_SM_Main_0__bdd_4_lut_4_lut_4_lut.LUT_INIT = 16'h7780;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n30189));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n45162));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_2198_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n41863), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2198_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n41862), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_8 (.CI(n41862), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n41863));
    SB_LUT4 r_Clock_Count_2198_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n41861), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_7 (.CI(n41861), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n41862));
    SB_LUT4 r_Clock_Count_2198_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n41860), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_6 (.CI(n41860), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n41861));
    SB_LUT4 r_Clock_Count_2198_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n41859), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_5 (.CI(n41859), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n41860));
    SB_LUT4 r_Clock_Count_2198_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n41858), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_4 (.CI(n41858), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n41859));
    SB_LUT4 r_Clock_Count_2198_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n41857), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_3 (.CI(n41857), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n41858));
    SB_LUT4 r_Clock_Count_2198_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2198_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2198_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n41857));
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3545[0]), .O(n29972));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_865 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3542[2] ), .O(n29701));
    defparam i1_3_lut_4_lut_adj_865.LUT_INIT = 16'h1101;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, pwm_setpoint, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input [23:0]pwm_setpoint;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire pwm_out_N_797;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n46962, n22, n15, n20, n24, n19, pwm_counter_23__N_795;
    wire [23:0]n101;
    
    wire n39, n41, n45, n43, n37, n29, n31, n23, n25, n35, 
        n33, n11, n13, n15_adj_4401, n27, n9, n17, n19_adj_4402, 
        n21, n51288, n51280, n12, n30, n51301, n51575, n51571, 
        n51890, n51704, n51937, n8, n6, n51736, n51737, n51224, 
        n16, n24_adj_4403, n10, n51271, n51226, n51796, n51506, 
        n4, n51728, n51729, n51275, n51860, n51508, n51965, n51966, 
        n51944, n51248, n51876, n51514, n51922, n41792, n41791, 
        n41790, n41789, n41788, n41787, n41786, n41785, n41784, 
        n41783, n41782, n41781, n41780, n41779, n41778, n41777, 
        n41776, n41775, n41774, n41773, n41772, n41771, n41770;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_797));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n46962));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[14]), .I2(pwm_counter[19]), 
            .I3(pwm_counter[17]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n46962), .I1(pwm_counter[22]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(pwm_counter[18]), .I3(pwm_counter[15]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[13]), .I1(pwm_counter[12]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i37092_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(pwm_counter_23__N_795));   // verilog/pwm.v(18[8:40])
    defparam i37092_4_lut.LUT_INIT = 16'h5554;
    SB_DFFSR pwm_counter_2189__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4401));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4402));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35654_4_lut (.I0(n21), .I1(n19_adj_4402), .I2(n17), .I3(n9), 
            .O(n51288));
    defparam i35654_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35646_4_lut (.I0(n27), .I1(n15_adj_4401), .I2(n13), .I3(n11), 
            .O(n51280));
    defparam i35646_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35940_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n51301), 
            .O(n51575));
    defparam i35940_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35936_4_lut (.I0(n19_adj_4402), .I1(n17), .I2(n15_adj_4401), 
            .I3(n51575), .O(n51571));
    defparam i35936_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36255_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n51571), 
            .O(n51890));
    defparam i36255_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36069_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n51890), 
            .O(n51704));
    defparam i36069_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36302_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n51704), 
            .O(n51937));
    defparam i36302_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36101_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n51736));   // verilog/pwm.v(21[8:24])
    defparam i36101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36102_3_lut (.I0(n51736), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n51737));   // verilog/pwm.v(21[8:24])
    defparam i36102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35590_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n51224));
    defparam i35590_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4403));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35637_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n51271));
    defparam i35637_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35592_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n51288), 
            .O(n51226));
    defparam i35592_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36161_4_lut (.I0(n24_adj_4403), .I1(n8), .I2(n45), .I3(n51224), 
            .O(n51796));   // verilog/pwm.v(21[8:24])
    defparam i36161_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35871_3_lut (.I0(n51737), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n51506));   // verilog/pwm.v(21[8:24])
    defparam i35871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i36093_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n51728));   // verilog/pwm.v(21[8:24])
    defparam i36093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36094_3_lut (.I0(n51728), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n51729));   // verilog/pwm.v(21[8:24])
    defparam i36094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35641_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n51280), 
            .O(n51275));
    defparam i35641_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36225_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n51271), 
            .O(n51860));   // verilog/pwm.v(21[8:24])
    defparam i36225_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35873_3_lut (.I0(n51729), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n51508));   // verilog/pwm.v(21[8:24])
    defparam i35873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36330_4_lut (.I0(n51508), .I1(n51860), .I2(n35), .I3(n51275), 
            .O(n51965));   // verilog/pwm.v(21[8:24])
    defparam i36330_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36331_3_lut (.I0(n51965), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n51966));   // verilog/pwm.v(21[8:24])
    defparam i36331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36309_3_lut (.I0(n51966), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n51944));   // verilog/pwm.v(21[8:24])
    defparam i36309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35614_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n51937), 
            .O(n51248));
    defparam i35614_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36241_4_lut (.I0(n51506), .I1(n51796), .I2(n45), .I3(n51226), 
            .O(n51876));   // verilog/pwm.v(21[8:24])
    defparam i36241_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35879_3_lut (.I0(n51944), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n51514));   // verilog/pwm.v(21[8:24])
    defparam i35879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36287_4_lut (.I0(n51514), .I1(n51876), .I2(n45), .I3(n51248), 
            .O(n51922));   // verilog/pwm.v(21[8:24])
    defparam i36287_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36288_3_lut (.I0(n51922), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_797));   // verilog/pwm.v(21[8:24])
    defparam i36288_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFSR pwm_counter_2189__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2189__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2189_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n41792), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2189_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n41791), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_24 (.CI(n41791), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n41792));
    SB_LUT4 pwm_counter_2189_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n41790), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_23 (.CI(n41790), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n41791));
    SB_LUT4 pwm_counter_2189_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n41789), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_22 (.CI(n41789), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n41790));
    SB_LUT4 pwm_counter_2189_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n41788), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_21 (.CI(n41788), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n41789));
    SB_LUT4 pwm_counter_2189_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n41787), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_20 (.CI(n41787), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n41788));
    SB_LUT4 pwm_counter_2189_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n41786), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_19 (.CI(n41786), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n41787));
    SB_LUT4 pwm_counter_2189_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n41785), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35667_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n51301));   // verilog/pwm.v(21[8:24])
    defparam i35667_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY pwm_counter_2189_add_4_18 (.CI(n41785), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n41786));
    SB_LUT4 pwm_counter_2189_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n41784), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_17 (.CI(n41784), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n41785));
    SB_LUT4 pwm_counter_2189_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n41783), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_16 (.CI(n41783), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n41784));
    SB_LUT4 pwm_counter_2189_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n41782), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_15 (.CI(n41782), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n41783));
    SB_LUT4 pwm_counter_2189_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n41781), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY pwm_counter_2189_add_4_14 (.CI(n41781), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n41782));
    SB_LUT4 pwm_counter_2189_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n41780), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_13 (.CI(n41780), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n41781));
    SB_LUT4 pwm_counter_2189_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n41779), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_12 (.CI(n41779), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n41780));
    SB_LUT4 pwm_counter_2189_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n41778), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_11 (.CI(n41778), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n41779));
    SB_LUT4 pwm_counter_2189_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n41777), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_10 (.CI(n41777), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n41778));
    SB_LUT4 pwm_counter_2189_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n41776), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_9 (.CI(n41776), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n41777));
    SB_LUT4 pwm_counter_2189_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n41775), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_8 (.CI(n41775), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n41776));
    SB_LUT4 pwm_counter_2189_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n41774), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_7 (.CI(n41774), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n41775));
    SB_LUT4 pwm_counter_2189_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n41773), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_6 (.CI(n41773), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n41774));
    SB_LUT4 pwm_counter_2189_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n41772), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_5 (.CI(n41772), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n41773));
    SB_LUT4 pwm_counter_2189_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n41771), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_4 (.CI(n41771), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n41772));
    SB_LUT4 pwm_counter_2189_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n41770), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_3 (.CI(n41770), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n41771));
    SB_LUT4 pwm_counter_2189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n41770));
    
endmodule
