// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 4 2020 19:52:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    input SDA;
    input SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__56636;
    wire N__56635;
    wire N__56634;
    wire N__56627;
    wire N__56626;
    wire N__56625;
    wire N__56618;
    wire N__56617;
    wire N__56616;
    wire N__56609;
    wire N__56608;
    wire N__56607;
    wire N__56600;
    wire N__56599;
    wire N__56598;
    wire N__56591;
    wire N__56590;
    wire N__56589;
    wire N__56582;
    wire N__56581;
    wire N__56580;
    wire N__56573;
    wire N__56572;
    wire N__56571;
    wire N__56564;
    wire N__56563;
    wire N__56562;
    wire N__56555;
    wire N__56554;
    wire N__56553;
    wire N__56546;
    wire N__56545;
    wire N__56544;
    wire N__56537;
    wire N__56536;
    wire N__56535;
    wire N__56528;
    wire N__56527;
    wire N__56526;
    wire N__56519;
    wire N__56518;
    wire N__56517;
    wire N__56510;
    wire N__56509;
    wire N__56508;
    wire N__56501;
    wire N__56500;
    wire N__56499;
    wire N__56492;
    wire N__56491;
    wire N__56490;
    wire N__56483;
    wire N__56482;
    wire N__56481;
    wire N__56474;
    wire N__56473;
    wire N__56472;
    wire N__56455;
    wire N__56452;
    wire N__56449;
    wire N__56446;
    wire N__56443;
    wire N__56440;
    wire N__56437;
    wire N__56436;
    wire N__56435;
    wire N__56434;
    wire N__56431;
    wire N__56430;
    wire N__56429;
    wire N__56424;
    wire N__56421;
    wire N__56418;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56404;
    wire N__56399;
    wire N__56392;
    wire N__56391;
    wire N__56390;
    wire N__56389;
    wire N__56388;
    wire N__56383;
    wire N__56382;
    wire N__56377;
    wire N__56376;
    wire N__56375;
    wire N__56374;
    wire N__56371;
    wire N__56368;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56354;
    wire N__56353;
    wire N__56350;
    wire N__56347;
    wire N__56344;
    wire N__56341;
    wire N__56336;
    wire N__56333;
    wire N__56330;
    wire N__56323;
    wire N__56320;
    wire N__56317;
    wire N__56314;
    wire N__56309;
    wire N__56302;
    wire N__56301;
    wire N__56300;
    wire N__56297;
    wire N__56296;
    wire N__56295;
    wire N__56294;
    wire N__56291;
    wire N__56286;
    wire N__56283;
    wire N__56278;
    wire N__56277;
    wire N__56276;
    wire N__56275;
    wire N__56272;
    wire N__56265;
    wire N__56260;
    wire N__56257;
    wire N__56256;
    wire N__56255;
    wire N__56254;
    wire N__56253;
    wire N__56252;
    wire N__56251;
    wire N__56250;
    wire N__56247;
    wire N__56244;
    wire N__56241;
    wire N__56238;
    wire N__56227;
    wire N__56224;
    wire N__56221;
    wire N__56216;
    wire N__56211;
    wire N__56206;
    wire N__56197;
    wire N__56196;
    wire N__56195;
    wire N__56194;
    wire N__56191;
    wire N__56188;
    wire N__56187;
    wire N__56184;
    wire N__56181;
    wire N__56180;
    wire N__56175;
    wire N__56174;
    wire N__56169;
    wire N__56166;
    wire N__56165;
    wire N__56162;
    wire N__56159;
    wire N__56156;
    wire N__56151;
    wire N__56146;
    wire N__56145;
    wire N__56142;
    wire N__56139;
    wire N__56134;
    wire N__56133;
    wire N__56130;
    wire N__56127;
    wire N__56124;
    wire N__56121;
    wire N__56118;
    wire N__56115;
    wire N__56112;
    wire N__56107;
    wire N__56098;
    wire N__56097;
    wire N__56096;
    wire N__56095;
    wire N__56094;
    wire N__56093;
    wire N__56092;
    wire N__56091;
    wire N__56090;
    wire N__56089;
    wire N__56088;
    wire N__56087;
    wire N__56086;
    wire N__56085;
    wire N__56084;
    wire N__56083;
    wire N__56082;
    wire N__56081;
    wire N__56080;
    wire N__56079;
    wire N__56078;
    wire N__56077;
    wire N__56076;
    wire N__56075;
    wire N__56074;
    wire N__56073;
    wire N__56072;
    wire N__56071;
    wire N__56070;
    wire N__56069;
    wire N__56068;
    wire N__56067;
    wire N__56066;
    wire N__56065;
    wire N__56064;
    wire N__56063;
    wire N__56062;
    wire N__56061;
    wire N__56060;
    wire N__56059;
    wire N__56058;
    wire N__56057;
    wire N__56056;
    wire N__56055;
    wire N__56054;
    wire N__56053;
    wire N__56052;
    wire N__56051;
    wire N__56050;
    wire N__56049;
    wire N__56048;
    wire N__56047;
    wire N__56046;
    wire N__56045;
    wire N__56044;
    wire N__56043;
    wire N__56042;
    wire N__56041;
    wire N__56040;
    wire N__56039;
    wire N__55918;
    wire N__55915;
    wire N__55912;
    wire N__55909;
    wire N__55908;
    wire N__55905;
    wire N__55902;
    wire N__55901;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55888;
    wire N__55887;
    wire N__55884;
    wire N__55879;
    wire N__55876;
    wire N__55873;
    wire N__55864;
    wire N__55861;
    wire N__55860;
    wire N__55859;
    wire N__55856;
    wire N__55855;
    wire N__55852;
    wire N__55849;
    wire N__55846;
    wire N__55843;
    wire N__55840;
    wire N__55837;
    wire N__55832;
    wire N__55829;
    wire N__55826;
    wire N__55823;
    wire N__55816;
    wire N__55813;
    wire N__55810;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55798;
    wire N__55795;
    wire N__55792;
    wire N__55789;
    wire N__55786;
    wire N__55783;
    wire N__55780;
    wire N__55777;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55767;
    wire N__55766;
    wire N__55763;
    wire N__55758;
    wire N__55755;
    wire N__55752;
    wire N__55747;
    wire N__55744;
    wire N__55741;
    wire N__55738;
    wire N__55735;
    wire N__55732;
    wire N__55729;
    wire N__55726;
    wire N__55723;
    wire N__55720;
    wire N__55717;
    wire N__55714;
    wire N__55713;
    wire N__55712;
    wire N__55711;
    wire N__55710;
    wire N__55709;
    wire N__55708;
    wire N__55707;
    wire N__55706;
    wire N__55703;
    wire N__55702;
    wire N__55701;
    wire N__55700;
    wire N__55699;
    wire N__55698;
    wire N__55697;
    wire N__55696;
    wire N__55695;
    wire N__55694;
    wire N__55685;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55673;
    wire N__55668;
    wire N__55657;
    wire N__55656;
    wire N__55655;
    wire N__55654;
    wire N__55653;
    wire N__55652;
    wire N__55651;
    wire N__55648;
    wire N__55645;
    wire N__55644;
    wire N__55641;
    wire N__55638;
    wire N__55633;
    wire N__55628;
    wire N__55623;
    wire N__55618;
    wire N__55615;
    wire N__55608;
    wire N__55605;
    wire N__55602;
    wire N__55599;
    wire N__55596;
    wire N__55587;
    wire N__55576;
    wire N__55567;
    wire N__55564;
    wire N__55563;
    wire N__55560;
    wire N__55557;
    wire N__55552;
    wire N__55549;
    wire N__55546;
    wire N__55543;
    wire N__55540;
    wire N__55537;
    wire N__55534;
    wire N__55531;
    wire N__55528;
    wire N__55525;
    wire N__55522;
    wire N__55519;
    wire N__55516;
    wire N__55515;
    wire N__55512;
    wire N__55509;
    wire N__55508;
    wire N__55507;
    wire N__55506;
    wire N__55501;
    wire N__55496;
    wire N__55495;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55483;
    wire N__55476;
    wire N__55471;
    wire N__55470;
    wire N__55469;
    wire N__55466;
    wire N__55463;
    wire N__55460;
    wire N__55457;
    wire N__55454;
    wire N__55451;
    wire N__55448;
    wire N__55447;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55426;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55414;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55392;
    wire N__55389;
    wire N__55386;
    wire N__55383;
    wire N__55382;
    wire N__55377;
    wire N__55374;
    wire N__55369;
    wire N__55366;
    wire N__55363;
    wire N__55362;
    wire N__55359;
    wire N__55356;
    wire N__55353;
    wire N__55352;
    wire N__55349;
    wire N__55346;
    wire N__55343;
    wire N__55336;
    wire N__55333;
    wire N__55330;
    wire N__55329;
    wire N__55326;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55316;
    wire N__55309;
    wire N__55306;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55296;
    wire N__55295;
    wire N__55292;
    wire N__55289;
    wire N__55286;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55272;
    wire N__55269;
    wire N__55268;
    wire N__55265;
    wire N__55262;
    wire N__55259;
    wire N__55252;
    wire N__55249;
    wire N__55248;
    wire N__55247;
    wire N__55246;
    wire N__55243;
    wire N__55240;
    wire N__55237;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55230;
    wire N__55229;
    wire N__55228;
    wire N__55227;
    wire N__55226;
    wire N__55225;
    wire N__55224;
    wire N__55223;
    wire N__55222;
    wire N__55221;
    wire N__55220;
    wire N__55219;
    wire N__55218;
    wire N__55217;
    wire N__55216;
    wire N__55215;
    wire N__55214;
    wire N__55213;
    wire N__55212;
    wire N__55211;
    wire N__55210;
    wire N__55209;
    wire N__55202;
    wire N__55193;
    wire N__55192;
    wire N__55191;
    wire N__55190;
    wire N__55189;
    wire N__55188;
    wire N__55187;
    wire N__55186;
    wire N__55185;
    wire N__55180;
    wire N__55175;
    wire N__55174;
    wire N__55173;
    wire N__55172;
    wire N__55169;
    wire N__55168;
    wire N__55167;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55163;
    wire N__55162;
    wire N__55161;
    wire N__55156;
    wire N__55153;
    wire N__55146;
    wire N__55145;
    wire N__55142;
    wire N__55141;
    wire N__55140;
    wire N__55137;
    wire N__55136;
    wire N__55135;
    wire N__55134;
    wire N__55133;
    wire N__55132;
    wire N__55131;
    wire N__55130;
    wire N__55129;
    wire N__55128;
    wire N__55127;
    wire N__55126;
    wire N__55125;
    wire N__55124;
    wire N__55123;
    wire N__55122;
    wire N__55121;
    wire N__55118;
    wire N__55117;
    wire N__55114;
    wire N__55113;
    wire N__55110;
    wire N__55109;
    wire N__55106;
    wire N__55103;
    wire N__55102;
    wire N__55099;
    wire N__55098;
    wire N__55095;
    wire N__55094;
    wire N__55091;
    wire N__55090;
    wire N__55089;
    wire N__55088;
    wire N__55087;
    wire N__55086;
    wire N__55085;
    wire N__55084;
    wire N__55083;
    wire N__55082;
    wire N__55081;
    wire N__55080;
    wire N__55079;
    wire N__55078;
    wire N__55077;
    wire N__55076;
    wire N__55073;
    wire N__55072;
    wire N__55071;
    wire N__55070;
    wire N__55069;
    wire N__55068;
    wire N__55067;
    wire N__55066;
    wire N__55065;
    wire N__55064;
    wire N__55063;
    wire N__55062;
    wire N__55061;
    wire N__55060;
    wire N__55057;
    wire N__55054;
    wire N__55047;
    wire N__55044;
    wire N__55041;
    wire N__55038;
    wire N__55035;
    wire N__55034;
    wire N__55031;
    wire N__55026;
    wire N__55019;
    wire N__55010;
    wire N__55001;
    wire N__54998;
    wire N__54997;
    wire N__54996;
    wire N__54995;
    wire N__54994;
    wire N__54993;
    wire N__54992;
    wire N__54991;
    wire N__54990;
    wire N__54989;
    wire N__54988;
    wire N__54987;
    wire N__54986;
    wire N__54985;
    wire N__54984;
    wire N__54983;
    wire N__54982;
    wire N__54981;
    wire N__54980;
    wire N__54979;
    wire N__54978;
    wire N__54977;
    wire N__54976;
    wire N__54975;
    wire N__54968;
    wire N__54959;
    wire N__54952;
    wire N__54951;
    wire N__54950;
    wire N__54949;
    wire N__54948;
    wire N__54947;
    wire N__54946;
    wire N__54945;
    wire N__54942;
    wire N__54941;
    wire N__54940;
    wire N__54939;
    wire N__54938;
    wire N__54937;
    wire N__54936;
    wire N__54935;
    wire N__54934;
    wire N__54931;
    wire N__54928;
    wire N__54927;
    wire N__54926;
    wire N__54925;
    wire N__54924;
    wire N__54923;
    wire N__54922;
    wire N__54921;
    wire N__54920;
    wire N__54917;
    wire N__54914;
    wire N__54911;
    wire N__54908;
    wire N__54905;
    wire N__54902;
    wire N__54899;
    wire N__54896;
    wire N__54893;
    wire N__54890;
    wire N__54889;
    wire N__54888;
    wire N__54887;
    wire N__54886;
    wire N__54885;
    wire N__54884;
    wire N__54883;
    wire N__54882;
    wire N__54881;
    wire N__54880;
    wire N__54879;
    wire N__54878;
    wire N__54877;
    wire N__54876;
    wire N__54875;
    wire N__54874;
    wire N__54873;
    wire N__54872;
    wire N__54871;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54867;
    wire N__54866;
    wire N__54865;
    wire N__54848;
    wire N__54831;
    wire N__54828;
    wire N__54827;
    wire N__54824;
    wire N__54823;
    wire N__54820;
    wire N__54819;
    wire N__54816;
    wire N__54815;
    wire N__54812;
    wire N__54809;
    wire N__54806;
    wire N__54803;
    wire N__54800;
    wire N__54797;
    wire N__54794;
    wire N__54791;
    wire N__54788;
    wire N__54785;
    wire N__54784;
    wire N__54779;
    wire N__54774;
    wire N__54773;
    wire N__54772;
    wire N__54771;
    wire N__54770;
    wire N__54769;
    wire N__54768;
    wire N__54767;
    wire N__54762;
    wire N__54759;
    wire N__54756;
    wire N__54749;
    wire N__54748;
    wire N__54745;
    wire N__54744;
    wire N__54743;
    wire N__54742;
    wire N__54741;
    wire N__54740;
    wire N__54739;
    wire N__54738;
    wire N__54735;
    wire N__54734;
    wire N__54733;
    wire N__54732;
    wire N__54731;
    wire N__54730;
    wire N__54729;
    wire N__54728;
    wire N__54727;
    wire N__54724;
    wire N__54717;
    wire N__54712;
    wire N__54703;
    wire N__54702;
    wire N__54701;
    wire N__54700;
    wire N__54699;
    wire N__54694;
    wire N__54689;
    wire N__54686;
    wire N__54683;
    wire N__54680;
    wire N__54679;
    wire N__54678;
    wire N__54677;
    wire N__54676;
    wire N__54673;
    wire N__54670;
    wire N__54669;
    wire N__54668;
    wire N__54665;
    wire N__54662;
    wire N__54659;
    wire N__54656;
    wire N__54653;
    wire N__54650;
    wire N__54649;
    wire N__54646;
    wire N__54643;
    wire N__54640;
    wire N__54637;
    wire N__54634;
    wire N__54631;
    wire N__54628;
    wire N__54625;
    wire N__54622;
    wire N__54621;
    wire N__54620;
    wire N__54619;
    wire N__54618;
    wire N__54617;
    wire N__54616;
    wire N__54615;
    wire N__54614;
    wire N__54613;
    wire N__54612;
    wire N__54611;
    wire N__54610;
    wire N__54609;
    wire N__54606;
    wire N__54605;
    wire N__54604;
    wire N__54603;
    wire N__54600;
    wire N__54599;
    wire N__54598;
    wire N__54597;
    wire N__54596;
    wire N__54595;
    wire N__54594;
    wire N__54593;
    wire N__54590;
    wire N__54589;
    wire N__54586;
    wire N__54585;
    wire N__54584;
    wire N__54583;
    wire N__54582;
    wire N__54581;
    wire N__54580;
    wire N__54573;
    wire N__54570;
    wire N__54567;
    wire N__54560;
    wire N__54549;
    wire N__54546;
    wire N__54539;
    wire N__54536;
    wire N__54535;
    wire N__54532;
    wire N__54531;
    wire N__54522;
    wire N__54521;
    wire N__54520;
    wire N__54519;
    wire N__54518;
    wire N__54517;
    wire N__54514;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54506;
    wire N__54505;
    wire N__54502;
    wire N__54501;
    wire N__54498;
    wire N__54495;
    wire N__54488;
    wire N__54479;
    wire N__54472;
    wire N__54471;
    wire N__54468;
    wire N__54465;
    wire N__54462;
    wire N__54459;
    wire N__54456;
    wire N__54453;
    wire N__54450;
    wire N__54447;
    wire N__54444;
    wire N__54441;
    wire N__54438;
    wire N__54435;
    wire N__54432;
    wire N__54431;
    wire N__54428;
    wire N__54425;
    wire N__54422;
    wire N__54419;
    wire N__54416;
    wire N__54413;
    wire N__54410;
    wire N__54407;
    wire N__54404;
    wire N__54403;
    wire N__54400;
    wire N__54397;
    wire N__54394;
    wire N__54389;
    wire N__54374;
    wire N__54367;
    wire N__54358;
    wire N__54347;
    wire N__54346;
    wire N__54345;
    wire N__54344;
    wire N__54343;
    wire N__54342;
    wire N__54341;
    wire N__54340;
    wire N__54339;
    wire N__54338;
    wire N__54337;
    wire N__54336;
    wire N__54331;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54321;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54308;
    wire N__54299;
    wire N__54292;
    wire N__54287;
    wire N__54284;
    wire N__54277;
    wire N__54272;
    wire N__54267;
    wire N__54266;
    wire N__54263;
    wire N__54260;
    wire N__54257;
    wire N__54256;
    wire N__54255;
    wire N__54254;
    wire N__54253;
    wire N__54252;
    wire N__54251;
    wire N__54250;
    wire N__54249;
    wire N__54248;
    wire N__54245;
    wire N__54242;
    wire N__54241;
    wire N__54240;
    wire N__54235;
    wire N__54230;
    wire N__54227;
    wire N__54220;
    wire N__54213;
    wire N__54204;
    wire N__54201;
    wire N__54198;
    wire N__54191;
    wire N__54186;
    wire N__54183;
    wire N__54172;
    wire N__54163;
    wire N__54154;
    wire N__54143;
    wire N__54134;
    wire N__54131;
    wire N__54124;
    wire N__54119;
    wire N__54116;
    wire N__54115;
    wire N__54112;
    wire N__54109;
    wire N__54106;
    wire N__54103;
    wire N__54100;
    wire N__54095;
    wire N__54090;
    wire N__54085;
    wire N__54084;
    wire N__54083;
    wire N__54082;
    wire N__54079;
    wire N__54078;
    wire N__54077;
    wire N__54070;
    wire N__54063;
    wire N__54060;
    wire N__54059;
    wire N__54058;
    wire N__54057;
    wire N__54042;
    wire N__54039;
    wire N__54034;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54018;
    wire N__54013;
    wire N__53998;
    wire N__53993;
    wire N__53992;
    wire N__53991;
    wire N__53990;
    wire N__53983;
    wire N__53974;
    wire N__53965;
    wire N__53958;
    wire N__53947;
    wire N__53938;
    wire N__53929;
    wire N__53920;
    wire N__53909;
    wire N__53906;
    wire N__53899;
    wire N__53892;
    wire N__53891;
    wire N__53890;
    wire N__53887;
    wire N__53884;
    wire N__53881;
    wire N__53878;
    wire N__53877;
    wire N__53872;
    wire N__53871;
    wire N__53870;
    wire N__53869;
    wire N__53866;
    wire N__53865;
    wire N__53862;
    wire N__53861;
    wire N__53860;
    wire N__53859;
    wire N__53858;
    wire N__53855;
    wire N__53852;
    wire N__53845;
    wire N__53842;
    wire N__53841;
    wire N__53840;
    wire N__53839;
    wire N__53838;
    wire N__53837;
    wire N__53836;
    wire N__53835;
    wire N__53834;
    wire N__53833;
    wire N__53832;
    wire N__53831;
    wire N__53830;
    wire N__53829;
    wire N__53828;
    wire N__53827;
    wire N__53822;
    wire N__53811;
    wire N__53808;
    wire N__53805;
    wire N__53796;
    wire N__53793;
    wire N__53792;
    wire N__53791;
    wire N__53790;
    wire N__53789;
    wire N__53786;
    wire N__53783;
    wire N__53780;
    wire N__53777;
    wire N__53774;
    wire N__53773;
    wire N__53770;
    wire N__53769;
    wire N__53768;
    wire N__53767;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53755;
    wire N__53742;
    wire N__53737;
    wire N__53736;
    wire N__53719;
    wire N__53714;
    wire N__53711;
    wire N__53702;
    wire N__53697;
    wire N__53690;
    wire N__53687;
    wire N__53682;
    wire N__53677;
    wire N__53676;
    wire N__53673;
    wire N__53672;
    wire N__53669;
    wire N__53668;
    wire N__53667;
    wire N__53666;
    wire N__53665;
    wire N__53664;
    wire N__53663;
    wire N__53662;
    wire N__53659;
    wire N__53654;
    wire N__53647;
    wire N__53630;
    wire N__53625;
    wire N__53622;
    wire N__53621;
    wire N__53620;
    wire N__53617;
    wire N__53616;
    wire N__53615;
    wire N__53612;
    wire N__53611;
    wire N__53608;
    wire N__53593;
    wire N__53584;
    wire N__53581;
    wire N__53570;
    wire N__53569;
    wire N__53566;
    wire N__53565;
    wire N__53564;
    wire N__53563;
    wire N__53562;
    wire N__53561;
    wire N__53560;
    wire N__53557;
    wire N__53554;
    wire N__53551;
    wire N__53550;
    wire N__53547;
    wire N__53536;
    wire N__53529;
    wire N__53524;
    wire N__53523;
    wire N__53514;
    wire N__53511;
    wire N__53510;
    wire N__53507;
    wire N__53504;
    wire N__53501;
    wire N__53500;
    wire N__53497;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53489;
    wire N__53486;
    wire N__53485;
    wire N__53484;
    wire N__53483;
    wire N__53482;
    wire N__53479;
    wire N__53472;
    wire N__53461;
    wire N__53458;
    wire N__53451;
    wire N__53444;
    wire N__53437;
    wire N__53426;
    wire N__53419;
    wire N__53418;
    wire N__53417;
    wire N__53416;
    wire N__53415;
    wire N__53408;
    wire N__53405;
    wire N__53400;
    wire N__53395;
    wire N__53388;
    wire N__53383;
    wire N__53374;
    wire N__53373;
    wire N__53370;
    wire N__53367;
    wire N__53366;
    wire N__53363;
    wire N__53362;
    wire N__53361;
    wire N__53360;
    wire N__53359;
    wire N__53358;
    wire N__53357;
    wire N__53356;
    wire N__53353;
    wire N__53352;
    wire N__53351;
    wire N__53350;
    wire N__53349;
    wire N__53348;
    wire N__53347;
    wire N__53344;
    wire N__53341;
    wire N__53340;
    wire N__53337;
    wire N__53330;
    wire N__53325;
    wire N__53318;
    wire N__53307;
    wire N__53296;
    wire N__53293;
    wire N__53284;
    wire N__53277;
    wire N__53274;
    wire N__53265;
    wire N__53258;
    wire N__53255;
    wire N__53252;
    wire N__53243;
    wire N__53232;
    wire N__53225;
    wire N__53222;
    wire N__53215;
    wire N__53210;
    wire N__53195;
    wire N__53192;
    wire N__53185;
    wire N__53180;
    wire N__53179;
    wire N__53178;
    wire N__53177;
    wire N__53172;
    wire N__53165;
    wire N__53154;
    wire N__53151;
    wire N__53144;
    wire N__53137;
    wire N__53126;
    wire N__53125;
    wire N__53124;
    wire N__53121;
    wire N__53118;
    wire N__53109;
    wire N__53108;
    wire N__53105;
    wire N__53098;
    wire N__53093;
    wire N__53088;
    wire N__53083;
    wire N__53066;
    wire N__53065;
    wire N__53064;
    wire N__53063;
    wire N__53054;
    wire N__53051;
    wire N__53044;
    wire N__53029;
    wire N__53020;
    wire N__53017;
    wire N__53016;
    wire N__53015;
    wire N__53014;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53008;
    wire N__53007;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52991;
    wire N__52986;
    wire N__52985;
    wire N__52982;
    wire N__52975;
    wire N__52968;
    wire N__52961;
    wire N__52950;
    wire N__52939;
    wire N__52934;
    wire N__52921;
    wire N__52918;
    wire N__52917;
    wire N__52914;
    wire N__52913;
    wire N__52910;
    wire N__52907;
    wire N__52904;
    wire N__52897;
    wire N__52896;
    wire N__52893;
    wire N__52890;
    wire N__52887;
    wire N__52884;
    wire N__52883;
    wire N__52882;
    wire N__52881;
    wire N__52876;
    wire N__52873;
    wire N__52870;
    wire N__52869;
    wire N__52866;
    wire N__52865;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52848;
    wire N__52845;
    wire N__52840;
    wire N__52835;
    wire N__52828;
    wire N__52827;
    wire N__52824;
    wire N__52823;
    wire N__52820;
    wire N__52817;
    wire N__52814;
    wire N__52811;
    wire N__52806;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52792;
    wire N__52789;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52776;
    wire N__52771;
    wire N__52770;
    wire N__52767;
    wire N__52764;
    wire N__52763;
    wire N__52760;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52748;
    wire N__52745;
    wire N__52742;
    wire N__52737;
    wire N__52732;
    wire N__52731;
    wire N__52728;
    wire N__52725;
    wire N__52722;
    wire N__52719;
    wire N__52714;
    wire N__52711;
    wire N__52708;
    wire N__52705;
    wire N__52702;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52694;
    wire N__52691;
    wire N__52688;
    wire N__52685;
    wire N__52678;
    wire N__52675;
    wire N__52674;
    wire N__52671;
    wire N__52670;
    wire N__52667;
    wire N__52664;
    wire N__52661;
    wire N__52654;
    wire N__52651;
    wire N__52650;
    wire N__52647;
    wire N__52644;
    wire N__52641;
    wire N__52640;
    wire N__52637;
    wire N__52634;
    wire N__52631;
    wire N__52624;
    wire N__52621;
    wire N__52618;
    wire N__52617;
    wire N__52616;
    wire N__52613;
    wire N__52610;
    wire N__52607;
    wire N__52604;
    wire N__52601;
    wire N__52594;
    wire N__52591;
    wire N__52590;
    wire N__52587;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52574;
    wire N__52571;
    wire N__52568;
    wire N__52561;
    wire N__52558;
    wire N__52555;
    wire N__52554;
    wire N__52551;
    wire N__52550;
    wire N__52547;
    wire N__52544;
    wire N__52541;
    wire N__52534;
    wire N__52531;
    wire N__52530;
    wire N__52527;
    wire N__52526;
    wire N__52523;
    wire N__52520;
    wire N__52517;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52494;
    wire N__52493;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52470;
    wire N__52467;
    wire N__52466;
    wire N__52463;
    wire N__52460;
    wire N__52457;
    wire N__52450;
    wire N__52447;
    wire N__52444;
    wire N__52443;
    wire N__52440;
    wire N__52437;
    wire N__52434;
    wire N__52433;
    wire N__52430;
    wire N__52427;
    wire N__52424;
    wire N__52417;
    wire N__52414;
    wire N__52411;
    wire N__52410;
    wire N__52407;
    wire N__52406;
    wire N__52403;
    wire N__52400;
    wire N__52397;
    wire N__52390;
    wire N__52387;
    wire N__52386;
    wire N__52383;
    wire N__52380;
    wire N__52377;
    wire N__52376;
    wire N__52373;
    wire N__52370;
    wire N__52367;
    wire N__52360;
    wire N__52357;
    wire N__52356;
    wire N__52353;
    wire N__52352;
    wire N__52349;
    wire N__52346;
    wire N__52343;
    wire N__52336;
    wire N__52333;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52325;
    wire N__52322;
    wire N__52319;
    wire N__52316;
    wire N__52309;
    wire N__52306;
    wire N__52305;
    wire N__52302;
    wire N__52301;
    wire N__52298;
    wire N__52295;
    wire N__52292;
    wire N__52285;
    wire N__52282;
    wire N__52281;
    wire N__52280;
    wire N__52277;
    wire N__52274;
    wire N__52271;
    wire N__52268;
    wire N__52265;
    wire N__52262;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52248;
    wire N__52245;
    wire N__52244;
    wire N__52241;
    wire N__52238;
    wire N__52235;
    wire N__52228;
    wire N__52225;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52205;
    wire N__52202;
    wire N__52199;
    wire N__52196;
    wire N__52189;
    wire N__52186;
    wire N__52183;
    wire N__52180;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52167;
    wire N__52164;
    wire N__52161;
    wire N__52158;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52141;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52133;
    wire N__52130;
    wire N__52127;
    wire N__52124;
    wire N__52119;
    wire N__52114;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52092;
    wire N__52089;
    wire N__52086;
    wire N__52083;
    wire N__52078;
    wire N__52077;
    wire N__52074;
    wire N__52071;
    wire N__52068;
    wire N__52063;
    wire N__52060;
    wire N__52057;
    wire N__52054;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52041;
    wire N__52040;
    wire N__52037;
    wire N__52032;
    wire N__52029;
    wire N__52026;
    wire N__52023;
    wire N__52020;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51997;
    wire N__51996;
    wire N__51993;
    wire N__51992;
    wire N__51989;
    wire N__51986;
    wire N__51983;
    wire N__51980;
    wire N__51975;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51942;
    wire N__51937;
    wire N__51934;
    wire N__51931;
    wire N__51930;
    wire N__51927;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51913;
    wire N__51910;
    wire N__51909;
    wire N__51906;
    wire N__51903;
    wire N__51900;
    wire N__51897;
    wire N__51894;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51880;
    wire N__51879;
    wire N__51876;
    wire N__51875;
    wire N__51872;
    wire N__51869;
    wire N__51866;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51843;
    wire N__51842;
    wire N__51839;
    wire N__51836;
    wire N__51833;
    wire N__51826;
    wire N__51823;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51808;
    wire N__51805;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51792;
    wire N__51789;
    wire N__51786;
    wire N__51783;
    wire N__51780;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51750;
    wire N__51749;
    wire N__51746;
    wire N__51743;
    wire N__51740;
    wire N__51735;
    wire N__51730;
    wire N__51727;
    wire N__51724;
    wire N__51721;
    wire N__51718;
    wire N__51715;
    wire N__51712;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51688;
    wire N__51685;
    wire N__51682;
    wire N__51679;
    wire N__51676;
    wire N__51673;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51663;
    wire N__51660;
    wire N__51657;
    wire N__51654;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51632;
    wire N__51629;
    wire N__51626;
    wire N__51623;
    wire N__51618;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51588;
    wire N__51585;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51555;
    wire N__51552;
    wire N__51549;
    wire N__51548;
    wire N__51545;
    wire N__51542;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51530;
    wire N__51523;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51498;
    wire N__51497;
    wire N__51494;
    wire N__51491;
    wire N__51488;
    wire N__51485;
    wire N__51482;
    wire N__51479;
    wire N__51476;
    wire N__51473;
    wire N__51466;
    wire N__51463;
    wire N__51460;
    wire N__51457;
    wire N__51454;
    wire N__51451;
    wire N__51448;
    wire N__51445;
    wire N__51444;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51434;
    wire N__51431;
    wire N__51428;
    wire N__51425;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51395;
    wire N__51392;
    wire N__51389;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51372;
    wire N__51367;
    wire N__51364;
    wire N__51361;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51348;
    wire N__51345;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51333;
    wire N__51330;
    wire N__51325;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51313;
    wire N__51310;
    wire N__51309;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51297;
    wire N__51294;
    wire N__51289;
    wire N__51286;
    wire N__51283;
    wire N__51280;
    wire N__51277;
    wire N__51274;
    wire N__51273;
    wire N__51272;
    wire N__51269;
    wire N__51266;
    wire N__51263;
    wire N__51260;
    wire N__51257;
    wire N__51254;
    wire N__51251;
    wire N__51248;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51222;
    wire N__51219;
    wire N__51216;
    wire N__51213;
    wire N__51212;
    wire N__51207;
    wire N__51204;
    wire N__51199;
    wire N__51196;
    wire N__51193;
    wire N__51190;
    wire N__51187;
    wire N__51184;
    wire N__51181;
    wire N__51180;
    wire N__51177;
    wire N__51176;
    wire N__51173;
    wire N__51170;
    wire N__51167;
    wire N__51164;
    wire N__51159;
    wire N__51156;
    wire N__51153;
    wire N__51150;
    wire N__51147;
    wire N__51144;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51127;
    wire N__51124;
    wire N__51121;
    wire N__51118;
    wire N__51117;
    wire N__51114;
    wire N__51111;
    wire N__51110;
    wire N__51107;
    wire N__51102;
    wire N__51099;
    wire N__51094;
    wire N__51091;
    wire N__51088;
    wire N__51085;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51073;
    wire N__51070;
    wire N__51069;
    wire N__51068;
    wire N__51065;
    wire N__51062;
    wire N__51059;
    wire N__51056;
    wire N__51053;
    wire N__51050;
    wire N__51047;
    wire N__51040;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51028;
    wire N__51025;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51013;
    wire N__51012;
    wire N__51011;
    wire N__51008;
    wire N__51003;
    wire N__50998;
    wire N__50995;
    wire N__50992;
    wire N__50989;
    wire N__50986;
    wire N__50983;
    wire N__50982;
    wire N__50979;
    wire N__50978;
    wire N__50975;
    wire N__50972;
    wire N__50969;
    wire N__50966;
    wire N__50963;
    wire N__50960;
    wire N__50953;
    wire N__50950;
    wire N__50947;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50935;
    wire N__50932;
    wire N__50929;
    wire N__50928;
    wire N__50925;
    wire N__50924;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50906;
    wire N__50903;
    wire N__50896;
    wire N__50893;
    wire N__50890;
    wire N__50887;
    wire N__50884;
    wire N__50881;
    wire N__50878;
    wire N__50877;
    wire N__50874;
    wire N__50871;
    wire N__50868;
    wire N__50865;
    wire N__50862;
    wire N__50859;
    wire N__50856;
    wire N__50855;
    wire N__50852;
    wire N__50849;
    wire N__50846;
    wire N__50839;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50827;
    wire N__50824;
    wire N__50821;
    wire N__50820;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50803;
    wire N__50800;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50788;
    wire N__50785;
    wire N__50782;
    wire N__50779;
    wire N__50776;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50764;
    wire N__50761;
    wire N__50760;
    wire N__50757;
    wire N__50754;
    wire N__50749;
    wire N__50746;
    wire N__50745;
    wire N__50742;
    wire N__50739;
    wire N__50734;
    wire N__50731;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50719;
    wire N__50716;
    wire N__50715;
    wire N__50712;
    wire N__50709;
    wire N__50706;
    wire N__50701;
    wire N__50698;
    wire N__50697;
    wire N__50694;
    wire N__50691;
    wire N__50688;
    wire N__50683;
    wire N__50680;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50668;
    wire N__50665;
    wire N__50662;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50650;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50638;
    wire N__50635;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50620;
    wire N__50617;
    wire N__50616;
    wire N__50613;
    wire N__50610;
    wire N__50605;
    wire N__50602;
    wire N__50601;
    wire N__50598;
    wire N__50595;
    wire N__50590;
    wire N__50587;
    wire N__50586;
    wire N__50583;
    wire N__50580;
    wire N__50575;
    wire N__50572;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50557;
    wire N__50554;
    wire N__50551;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50539;
    wire N__50536;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50524;
    wire N__50521;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50509;
    wire N__50506;
    wire N__50503;
    wire N__50500;
    wire N__50497;
    wire N__50494;
    wire N__50493;
    wire N__50488;
    wire N__50485;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50473;
    wire N__50470;
    wire N__50469;
    wire N__50466;
    wire N__50465;
    wire N__50462;
    wire N__50457;
    wire N__50452;
    wire N__50449;
    wire N__50448;
    wire N__50447;
    wire N__50440;
    wire N__50437;
    wire N__50436;
    wire N__50433;
    wire N__50432;
    wire N__50431;
    wire N__50428;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50416;
    wire N__50411;
    wire N__50408;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50393;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50377;
    wire N__50376;
    wire N__50373;
    wire N__50372;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50347;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50334;
    wire N__50333;
    wire N__50330;
    wire N__50325;
    wire N__50320;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50311;
    wire N__50310;
    wire N__50309;
    wire N__50306;
    wire N__50303;
    wire N__50298;
    wire N__50293;
    wire N__50290;
    wire N__50281;
    wire N__50278;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50265;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50238;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50220;
    wire N__50217;
    wire N__50214;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50173;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50155;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50113;
    wire N__50110;
    wire N__50109;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50105;
    wire N__50098;
    wire N__50097;
    wire N__50096;
    wire N__50095;
    wire N__50090;
    wire N__50087;
    wire N__50086;
    wire N__50085;
    wire N__50082;
    wire N__50079;
    wire N__50078;
    wire N__50077;
    wire N__50074;
    wire N__50073;
    wire N__50072;
    wire N__50071;
    wire N__50070;
    wire N__50069;
    wire N__50068;
    wire N__50065;
    wire N__50058;
    wire N__50053;
    wire N__50048;
    wire N__50045;
    wire N__50042;
    wire N__50033;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50025;
    wire N__50024;
    wire N__50023;
    wire N__50020;
    wire N__50019;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50013;
    wire N__50010;
    wire N__50005;
    wire N__50002;
    wire N__49999;
    wire N__49992;
    wire N__49989;
    wire N__49980;
    wire N__49977;
    wire N__49972;
    wire N__49963;
    wire N__49958;
    wire N__49955;
    wire N__49950;
    wire N__49933;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49925;
    wire N__49922;
    wire N__49919;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49907;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49876;
    wire N__49875;
    wire N__49872;
    wire N__49871;
    wire N__49868;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49860;
    wire N__49857;
    wire N__49856;
    wire N__49853;
    wire N__49852;
    wire N__49849;
    wire N__49848;
    wire N__49845;
    wire N__49844;
    wire N__49841;
    wire N__49840;
    wire N__49837;
    wire N__49836;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49812;
    wire N__49795;
    wire N__49778;
    wire N__49777;
    wire N__49774;
    wire N__49773;
    wire N__49770;
    wire N__49769;
    wire N__49766;
    wire N__49765;
    wire N__49758;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49702;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49689;
    wire N__49688;
    wire N__49685;
    wire N__49682;
    wire N__49679;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49656;
    wire N__49655;
    wire N__49652;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49640;
    wire N__49637;
    wire N__49634;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49618;
    wire N__49617;
    wire N__49616;
    wire N__49615;
    wire N__49614;
    wire N__49613;
    wire N__49612;
    wire N__49609;
    wire N__49608;
    wire N__49607;
    wire N__49606;
    wire N__49605;
    wire N__49604;
    wire N__49593;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49585;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49578;
    wire N__49577;
    wire N__49574;
    wire N__49573;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49554;
    wire N__49551;
    wire N__49546;
    wire N__49543;
    wire N__49530;
    wire N__49519;
    wire N__49506;
    wire N__49495;
    wire N__49490;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49463;
    wire N__49458;
    wire N__49455;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49424;
    wire N__49421;
    wire N__49418;
    wire N__49413;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49387;
    wire N__49386;
    wire N__49383;
    wire N__49380;
    wire N__49375;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49371;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49355;
    wire N__49354;
    wire N__49353;
    wire N__49350;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49340;
    wire N__49337;
    wire N__49336;
    wire N__49333;
    wire N__49330;
    wire N__49327;
    wire N__49326;
    wire N__49325;
    wire N__49324;
    wire N__49321;
    wire N__49320;
    wire N__49317;
    wire N__49316;
    wire N__49313;
    wire N__49312;
    wire N__49303;
    wire N__49302;
    wire N__49299;
    wire N__49298;
    wire N__49297;
    wire N__49296;
    wire N__49295;
    wire N__49294;
    wire N__49293;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49281;
    wire N__49274;
    wire N__49273;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49255;
    wire N__49252;
    wire N__49245;
    wire N__49232;
    wire N__49223;
    wire N__49220;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49174;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49162;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49118;
    wire N__49115;
    wire N__49112;
    wire N__49109;
    wire N__49106;
    wire N__49101;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49073;
    wire N__49070;
    wire N__49069;
    wire N__49066;
    wire N__49065;
    wire N__49064;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49044;
    wire N__49043;
    wire N__49042;
    wire N__49041;
    wire N__49040;
    wire N__49039;
    wire N__49036;
    wire N__49031;
    wire N__49026;
    wire N__49021;
    wire N__49020;
    wire N__49019;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48996;
    wire N__48995;
    wire N__48992;
    wire N__48989;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48981;
    wire N__48980;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48954;
    wire N__48945;
    wire N__48938;
    wire N__48929;
    wire N__48924;
    wire N__48907;
    wire N__48906;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48896;
    wire N__48893;
    wire N__48890;
    wire N__48887;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48865;
    wire N__48864;
    wire N__48863;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48851;
    wire N__48848;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48804;
    wire N__48801;
    wire N__48800;
    wire N__48795;
    wire N__48792;
    wire N__48789;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48759;
    wire N__48756;
    wire N__48753;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48741;
    wire N__48738;
    wire N__48735;
    wire N__48734;
    wire N__48729;
    wire N__48726;
    wire N__48723;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48672;
    wire N__48669;
    wire N__48666;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48639;
    wire N__48636;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48623;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48585;
    wire N__48582;
    wire N__48579;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48533;
    wire N__48528;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48494;
    wire N__48489;
    wire N__48486;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48429;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48410;
    wire N__48407;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48377;
    wire N__48374;
    wire N__48371;
    wire N__48368;
    wire N__48365;
    wire N__48362;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48336;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48324;
    wire N__48321;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48291;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48274;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48264;
    wire N__48263;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48224;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48210;
    wire N__48207;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48187;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48119;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48080;
    wire N__48077;
    wire N__48074;
    wire N__48071;
    wire N__48064;
    wire N__48061;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48042;
    wire N__48039;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48029;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48003;
    wire N__48000;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47983;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47973;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47952;
    wire N__47951;
    wire N__47948;
    wire N__47943;
    wire N__47940;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47918;
    wire N__47913;
    wire N__47910;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47890;
    wire N__47889;
    wire N__47886;
    wire N__47883;
    wire N__47882;
    wire N__47879;
    wire N__47874;
    wire N__47871;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47850;
    wire N__47847;
    wire N__47846;
    wire N__47843;
    wire N__47840;
    wire N__47837;
    wire N__47834;
    wire N__47831;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47815;
    wire N__47814;
    wire N__47811;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47796;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47726;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47689;
    wire N__47686;
    wire N__47683;
    wire N__47682;
    wire N__47679;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47630;
    wire N__47629;
    wire N__47628;
    wire N__47627;
    wire N__47626;
    wire N__47625;
    wire N__47620;
    wire N__47617;
    wire N__47616;
    wire N__47613;
    wire N__47608;
    wire N__47607;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47603;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47595;
    wire N__47594;
    wire N__47589;
    wire N__47586;
    wire N__47581;
    wire N__47578;
    wire N__47577;
    wire N__47574;
    wire N__47573;
    wire N__47572;
    wire N__47569;
    wire N__47568;
    wire N__47567;
    wire N__47564;
    wire N__47563;
    wire N__47562;
    wire N__47559;
    wire N__47558;
    wire N__47555;
    wire N__47554;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47523;
    wire N__47516;
    wire N__47511;
    wire N__47500;
    wire N__47495;
    wire N__47488;
    wire N__47473;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47434;
    wire N__47431;
    wire N__47430;
    wire N__47427;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47410;
    wire N__47407;
    wire N__47406;
    wire N__47403;
    wire N__47400;
    wire N__47397;
    wire N__47396;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47377;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47361;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47314;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47303;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47289;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47249;
    wire N__47244;
    wire N__47241;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47211;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47171;
    wire N__47166;
    wire N__47163;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47149;
    wire N__47148;
    wire N__47145;
    wire N__47142;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47103;
    wire N__47102;
    wire N__47099;
    wire N__47094;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47082;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47065;
    wire N__47062;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47029;
    wire N__47026;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46927;
    wire N__46926;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46913;
    wire N__46906;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46882;
    wire N__46877;
    wire N__46874;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46843;
    wire N__46842;
    wire N__46841;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46829;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46809;
    wire N__46804;
    wire N__46801;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46774;
    wire N__46771;
    wire N__46768;
    wire N__46767;
    wire N__46766;
    wire N__46763;
    wire N__46760;
    wire N__46757;
    wire N__46754;
    wire N__46747;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46696;
    wire N__46695;
    wire N__46690;
    wire N__46687;
    wire N__46684;
    wire N__46681;
    wire N__46678;
    wire N__46677;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46645;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46633;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46618;
    wire N__46615;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46560;
    wire N__46557;
    wire N__46554;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46521;
    wire N__46518;
    wire N__46515;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46174;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46144;
    wire N__46141;
    wire N__46138;
    wire N__46135;
    wire N__46134;
    wire N__46133;
    wire N__46130;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46107;
    wire N__46106;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46006;
    wire N__46003;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45970;
    wire N__45967;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45943;
    wire N__45940;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45919;
    wire N__45916;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45889;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45838;
    wire N__45837;
    wire N__45834;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45769;
    wire N__45766;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45758;
    wire N__45753;
    wire N__45750;
    wire N__45745;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45705;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45670;
    wire N__45669;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45654;
    wire N__45651;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45621;
    wire N__45618;
    wire N__45615;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45601;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45569;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45495;
    wire N__45492;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45423;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45413;
    wire N__45408;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45379;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45338;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45322;
    wire N__45319;
    wire N__45316;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45273;
    wire N__45270;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45252;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45225;
    wire N__45222;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45154;
    wire N__45151;
    wire N__45150;
    wire N__45147;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45117;
    wire N__45114;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45087;
    wire N__45084;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45035;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45012;
    wire N__45009;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44943;
    wire N__44940;
    wire N__44939;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44923;
    wire N__44920;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44912;
    wire N__44907;
    wire N__44904;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44892;
    wire N__44889;
    wire N__44888;
    wire N__44885;
    wire N__44882;
    wire N__44879;
    wire N__44876;
    wire N__44873;
    wire N__44870;
    wire N__44867;
    wire N__44864;
    wire N__44861;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44810;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44733;
    wire N__44732;
    wire N__44729;
    wire N__44726;
    wire N__44723;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44684;
    wire N__44681;
    wire N__44678;
    wire N__44675;
    wire N__44668;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44654;
    wire N__44651;
    wire N__44648;
    wire N__44645;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44629;
    wire N__44626;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44615;
    wire N__44610;
    wire N__44607;
    wire N__44602;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44557;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44545;
    wire N__44544;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44528;
    wire N__44523;
    wire N__44520;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44461;
    wire N__44460;
    wire N__44457;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44409;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44385;
    wire N__44382;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44287;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44275;
    wire N__44274;
    wire N__44271;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44256;
    wire N__44251;
    wire N__44250;
    wire N__44247;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44229;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44193;
    wire N__44190;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44177;
    wire N__44170;
    wire N__44167;
    wire N__44166;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44148;
    wire N__44143;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44115;
    wire N__44112;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44061;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44051;
    wire N__44046;
    wire N__44041;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44031;
    wire N__44030;
    wire N__44027;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44008;
    wire N__44005;
    wire N__44004;
    wire N__44001;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43974;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43950;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43647;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43620;
    wire N__43619;
    wire N__43616;
    wire N__43611;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43545;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43528;
    wire N__43527;
    wire N__43524;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43498;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43482;
    wire N__43479;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43380;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43341;
    wire N__43338;
    wire N__43337;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43302;
    wire N__43299;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43229;
    wire N__43224;
    wire N__43221;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43203;
    wire N__43200;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43167;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43131;
    wire N__43130;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43005;
    wire N__43004;
    wire N__43003;
    wire N__43002;
    wire N__43001;
    wire N__43000;
    wire N__42999;
    wire N__42998;
    wire N__42997;
    wire N__42996;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42990;
    wire N__42981;
    wire N__42980;
    wire N__42979;
    wire N__42976;
    wire N__42975;
    wire N__42972;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42964;
    wire N__42963;
    wire N__42962;
    wire N__42961;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42946;
    wire N__42945;
    wire N__42942;
    wire N__42941;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42920;
    wire N__42913;
    wire N__42906;
    wire N__42897;
    wire N__42888;
    wire N__42881;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42822;
    wire N__42819;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42792;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42765;
    wire N__42762;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42687;
    wire N__42684;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42595;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42532;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42524;
    wire N__42519;
    wire N__42516;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42474;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42448;
    wire N__42445;
    wire N__42444;
    wire N__42443;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42430;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42423;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42405;
    wire N__42404;
    wire N__42403;
    wire N__42402;
    wire N__42399;
    wire N__42398;
    wire N__42397;
    wire N__42396;
    wire N__42395;
    wire N__42392;
    wire N__42391;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42383;
    wire N__42382;
    wire N__42375;
    wire N__42368;
    wire N__42357;
    wire N__42346;
    wire N__42341;
    wire N__42336;
    wire N__42325;
    wire N__42310;
    wire N__42309;
    wire N__42306;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42288;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42232;
    wire N__42231;
    wire N__42228;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42207;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42173;
    wire N__42168;
    wire N__42165;
    wire N__42160;
    wire N__42157;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42131;
    wire N__42126;
    wire N__42123;
    wire N__42118;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42064;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41985;
    wire N__41982;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41962;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41951;
    wire N__41946;
    wire N__41943;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41856;
    wire N__41853;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41833;
    wire N__41832;
    wire N__41829;
    wire N__41828;
    wire N__41825;
    wire N__41820;
    wire N__41817;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41799;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41767;
    wire N__41764;
    wire N__41763;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41716;
    wire N__41713;
    wire N__41712;
    wire N__41711;
    wire N__41708;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41692;
    wire N__41691;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41674;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41657;
    wire N__41650;
    wire N__41647;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41593;
    wire N__41590;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41568;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41544;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41532;
    wire N__41531;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41519;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41479;
    wire N__41476;
    wire N__41475;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41429;
    wire N__41424;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41400;
    wire N__41399;
    wire N__41396;
    wire N__41391;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41373;
    wire N__41368;
    wire N__41365;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41343;
    wire N__41342;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41324;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41293;
    wire N__41292;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41280;
    wire N__41275;
    wire N__41272;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41235;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41202;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41190;
    wire N__41187;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41165;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41143;
    wire N__41142;
    wire N__41141;
    wire N__41140;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41132;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41124;
    wire N__41121;
    wire N__41116;
    wire N__41107;
    wire N__41104;
    wire N__41095;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41068;
    wire N__41067;
    wire N__41066;
    wire N__41061;
    wire N__41060;
    wire N__41059;
    wire N__41058;
    wire N__41057;
    wire N__41056;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41035;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41019;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40996;
    wire N__40993;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40974;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40893;
    wire N__40892;
    wire N__40889;
    wire N__40884;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40869;
    wire N__40868;
    wire N__40867;
    wire N__40864;
    wire N__40863;
    wire N__40860;
    wire N__40859;
    wire N__40856;
    wire N__40855;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40786;
    wire N__40783;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40768;
    wire N__40767;
    wire N__40766;
    wire N__40763;
    wire N__40758;
    wire N__40753;
    wire N__40750;
    wire N__40749;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40722;
    wire N__40719;
    wire N__40718;
    wire N__40715;
    wire N__40712;
    wire N__40709;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40534;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40522;
    wire N__40519;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40470;
    wire N__40467;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40366;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40341;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40216;
    wire N__40213;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40177;
    wire N__40176;
    wire N__40175;
    wire N__40170;
    wire N__40169;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40134;
    wire N__40131;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40096;
    wire N__40093;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40081;
    wire N__40078;
    wire N__40077;
    wire N__40074;
    wire N__40071;
    wire N__40066;
    wire N__40063;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40048;
    wire N__40045;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40005;
    wire N__40004;
    wire N__40001;
    wire N__39996;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39951;
    wire N__39948;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39849;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39822;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39564;
    wire N__39563;
    wire N__39562;
    wire N__39559;
    wire N__39558;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39548;
    wire N__39547;
    wire N__39546;
    wire N__39543;
    wire N__39542;
    wire N__39539;
    wire N__39536;
    wire N__39535;
    wire N__39534;
    wire N__39533;
    wire N__39532;
    wire N__39531;
    wire N__39530;
    wire N__39529;
    wire N__39528;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39497;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39487;
    wire N__39486;
    wire N__39485;
    wire N__39482;
    wire N__39481;
    wire N__39480;
    wire N__39477;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39471;
    wire N__39468;
    wire N__39467;
    wire N__39466;
    wire N__39465;
    wire N__39462;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39445;
    wire N__39444;
    wire N__39443;
    wire N__39442;
    wire N__39437;
    wire N__39434;
    wire N__39429;
    wire N__39422;
    wire N__39419;
    wire N__39408;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39391;
    wire N__39386;
    wire N__39379;
    wire N__39374;
    wire N__39367;
    wire N__39364;
    wire N__39349;
    wire N__39342;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39179;
    wire N__39174;
    wire N__39171;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39150;
    wire N__39149;
    wire N__39146;
    wire N__39145;
    wire N__39144;
    wire N__39143;
    wire N__39140;
    wire N__39139;
    wire N__39138;
    wire N__39135;
    wire N__39134;
    wire N__39133;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39119;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39105;
    wire N__39104;
    wire N__39099;
    wire N__39098;
    wire N__39097;
    wire N__39096;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39072;
    wire N__39071;
    wire N__39068;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39056;
    wire N__39051;
    wire N__39042;
    wire N__39037;
    wire N__39028;
    wire N__39013;
    wire N__39012;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38936;
    wire N__38935;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38931;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38909;
    wire N__38908;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38900;
    wire N__38899;
    wire N__38898;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38869;
    wire N__38868;
    wire N__38863;
    wire N__38862;
    wire N__38861;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38838;
    wire N__38835;
    wire N__38828;
    wire N__38825;
    wire N__38820;
    wire N__38807;
    wire N__38794;
    wire N__38791;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38776;
    wire N__38775;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38737;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38712;
    wire N__38707;
    wire N__38704;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38679;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38624;
    wire N__38619;
    wire N__38616;
    wire N__38611;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38586;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38550;
    wire N__38549;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38537;
    wire N__38532;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38487;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38469;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38442;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38394;
    wire N__38393;
    wire N__38390;
    wire N__38385;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38283;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38262;
    wire N__38261;
    wire N__38258;
    wire N__38257;
    wire N__38252;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38199;
    wire N__38198;
    wire N__38193;
    wire N__38192;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38172;
    wire N__38171;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38155;
    wire N__38154;
    wire N__38151;
    wire N__38150;
    wire N__38149;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38088;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38070;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38048;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37776;
    wire N__37773;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37758;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37713;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37690;
    wire N__37687;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37679;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37632;
    wire N__37629;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37603;
    wire N__37600;
    wire N__37599;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37581;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37516;
    wire N__37513;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37505;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37483;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37467;
    wire N__37464;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37426;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37296;
    wire N__37293;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37245;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37218;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37191;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37164;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37122;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37027;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36925;
    wire N__36918;
    wire N__36915;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36882;
    wire N__36879;
    wire N__36876;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36855;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36832;
    wire N__36831;
    wire N__36826;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36814;
    wire N__36813;
    wire N__36810;
    wire N__36805;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36793;
    wire N__36790;
    wire N__36789;
    wire N__36784;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36745;
    wire N__36744;
    wire N__36743;
    wire N__36740;
    wire N__36739;
    wire N__36734;
    wire N__36733;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36725;
    wire N__36722;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36716;
    wire N__36715;
    wire N__36712;
    wire N__36711;
    wire N__36708;
    wire N__36703;
    wire N__36700;
    wire N__36695;
    wire N__36684;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36629;
    wire N__36628;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36604;
    wire N__36601;
    wire N__36590;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36553;
    wire N__36550;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36542;
    wire N__36541;
    wire N__36540;
    wire N__36539;
    wire N__36538;
    wire N__36537;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36515;
    wire N__36512;
    wire N__36503;
    wire N__36490;
    wire N__36487;
    wire N__36486;
    wire N__36485;
    wire N__36484;
    wire N__36483;
    wire N__36482;
    wire N__36481;
    wire N__36480;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36476;
    wire N__36475;
    wire N__36474;
    wire N__36473;
    wire N__36472;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36406;
    wire N__36403;
    wire N__36388;
    wire N__36379;
    wire N__36376;
    wire N__36367;
    wire N__36362;
    wire N__36349;
    wire N__36342;
    wire N__36339;
    wire N__36332;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36261;
    wire N__36260;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36211;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36177;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36169;
    wire N__36168;
    wire N__36163;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36136;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36118;
    wire N__36113;
    wire N__36104;
    wire N__36097;
    wire N__36094;
    wire N__36089;
    wire N__36076;
    wire N__36073;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36049;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36032;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36015;
    wire N__36012;
    wire N__36007;
    wire N__35998;
    wire N__35995;
    wire N__35994;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35988;
    wire N__35987;
    wire N__35986;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35978;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35950;
    wire N__35941;
    wire N__35938;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35894;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35875;
    wire N__35874;
    wire N__35873;
    wire N__35872;
    wire N__35871;
    wire N__35870;
    wire N__35869;
    wire N__35868;
    wire N__35867;
    wire N__35864;
    wire N__35863;
    wire N__35862;
    wire N__35859;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35825;
    wire N__35812;
    wire N__35807;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35766;
    wire N__35765;
    wire N__35762;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35751;
    wire N__35748;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35734;
    wire N__35733;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35727;
    wire N__35726;
    wire N__35725;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35689;
    wire N__35680;
    wire N__35675;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35629;
    wire N__35628;
    wire N__35625;
    wire N__35624;
    wire N__35623;
    wire N__35622;
    wire N__35621;
    wire N__35620;
    wire N__35619;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35600;
    wire N__35599;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35585;
    wire N__35584;
    wire N__35581;
    wire N__35574;
    wire N__35571;
    wire N__35566;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35543;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35493;
    wire N__35492;
    wire N__35491;
    wire N__35488;
    wire N__35487;
    wire N__35486;
    wire N__35485;
    wire N__35484;
    wire N__35483;
    wire N__35482;
    wire N__35481;
    wire N__35480;
    wire N__35477;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35469;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35455;
    wire N__35446;
    wire N__35433;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35389;
    wire N__35388;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35382;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35361;
    wire N__35356;
    wire N__35353;
    wire N__35342;
    wire N__35331;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35286;
    wire N__35283;
    wire N__35282;
    wire N__35281;
    wire N__35280;
    wire N__35279;
    wire N__35276;
    wire N__35275;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35256;
    wire N__35251;
    wire N__35248;
    wire N__35247;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35215;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35106;
    wire N__35105;
    wire N__35104;
    wire N__35103;
    wire N__35102;
    wire N__35101;
    wire N__35098;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35085;
    wire N__35084;
    wire N__35081;
    wire N__35076;
    wire N__35075;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35054;
    wire N__35053;
    wire N__35052;
    wire N__35049;
    wire N__35048;
    wire N__35047;
    wire N__35046;
    wire N__35039;
    wire N__35034;
    wire N__35031;
    wire N__35026;
    wire N__35023;
    wire N__35018;
    wire N__35015;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__34997;
    wire N__34994;
    wire N__34989;
    wire N__34978;
    wire N__34975;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34939;
    wire N__34936;
    wire N__34935;
    wire N__34932;
    wire N__34931;
    wire N__34930;
    wire N__34929;
    wire N__34928;
    wire N__34927;
    wire N__34926;
    wire N__34925;
    wire N__34924;
    wire N__34921;
    wire N__34920;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34906;
    wire N__34905;
    wire N__34904;
    wire N__34901;
    wire N__34900;
    wire N__34897;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34891;
    wire N__34890;
    wire N__34885;
    wire N__34882;
    wire N__34877;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34861;
    wire N__34852;
    wire N__34847;
    wire N__34838;
    wire N__34835;
    wire N__34830;
    wire N__34823;
    wire N__34818;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34581;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34522;
    wire N__34519;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34497;
    wire N__34494;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34444;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34251;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34225;
    wire N__34224;
    wire N__34223;
    wire N__34220;
    wire N__34219;
    wire N__34216;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34206;
    wire N__34199;
    wire N__34192;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34174;
    wire N__34171;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34147;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34129;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34038;
    wire N__34035;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34018;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34004;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33985;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33969;
    wire N__33966;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33928;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33874;
    wire N__33873;
    wire N__33870;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33853;
    wire N__33850;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33771;
    wire N__33770;
    wire N__33767;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33738;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33712;
    wire N__33709;
    wire N__33708;
    wire N__33707;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33617;
    wire N__33612;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33573;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33558;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33522;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33462;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33411;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33393;
    wire N__33392;
    wire N__33389;
    wire N__33388;
    wire N__33383;
    wire N__33378;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33354;
    wire N__33351;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32799;
    wire N__32796;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32776;
    wire N__32775;
    wire N__32772;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32737;
    wire N__32734;
    wire N__32733;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32695;
    wire N__32694;
    wire N__32691;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32641;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32582;
    wire N__32577;
    wire N__32572;
    wire N__32569;
    wire N__32568;
    wire N__32565;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32475;
    wire N__32472;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32455;
    wire N__32452;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32433;
    wire N__32430;
    wire N__32425;
    wire N__32422;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32395;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32362;
    wire N__32359;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32343;
    wire N__32340;
    wire N__32335;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32302;
    wire N__32299;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32281;
    wire N__32278;
    wire N__32277;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32256;
    wire N__32253;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32209;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32161;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32149;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32079;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32022;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31974;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31734;
    wire N__31731;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31623;
    wire N__31620;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31548;
    wire N__31547;
    wire N__31544;
    wire N__31539;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31521;
    wire N__31518;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31503;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31437;
    wire N__31434;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31422;
    wire N__31419;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31396;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31362;
    wire N__31359;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31293;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31275;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31194;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31170;
    wire N__31169;
    wire N__31166;
    wire N__31161;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31033;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31019;
    wire N__31014;
    wire N__31011;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30976;
    wire N__30973;
    wire N__30972;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30784;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30682;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30670;
    wire N__30669;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30602;
    wire N__30597;
    wire N__30594;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30517;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30493;
    wire N__30492;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30453;
    wire N__30450;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30418;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30407;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30391;
    wire N__30390;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30318;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30276;
    wire N__30273;
    wire N__30272;
    wire N__30271;
    wire N__30268;
    wire N__30263;
    wire N__30260;
    wire N__30255;
    wire N__30250;
    wire N__30249;
    wire N__30246;
    wire N__30245;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30121;
    wire N__30120;
    wire N__30117;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30068;
    wire N__30065;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30043;
    wire N__30040;
    wire N__30037;
    wire N__30036;
    wire N__30035;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29976;
    wire N__29975;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29959;
    wire N__29956;
    wire N__29955;
    wire N__29952;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29932;
    wire N__29929;
    wire N__29928;
    wire N__29923;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29901;
    wire N__29898;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29880;
    wire N__29875;
    wire N__29872;
    wire N__29871;
    wire N__29866;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29705;
    wire N__29700;
    wire N__29697;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29677;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29665;
    wire N__29662;
    wire N__29661;
    wire N__29658;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29505;
    wire N__29502;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29425;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29406;
    wire N__29403;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29370;
    wire N__29367;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29322;
    wire N__29321;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29280;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29181;
    wire N__29178;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29102;
    wire N__29097;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29073;
    wire N__29070;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29058;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29001;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28789;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28758;
    wire N__28755;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28706;
    wire N__28703;
    wire N__28698;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28683;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28663;
    wire N__28660;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28633;
    wire N__28630;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28537;
    wire N__28536;
    wire N__28533;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28450;
    wire N__28447;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28390;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28366;
    wire N__28363;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28282;
    wire N__28279;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28267;
    wire N__28264;
    wire N__28263;
    wire N__28260;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28147;
    wire N__28144;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28120;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28098;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28024;
    wire N__28021;
    wire N__28020;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27994;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27945;
    wire N__27944;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27932;
    wire N__27925;
    wire N__27922;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27886;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27872;
    wire N__27867;
    wire N__27864;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27835;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27821;
    wire N__27816;
    wire N__27813;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27798;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27725;
    wire N__27720;
    wire N__27717;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27685;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27635;
    wire N__27630;
    wire N__27627;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27582;
    wire N__27579;
    wire N__27574;
    wire N__27571;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27563;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27414;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27325;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27310;
    wire N__27307;
    wire N__27306;
    wire N__27303;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27285;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27273;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27244;
    wire N__27241;
    wire N__27240;
    wire N__27237;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27164;
    wire N__27159;
    wire N__27156;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27132;
    wire N__27129;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27091;
    wire N__27088;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27057;
    wire N__27054;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26960;
    wire N__26955;
    wire N__26952;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26901;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26861;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26845;
    wire N__26842;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26773;
    wire N__26770;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26748;
    wire N__26743;
    wire N__26740;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26718;
    wire N__26713;
    wire N__26710;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26693;
    wire N__26688;
    wire N__26685;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26256;
    wire N__26253;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26220;
    wire N__26217;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26164;
    wire N__26161;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26133;
    wire N__26130;
    wire N__26125;
    wire N__26122;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26110;
    wire N__26109;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26092;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26079;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26019;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25938;
    wire N__25935;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25845;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25725;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25492;
    wire N__25489;
    wire N__25488;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25437;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25386;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25374;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25353;
    wire N__25352;
    wire N__25349;
    wire N__25344;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25245;
    wire N__25242;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25173;
    wire N__25170;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25134;
    wire N__25133;
    wire N__25130;
    wire N__25125;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25004;
    wire N__24999;
    wire N__24996;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24928;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24798;
    wire N__24795;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24729;
    wire N__24726;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24628;
    wire N__24625;
    wire N__24624;
    wire N__24621;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24561;
    wire N__24558;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24541;
    wire N__24538;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24530;
    wire N__24527;
    wire N__24522;
    wire N__24519;
    wire N__24514;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24499;
    wire N__24498;
    wire N__24495;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24378;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24330;
    wire N__24329;
    wire N__24326;
    wire N__24321;
    wire N__24316;
    wire N__24313;
    wire N__24312;
    wire N__24309;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24294;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24241;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24224;
    wire N__24219;
    wire N__24216;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24166;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24108;
    wire N__24105;
    wire N__24104;
    wire N__24101;
    wire N__24096;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23925;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23664;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23578;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23532;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23506;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23498;
    wire N__23493;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23452;
    wire N__23449;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23409;
    wire N__23408;
    wire N__23405;
    wire N__23400;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23388;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23373;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23253;
    wire N__23250;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23238;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23164;
    wire N__23161;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22980;
    wire N__22977;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22890;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22672;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22344;
    wire N__22339;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22331;
    wire N__22326;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22122;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22048;
    wire N__22045;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21986;
    wire N__21981;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21904;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21889;
    wire N__21886;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21871;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21841;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_17_0_;
    wire n12257;
    wire n12258;
    wire n12259;
    wire n12260;
    wire n12261;
    wire n12262;
    wire n12263;
    wire n12264;
    wire bfn_1_18_0_;
    wire n12265;
    wire n12266;
    wire n12267;
    wire n12268;
    wire n12269;
    wire n12270;
    wire n12271;
    wire n12272;
    wire bfn_1_19_0_;
    wire n12273;
    wire n12274;
    wire n12275;
    wire bfn_1_20_0_;
    wire n12239;
    wire n12240;
    wire n12241;
    wire n12242;
    wire n12243;
    wire n12244;
    wire n12245;
    wire n12246;
    wire bfn_1_21_0_;
    wire n12247;
    wire n12248;
    wire n12249;
    wire n12250;
    wire n12251;
    wire n12252;
    wire n12253;
    wire n12254;
    wire bfn_1_22_0_;
    wire n12255;
    wire n12256;
    wire bfn_1_23_0_;
    wire n12206;
    wire n12207;
    wire n12208;
    wire n12209;
    wire n12210;
    wire n12211;
    wire n12212;
    wire n12213;
    wire bfn_1_24_0_;
    wire n12214;
    wire n12215;
    wire n12216;
    wire n12217;
    wire n12218;
    wire n12219;
    wire n12220;
    wire n12221;
    wire bfn_1_25_0_;
    wire bfn_1_26_0_;
    wire n12177;
    wire n12178;
    wire n12179;
    wire n12180;
    wire n12181;
    wire n12182;
    wire n12183;
    wire n12184;
    wire bfn_1_27_0_;
    wire n12185;
    wire n12186;
    wire n12187;
    wire n12188;
    wire n12189;
    wire n12190;
    wire n1427_cascade_;
    wire n1430_cascade_;
    wire n11638;
    wire bfn_1_29_0_;
    wire \debounce.n12654 ;
    wire \debounce.n12655 ;
    wire \debounce.n12656 ;
    wire \debounce.n12657 ;
    wire \debounce.n12658 ;
    wire \debounce.n12659 ;
    wire \debounce.n12660 ;
    wire \debounce.n12661 ;
    wire bfn_1_30_0_;
    wire \debounce.n12662 ;
    wire bfn_1_31_0_;
    wire n12122;
    wire n12123;
    wire n12124;
    wire n12125;
    wire n12126;
    wire n12127;
    wire n12128;
    wire n12129;
    wire bfn_1_32_0_;
    wire n12130;
    wire \debounce.cnt_reg_3 ;
    wire \debounce.cnt_reg_9 ;
    wire \debounce.cnt_reg_5 ;
    wire \debounce.cnt_reg_8 ;
    wire \debounce.cnt_reg_1 ;
    wire \debounce.cnt_reg_2 ;
    wire \debounce.n14472_cascade_ ;
    wire n2095;
    wire n2094;
    wire n2101;
    wire n2200;
    wire n2133_cascade_;
    wire n2232_cascade_;
    wire n2331_cascade_;
    wire n2089;
    wire n2188;
    wire n2121_cascade_;
    wire n2220_cascade_;
    wire n2319_cascade_;
    wire n2097;
    wire n2049_cascade_;
    wire n2183;
    wire n2184;
    wire n2084;
    wire n2116;
    wire n2115;
    wire n2116_cascade_;
    wire n2148_cascade_;
    wire n2195;
    wire n2087;
    wire n2093;
    wire n2085;
    wire n2117;
    wire bfn_2_21_0_;
    wire n12222;
    wire n12223;
    wire n12224;
    wire n12225;
    wire n12226;
    wire n12227;
    wire n12228;
    wire n12229;
    wire bfn_2_22_0_;
    wire n12230;
    wire n12231;
    wire n12232;
    wire n12233;
    wire n12234;
    wire n12235;
    wire n12236;
    wire n12237;
    wire bfn_2_23_0_;
    wire n12238;
    wire n2016;
    wire n1888;
    wire n1985;
    wire n2017;
    wire n1700;
    wire n1699;
    wire n1731_cascade_;
    wire n1697;
    wire n1729_cascade_;
    wire n1701;
    wire n1733_cascade_;
    wire n1886;
    wire n1698;
    wire n1696;
    wire n1728_cascade_;
    wire n1695;
    wire n1694;
    wire n1689;
    wire n1630;
    wire n13986_cascade_;
    wire n1554_cascade_;
    wire n1629;
    wire n1631;
    wire bfn_2_27_0_;
    wire n12152;
    wire n12153;
    wire n12154;
    wire n12155;
    wire n12156;
    wire n12157;
    wire n12158;
    wire n12159;
    wire bfn_2_28_0_;
    wire n12160;
    wire n12161;
    wire n12162;
    wire n12163;
    wire n1491;
    wire n26_adj_678;
    wire bfn_2_29_0_;
    wire n25_adj_677;
    wire n12717;
    wire n24_adj_676;
    wire n12718;
    wire n23_adj_675;
    wire n12719;
    wire n22_adj_674;
    wire n12720;
    wire n21_adj_673;
    wire n12721;
    wire n20_adj_672;
    wire n12722;
    wire n19_adj_671;
    wire n12723;
    wire n12724;
    wire n18_adj_670;
    wire bfn_2_30_0_;
    wire n17_adj_669;
    wire n12725;
    wire n16_adj_668;
    wire n12726;
    wire n15_adj_667;
    wire n12727;
    wire n14_adj_666;
    wire n12728;
    wire n13_adj_665;
    wire n12729;
    wire n12_adj_664;
    wire n12730;
    wire n11_adj_663;
    wire n12731;
    wire n12732;
    wire n10_adj_662;
    wire bfn_2_31_0_;
    wire n9_adj_661;
    wire n12733;
    wire n8_adj_660;
    wire n12734;
    wire n7_adj_659;
    wire n12735;
    wire n6_adj_658;
    wire n12736;
    wire n12737;
    wire n12738;
    wire n12739;
    wire n12740;
    wire bfn_2_32_0_;
    wire n12741;
    wire \debounce.cnt_reg_4 ;
    wire \debounce.cnt_reg_6 ;
    wire \debounce.cnt_reg_0 ;
    wire \debounce.cnt_reg_7 ;
    wire \debounce.n13 ;
    wire bfn_3_17_0_;
    wire n12296;
    wire n12297;
    wire n2398;
    wire n12298;
    wire n12299;
    wire n12300;
    wire n12301;
    wire n12302;
    wire n12303;
    wire bfn_3_18_0_;
    wire n12304;
    wire n12305;
    wire n12306;
    wire n12307;
    wire n12308;
    wire n12309;
    wire n2386;
    wire n12310;
    wire n12311;
    wire bfn_3_19_0_;
    wire n12312;
    wire n12313;
    wire n12314;
    wire n12315;
    wire n12316;
    wire n2098;
    wire n2392;
    wire n2096;
    wire n2197;
    wire n1996;
    wire n2196;
    wire n2201;
    wire n14160;
    wire n2186;
    wire n2028;
    wire n1989;
    wire n1998;
    wire n1994;
    wire n2026;
    wire n1887;
    wire n1986;
    wire n1919_cascade_;
    wire n2018;
    wire n1988;
    wire n2020;
    wire n1987;
    wire n1991;
    wire n1892;
    wire n1924;
    wire n1924_cascade_;
    wire n1893;
    wire n1891;
    wire n1923_cascade_;
    wire n1896;
    wire n1899;
    wire n1822_cascade_;
    wire n1894;
    wire n1688;
    wire n1720_cascade_;
    wire n1820;
    wire n1752_cascade_;
    wire n1821;
    wire n13343;
    wire n14110_cascade_;
    wire n1653_cascade_;
    wire n1691;
    wire n13962;
    wire n11694;
    wire n13968_cascade_;
    wire n14116;
    wire n13972;
    wire n1690;
    wire n1628;
    wire n14104;
    wire n1624;
    wire n1692;
    wire n1626;
    wire n1693;
    wire n1632;
    wire n1632_cascade_;
    wire n1633;
    wire n11634;
    wire n1625;
    wire n1623;
    wire n1499;
    wire n1531_cascade_;
    wire n11698;
    wire n1627;
    wire n1430;
    wire n1497;
    wire n1498;
    wire n1622;
    wire n300;
    wire n1501;
    wire n300_cascade_;
    wire n1490;
    wire n1522_cascade_;
    wire n1621;
    wire n1495;
    wire n1496;
    wire n1528_cascade_;
    wire n13978_cascade_;
    wire n13984;
    wire n1432;
    wire n14088;
    wire n1433;
    wire n1433_cascade_;
    wire n1500;
    wire n1401;
    wire bfn_3_29_0_;
    wire n1400;
    wire n12141;
    wire n12142;
    wire n1398;
    wire n12143;
    wire n12144;
    wire n12145;
    wire n1395;
    wire n12146;
    wire n12147;
    wire n12148;
    wire bfn_3_30_0_;
    wire n12149;
    wire n12150;
    wire n12151;
    wire bfn_3_31_0_;
    wire n12131;
    wire n1299;
    wire n12132;
    wire n1298;
    wire n12133;
    wire n12134;
    wire n12135;
    wire n12136;
    wire n12137;
    wire n12138;
    wire bfn_3_32_0_;
    wire n12139;
    wire n12140;
    wire reg_B_2;
    wire \debounce.n6 ;
    wire \debounce.reg_A_2 ;
    wire \debounce.cnt_next_9__N_418 ;
    wire n1193;
    wire n2198;
    wire n2230_cascade_;
    wire n2189;
    wire n2221_cascade_;
    wire n2320_cascade_;
    wire n2387;
    wire n2399;
    wire n2397;
    wire n2429_cascade_;
    wire n14210_cascade_;
    wire n14214_cascade_;
    wire n13423;
    wire n2396;
    wire n2329;
    wire n14016_cascade_;
    wire n14022_cascade_;
    wire n2395;
    wire n2346_cascade_;
    wire n2384;
    wire n2385;
    wire n2389;
    wire n2317;
    wire n14410;
    wire n11774_cascade_;
    wire n14188_cascade_;
    wire n2187;
    wire n2219_cascade_;
    wire n2318;
    wire n2330;
    wire n2099;
    wire n1997;
    wire n2029;
    wire n2030;
    wire n2029_cascade_;
    wire n14154;
    wire n1990;
    wire n1923;
    wire n2022;
    wire n2022_cascade_;
    wire n14146;
    wire n14152;
    wire n1928;
    wire n1995;
    wire n2027;
    wire n2023;
    wire n2090;
    wire n2122;
    wire n2128;
    wire n2122_cascade_;
    wire n1918;
    wire n1919;
    wire n1926;
    wire n1950_cascade_;
    wire n1993;
    wire n1999;
    wire n2031;
    wire n2031_cascade_;
    wire n11680;
    wire n1992;
    wire n1925;
    wire n1819;
    wire n14134;
    wire n1851_cascade_;
    wire n1895;
    wire n1927;
    wire n1890;
    wire n1922;
    wire n13772;
    wire n1922_cascade_;
    wire n13770;
    wire n1920;
    wire n13778_cascade_;
    wire n13782;
    wire bfn_4_24_0_;
    wire n1733;
    wire n1800;
    wire n12191;
    wire n1732;
    wire n1799;
    wire n12192;
    wire n1731;
    wire n1798;
    wire n12193;
    wire n1730;
    wire n1797;
    wire n12194;
    wire n12195;
    wire n1728;
    wire n1795;
    wire n12196;
    wire n1727;
    wire n1794;
    wire n12197;
    wire n12198;
    wire bfn_4_25_0_;
    wire n1725;
    wire n1792;
    wire n12199;
    wire n12200;
    wire n1723;
    wire n1790;
    wire n12201;
    wire n1722;
    wire n1789;
    wire n12202;
    wire n1721;
    wire n1788;
    wire n12203;
    wire n1720;
    wire n1787;
    wire n12204;
    wire n1719;
    wire n12205;
    wire n1601;
    wire bfn_4_26_0_;
    wire n1533;
    wire n1600;
    wire n12164;
    wire n1532;
    wire n1599;
    wire n12165;
    wire n1531;
    wire n1598;
    wire n12166;
    wire n1530;
    wire n1597;
    wire n12167;
    wire n1529;
    wire n1596;
    wire n12168;
    wire n1528;
    wire n1595;
    wire n12169;
    wire n1527;
    wire n1594;
    wire n12170;
    wire n12171;
    wire n1593;
    wire bfn_4_27_0_;
    wire n1592;
    wire n12172;
    wire n1591;
    wire n12173;
    wire n1523;
    wire n1590;
    wire n12174;
    wire n1522;
    wire n1589;
    wire n12175;
    wire n1521;
    wire n12176;
    wire n1620;
    wire n1427;
    wire n1494;
    wire n1526;
    wire n1493;
    wire n1525;
    wire n1396;
    wire n1428;
    wire n1393;
    wire n1394;
    wire n1426;
    wire n1399;
    wire n1431;
    wire n1391;
    wire n1423;
    wire n1422;
    wire n13334;
    wire n1423_cascade_;
    wire n14094;
    wire n1425;
    wire n1455_cascade_;
    wire n1492;
    wire n1524;
    wire n1301;
    wire n1333;
    wire n1333_cascade_;
    wire n11640_cascade_;
    wire n1331;
    wire n1323;
    wire n13315_cascade_;
    wire n1356_cascade_;
    wire n1392;
    wire n1424;
    wire n299;
    wire n1330;
    wire n1397;
    wire n1429;
    wire n1297;
    wire n1329;
    wire n1295;
    wire n1294;
    wire n1224;
    wire n1257_cascade_;
    wire n1201;
    wire n1300;
    wire n1233_cascade_;
    wire n1332;
    wire n1296;
    wire n1194;
    wire n1200;
    wire n1225;
    wire n1292;
    wire n1324;
    wire n1158_cascade_;
    wire n1199;
    wire n1197;
    wire n1130;
    wire n1130_cascade_;
    wire n14068;
    wire n11706;
    wire n2527_cascade_;
    wire n13798;
    wire n13796_cascade_;
    wire n14354_cascade_;
    wire n14220;
    wire n14224_cascade_;
    wire n2445_cascade_;
    wire n2517_cascade_;
    wire n13804;
    wire n2185;
    wire n2390;
    wire n2401;
    wire n2433_cascade_;
    wire n11670;
    wire n2383;
    wire n2314;
    wire n2381;
    wire n2314_cascade_;
    wire n2326_cascade_;
    wire n2393;
    wire n2400;
    wire n14194;
    wire n2247_cascade_;
    wire n2333;
    wire n2332;
    wire n2333_cascade_;
    wire n2331;
    wire n11766;
    wire n2190;
    wire n2133;
    wire n2129;
    wire n2130;
    wire n11616_cascade_;
    wire n2131;
    wire n2001;
    wire n2033;
    wire n2100;
    wire n2033_cascade_;
    wire n2132;
    wire n2199;
    wire n2132_cascade_;
    wire n2000;
    wire n2032;
    wire n2091;
    wire n2024;
    wire n2123;
    wire n2123_cascade_;
    wire n2121;
    wire n13746_cascade_;
    wire n13748;
    wire n2119;
    wire n13754_cascade_;
    wire n13382;
    wire n13760;
    wire n1822;
    wire n1889;
    wire n1921;
    wire n1900;
    wire n1932;
    wire n1932_cascade_;
    wire n1931;
    wire n11686;
    wire n1897;
    wire n1929;
    wire n1929_cascade_;
    wire n14136;
    wire n1901;
    wire n1933;
    wire n1898;
    wire n1930;
    wire n1885;
    wire n1818;
    wire n1917;
    wire n1791;
    wire n1724;
    wire n1823;
    wire n1824;
    wire n1823_cascade_;
    wire n1830;
    wire n1829;
    wire n14126_cascade_;
    wire n14128;
    wire n1793;
    wire n1726;
    wire n1825;
    wire n1827;
    wire n1826;
    wire n1825_cascade_;
    wire n14122;
    wire n1729;
    wire n1796;
    wire n1828;
    wire n1832;
    wire n1831;
    wire n11688;
    wire n2021;
    wire n2088;
    wire n2120;
    wire n301;
    wire n1801;
    wire n303;
    wire n1833;
    wire n307;
    wire n13490;
    wire n306;
    wire n13257_cascade_;
    wire n302;
    wire bfn_5_28_0_;
    wire n12096;
    wire n12097;
    wire n2287;
    wire n12098;
    wire n12099;
    wire n402;
    wire n12100;
    wire n2289;
    wire n13261_cascade_;
    wire n297;
    wire \debounce.reg_A_1 ;
    wire reg_B_1;
    wire \debounce.reg_A_0 ;
    wire reg_B_0;
    wire n2288;
    wire n1293;
    wire n1325;
    wire n1326;
    wire n1327;
    wire n1325_cascade_;
    wire n1328;
    wire n13734;
    wire n298;
    wire n1233;
    wire n298_cascade_;
    wire n1232;
    wire n1196;
    wire n1228;
    wire n1228_cascade_;
    wire n1226;
    wire n14078;
    wire n1132;
    wire n1129;
    wire n1133;
    wire n1195;
    wire n1227;
    wire n1198;
    wire n1230;
    wire n1229;
    wire n1231;
    wire n1230_cascade_;
    wire n11642;
    wire n13318;
    wire n1125;
    wire n1126;
    wire n1126_cascade_;
    wire n1127;
    wire n13994;
    wire bfn_6_14_0_;
    wire n12339;
    wire n12340;
    wire n12341;
    wire n12342;
    wire n12343;
    wire n12344;
    wire n12345;
    wire n12346;
    wire bfn_6_15_0_;
    wire n12347;
    wire n12348;
    wire n12349;
    wire n12350;
    wire n12351;
    wire n12352;
    wire n12353;
    wire n12354;
    wire bfn_6_16_0_;
    wire n12355;
    wire n12356;
    wire n12357;
    wire n2581;
    wire n12358;
    wire n12359;
    wire n12360;
    wire n12361;
    wire bfn_6_17_0_;
    wire n12317;
    wire n12318;
    wire n12319;
    wire n2430;
    wire n2497;
    wire n12320;
    wire n2429;
    wire n2496;
    wire n12321;
    wire n2428;
    wire n2495;
    wire n12322;
    wire n2427;
    wire n2494;
    wire n12323;
    wire n12324;
    wire n2493;
    wire bfn_6_18_0_;
    wire n12325;
    wire n12326;
    wire n2490;
    wire n12327;
    wire n2422;
    wire n2489;
    wire n12328;
    wire n12329;
    wire n12330;
    wire n2419;
    wire n2486;
    wire n12331;
    wire n12332;
    wire n2418;
    wire n2485;
    wire bfn_6_19_0_;
    wire n12333;
    wire n12334;
    wire n2415;
    wire n2482;
    wire n12335;
    wire n12336;
    wire n12337;
    wire n2412;
    wire n12338;
    wire n2421;
    wire n2488;
    wire n2126;
    wire n2193;
    wire n2192;
    wire n2125;
    wire n2224_cascade_;
    wire n14174_cascade_;
    wire n14178_cascade_;
    wire n14184;
    wire n2500;
    wire n2433;
    wire n2431;
    wire n2498;
    wire n2194;
    wire n2127;
    wire n2501;
    wire n2533_cascade_;
    wire n11682_cascade_;
    wire n13397;
    wire n2086;
    wire n2019;
    wire n2118;
    wire n2432;
    wire n2499;
    wire n2025;
    wire n2092;
    wire n2124;
    wire n2191;
    wire n2124_cascade_;
    wire n2223_cascade_;
    wire n2315;
    wire n2382;
    wire n2315_cascade_;
    wire n2414;
    wire n2414_cascade_;
    wire n2481;
    wire bfn_6_23_0_;
    wire \quad_counter0.n12623 ;
    wire \quad_counter0.n12624 ;
    wire \quad_counter0.n12625 ;
    wire \quad_counter0.n12626 ;
    wire \quad_counter0.n12627 ;
    wire \quad_counter0.n12628 ;
    wire \quad_counter0.n12629 ;
    wire \quad_counter0.n12630 ;
    wire bfn_6_24_0_;
    wire \quad_counter0.n12631 ;
    wire \quad_counter0.n12632 ;
    wire \quad_counter0.n12633 ;
    wire encoder0_position_12;
    wire \quad_counter0.n12634 ;
    wire \quad_counter0.n12635 ;
    wire \quad_counter0.n12636 ;
    wire \quad_counter0.n12637 ;
    wire \quad_counter0.n12638 ;
    wire bfn_6_25_0_;
    wire encoder0_position_17;
    wire \quad_counter0.n12639 ;
    wire encoder0_position_18;
    wire \quad_counter0.n12640 ;
    wire encoder0_position_19;
    wire \quad_counter0.n12641 ;
    wire encoder0_position_20;
    wire \quad_counter0.n12642 ;
    wire encoder0_position_21;
    wire \quad_counter0.n12643 ;
    wire encoder0_position_22;
    wire \quad_counter0.n12644 ;
    wire \quad_counter0.n12645 ;
    wire \quad_counter0.n12646 ;
    wire bfn_6_26_0_;
    wire \quad_counter0.n12647 ;
    wire \quad_counter0.n12648 ;
    wire \quad_counter0.n12649 ;
    wire \quad_counter0.n12650 ;
    wire \quad_counter0.n12651 ;
    wire \quad_counter0.n12652 ;
    wire \quad_counter0.n12653 ;
    wire encoder0_position_16;
    wire encoder0_position_27;
    wire n175;
    wire encoder0_position_29;
    wire n404;
    wire n14170_cascade_;
    wire n2285;
    wire n293;
    wire n293_cascade_;
    wire n5_adj_697;
    wire n5_adj_697_cascade_;
    wire n2290;
    wire n13254_cascade_;
    wire n13259;
    wire n13263;
    wire n174;
    wire n13254;
    wire n2286;
    wire n13255_cascade_;
    wire encoder0_position_26;
    wire encoder0_position_30;
    wire n403;
    wire n11712_cascade_;
    wire n861_cascade_;
    wire encoder0_position_24;
    wire n1101;
    wire bfn_6_31_0_;
    wire n1100;
    wire n12114;
    wire n12115;
    wire n1098;
    wire n12116;
    wire n1097;
    wire n12117;
    wire n12118;
    wire n1095;
    wire n12119;
    wire n1094;
    wire n12120;
    wire n12121;
    wire bfn_6_32_0_;
    wire n1093;
    wire n1096;
    wire n1128;
    wire n1028;
    wire n1027;
    wire n1059_cascade_;
    wire n1099;
    wire n1131;
    wire encoder0_position_23;
    wire n2590;
    wire n2592;
    wire n2525;
    wire n2517;
    wire n2584;
    wire n2595;
    wire n2528;
    wire n2491;
    wire n2424;
    wire n2523;
    wire n2583;
    wire n2596;
    wire n2529;
    wire n2628_cascade_;
    wire n2585;
    wire n2518;
    wire n2417;
    wire n2484;
    wire n2516;
    wire n2514;
    wire n2516_cascade_;
    wire n13810;
    wire n13816_cascade_;
    wire n2511;
    wire n2582;
    wire n2544_cascade_;
    wire n2579;
    wire n2425;
    wire n2492;
    wire n2524;
    wire n2591;
    wire n2524_cascade_;
    wire n2391;
    wire n2423;
    wire n2601;
    wire n2394;
    wire n2426;
    wire n2480;
    wire n2413;
    wire n2512;
    wire n2388;
    wire n2420;
    wire n2487;
    wire n2420_cascade_;
    wire n2519;
    wire n2519_cascade_;
    wire n2586;
    wire n2532;
    wire n2599;
    wire n2483;
    wire n2416;
    wire n2515;
    wire n2301;
    wire bfn_7_20_0_;
    wire n2233;
    wire n2300;
    wire n12276;
    wire n2232;
    wire n2299;
    wire n12277;
    wire n2231;
    wire n2298;
    wire n12278;
    wire n2230;
    wire n2297;
    wire n12279;
    wire n2229;
    wire n2296;
    wire n12280;
    wire n12281;
    wire n2227;
    wire n2294;
    wire n12282;
    wire n12283;
    wire n2226;
    wire n2293;
    wire bfn_7_21_0_;
    wire n12284;
    wire n12285;
    wire n2223;
    wire n2290_adj_604;
    wire n12286;
    wire n2222;
    wire n2289_adj_603;
    wire n12287;
    wire n2221;
    wire n2288_adj_602;
    wire n12288;
    wire n2220;
    wire n2287_adj_601;
    wire n12289;
    wire n2219;
    wire n2286_adj_600;
    wire n12290;
    wire n12291;
    wire n2218;
    wire n2285_adj_599;
    wire bfn_7_22_0_;
    wire n12292;
    wire n2216;
    wire n2283;
    wire n12293;
    wire n2215;
    wire n2282;
    wire n12294;
    wire n2214;
    wire n12295;
    wire n2313;
    wire n2225;
    wire n2292;
    wire n2224;
    wire n2291;
    wire n2295;
    wire n2228;
    wire encoder0_position_2;
    wire n2321;
    wire n2324;
    wire n2328;
    wire n2327;
    wire n2322;
    wire n2326;
    wire n2325;
    wire n2323;
    wire encoder0_position_3;
    wire encoder0_position_11;
    wire n308;
    wire encoder0_position_8;
    wire n311;
    wire encoder0_position_5;
    wire encoder0_position_15;
    wire n304;
    wire n2320;
    wire n2319;
    wire n14008;
    wire n14006;
    wire n14014;
    wire encoder0_position_1;
    wire encoder0_position_0;
    wire n33_adj_657;
    wire n33;
    wire bfn_7_25_0_;
    wire n32_adj_656;
    wire n32;
    wire n12575;
    wire n31_adj_655;
    wire n31;
    wire n12576;
    wire n30_adj_654;
    wire n30;
    wire n12577;
    wire n29_adj_653;
    wire n12578;
    wire n28_adj_652;
    wire n28;
    wire n12579;
    wire n27;
    wire n12580;
    wire n26_adj_650;
    wire n12581;
    wire n12582;
    wire n25_adj_649;
    wire n25;
    wire bfn_7_26_0_;
    wire n24_adj_648;
    wire n12583;
    wire n23_adj_647;
    wire n12584;
    wire n22_adj_646;
    wire n22;
    wire n12585;
    wire n21_adj_645;
    wire n21;
    wire n12586;
    wire n20;
    wire n12587;
    wire n19_adj_643;
    wire n12588;
    wire n18_adj_642;
    wire n18;
    wire n12589;
    wire n12590;
    wire n17_adj_641;
    wire n17;
    wire bfn_7_27_0_;
    wire n16_adj_640;
    wire n16;
    wire n12591;
    wire n15_adj_639;
    wire n15;
    wire n12592;
    wire n14_adj_638;
    wire n14;
    wire n12593;
    wire n13_adj_637;
    wire n13;
    wire n12594;
    wire n12_adj_636;
    wire n12;
    wire n12595;
    wire n11_adj_635;
    wire n11;
    wire n12596;
    wire n10_adj_634;
    wire n10;
    wire n12597;
    wire n12598;
    wire n9_adj_633;
    wire n9;
    wire bfn_7_28_0_;
    wire n8_adj_632;
    wire n12599;
    wire n7_adj_631;
    wire n7;
    wire n12600;
    wire n6_adj_630;
    wire n6;
    wire n12601;
    wire n5;
    wire n12602;
    wire n4_adj_628;
    wire n4;
    wire n12603;
    wire n3_adj_627;
    wire n3_adj_567;
    wire n12604;
    wire n12605;
    wire n2_adj_568;
    wire n901;
    wire bfn_7_29_0_;
    wire n12101;
    wire n832;
    wire n899;
    wire n12102;
    wire n12103;
    wire n830;
    wire n897;
    wire n12104;
    wire n829;
    wire n896;
    wire n12105;
    wire n828;
    wire n12106;
    wire n900;
    wire n833;
    wire bfn_7_30_0_;
    wire n12107;
    wire n12108;
    wire n12109;
    wire n12110;
    wire n996;
    wire n12111;
    wire n995;
    wire n12112;
    wire n12113;
    wire n1026;
    wire n997;
    wire n999;
    wire n932;
    wire n898;
    wire n831;
    wire n861;
    wire n930;
    wire n930_cascade_;
    wire n929;
    wire n927;
    wire n928;
    wire n13726_cascade_;
    wire n11710;
    wire n1000;
    wire n960_cascade_;
    wire n933;
    wire n295;
    wire n1001;
    wire n931;
    wire n960;
    wire n998;
    wire n1032;
    wire n296;
    wire n1033;
    wire n1031;
    wire n1029;
    wire n11646_cascade_;
    wire n1030;
    wire n13323;
    wire n2531;
    wire n2598;
    wire n2630_cascade_;
    wire n14288_cascade_;
    wire n2527;
    wire n2594;
    wire n2626_cascade_;
    wire n14278;
    wire n14280_cascade_;
    wire n14286;
    wire n2522;
    wire n2589;
    wire n2597;
    wire n2530;
    wire n2520;
    wire n2587;
    wire n2580;
    wire n2513;
    wire n2721_cascade_;
    wire n2526;
    wire n2593;
    wire n2625_cascade_;
    wire bfn_9_19_0_;
    wire n12362;
    wire n12363;
    wire n12364;
    wire n12365;
    wire n12366;
    wire n12367;
    wire n12368;
    wire n12369;
    wire bfn_9_20_0_;
    wire n2625;
    wire n2692;
    wire n12370;
    wire n12371;
    wire n12372;
    wire n2622;
    wire n2689;
    wire n12373;
    wire n12374;
    wire n12375;
    wire n12376;
    wire n12377;
    wire bfn_9_21_0_;
    wire n12378;
    wire n12379;
    wire n12380;
    wire n12381;
    wire n12382;
    wire n12383;
    wire n12384;
    wire n12385;
    wire bfn_9_22_0_;
    wire n11750_cascade_;
    wire n13900_cascade_;
    wire n3232_cascade_;
    wire n13906;
    wire n13912_cascade_;
    wire n3138_cascade_;
    wire n3229_cascade_;
    wire n11658;
    wire bfn_9_25_0_;
    wire n12552;
    wire n12553;
    wire n12554;
    wire n12555;
    wire n12556;
    wire n12557;
    wire n15437;
    wire n12558;
    wire n12559;
    wire n15401;
    wire bfn_9_26_0_;
    wire n15375;
    wire n2445;
    wire n12560;
    wire n15348;
    wire n2346;
    wire n12561;
    wire n15322;
    wire n12562;
    wire n15059;
    wire n2148;
    wire n12563;
    wire n15035;
    wire n2049;
    wire n12564;
    wire n15012;
    wire n1950;
    wire n12565;
    wire n14990;
    wire n1851;
    wire n12566;
    wire n12567;
    wire n14969;
    wire n1752;
    wire bfn_9_27_0_;
    wire n14949;
    wire n1653;
    wire n12568;
    wire n15292;
    wire n1554;
    wire n12569;
    wire n15276;
    wire n1455;
    wire n12570;
    wire n15259;
    wire n1356;
    wire n12571;
    wire n15243;
    wire n1257;
    wire n12572;
    wire n15224;
    wire n1158;
    wire n12573;
    wire n2_adj_626;
    wire n12574;
    wire encoder0_position_scaled_17;
    wire encoder0_position_scaled_20;
    wire encoder0_position_25;
    wire n8;
    wire n294;
    wire encoder0_position_scaled_23;
    wire ENCODER0_A_N;
    wire n1059;
    wire n15210;
    wire n14536_cascade_;
    wire blink_counter_25;
    wire LED_c;
    wire blink_counter_24;
    wire blink_counter_21;
    wire blink_counter_22;
    wire blink_counter_23;
    wire n14535;
    wire n14294;
    wire n2693;
    wire n2626;
    wire n2725_cascade_;
    wire n14040_cascade_;
    wire n2629;
    wire n2696;
    wire n2630;
    wire n2697;
    wire n2695;
    wire n2628;
    wire n2619;
    wire n2686;
    wire n2627;
    wire n2694;
    wire n2521;
    wire n2588;
    wire n2620;
    wire n2687;
    wire n2620_cascade_;
    wire n2610;
    wire n14300;
    wire n2621;
    wire n2643_cascade_;
    wire n2688;
    wire n2720_cascade_;
    wire n14038_cascade_;
    wire n14042;
    wire n2614;
    wire n2681;
    wire n2685;
    wire n2618;
    wire encoder0_position_6;
    wire n27_adj_651;
    wire n24;
    wire encoder0_position_9;
    wire n310;
    wire n19;
    wire encoder0_position_14;
    wire n305;
    wire n23;
    wire encoder0_position_10;
    wire n309;
    wire n2616;
    wire n2683;
    wire n13884_cascade_;
    wire n3117_cascade_;
    wire n13888;
    wire n13886;
    wire bfn_10_21_0_;
    wire n12437;
    wire n12438;
    wire n12439;
    wire n12440;
    wire n12441;
    wire n12442;
    wire n12443;
    wire n12444;
    wire bfn_10_22_0_;
    wire n12445;
    wire n12446;
    wire n12447;
    wire n12448;
    wire n12449;
    wire n12450;
    wire n12451;
    wire n12452;
    wire bfn_10_23_0_;
    wire n12453;
    wire n12454;
    wire n12455;
    wire n12456;
    wire n12457;
    wire n12458;
    wire n12459;
    wire n12460;
    wire bfn_10_24_0_;
    wire n12461;
    wire n12462;
    wire n12463;
    wire n15197;
    wire n11593_cascade_;
    wire n59_cascade_;
    wire n11838;
    wire encoder0_position_scaled_0;
    wire encoder0_position_scaled_15;
    wire encoder0_position_scaled_12;
    wire encoder0_position_scaled_2;
    wire encoder0_position_scaled_4;
    wire dti_N_333_cascade_;
    wire encoder0_position_scaled_22;
    wire n26;
    wire encoder0_position_7;
    wire encoder0_position_scaled_19;
    wire encoder0_position_scaled_21;
    wire encoder0_position_scaled_13;
    wire n4828;
    wire encoder0_position_13;
    wire n20_adj_644;
    wire encoder0_position_28;
    wire n5_adj_629;
    wire encoder0_position_scaled_9;
    wire encoder0_position_scaled_10;
    wire h2;
    wire h3;
    wire h1;
    wire n6_adj_592;
    wire commutation_state_7__N_261;
    wire n41_cascade_;
    wire n41;
    wire n14715_cascade_;
    wire n40;
    wire n14866_cascade_;
    wire n12_adj_598_cascade_;
    wire n45_cascade_;
    wire n16_adj_614;
    wire n14843_cascade_;
    wire n24_adj_619;
    wire n14711_cascade_;
    wire n8_adj_607;
    wire n45;
    wire n14826_cascade_;
    wire n14779;
    wire n14864;
    wire n43;
    wire n14713;
    wire n2700;
    wire n2732_cascade_;
    wire n11666_cascade_;
    wire n2691;
    wire n2624;
    wire n2617;
    wire n2684;
    wire n2701;
    wire n2613;
    wire n2680;
    wire n2611;
    wire n2678;
    wire n2615;
    wire n2682;
    wire n2714_cascade_;
    wire n2623;
    wire n2690;
    wire n2698;
    wire n2699;
    wire n2217;
    wire n2284;
    wire n2247;
    wire n2316;
    wire n2533;
    wire n2600;
    wire n2544;
    wire n2632;
    wire n312;
    wire n2633;
    wire n2632_cascade_;
    wire n2631;
    wire n11760;
    wire n2817_cascade_;
    wire n3000;
    wire n3032_cascade_;
    wire n11660_cascade_;
    wire n2986;
    wire n2997;
    wire n3029_cascade_;
    wire encoder0_position_31;
    wire n29;
    wire encoder0_position_4;
    wire n3001;
    wire n315_cascade_;
    wire n2998;
    wire n3115_cascade_;
    wire n13894;
    wire n13898;
    wire n2988;
    wire n2987;
    wire n3019_cascade_;
    wire n2983;
    wire n2981;
    wire n2984;
    wire n2912_cascade_;
    wire n2979;
    wire n2975;
    wire n2980;
    wire n2976;
    wire n2978;
    wire n3010_cascade_;
    wire n15090;
    wire n14392_cascade_;
    wire n13470;
    wire n14380_cascade_;
    wire n14386;
    wire n14398;
    wire n3237_cascade_;
    wire n61;
    wire n13856_cascade_;
    wire n13858_cascade_;
    wire n13860_cascade_;
    wire n13862_cascade_;
    wire n13864_cascade_;
    wire n13866;
    wire encoder0_position_scaled_5;
    wire encoder0_position_scaled_8;
    wire encoder0_position_scaled_11;
    wire encoder0_position_scaled_7;
    wire encoder0_position_scaled_1;
    wire n4_adj_698_cascade_;
    wire pwm_setpoint_21;
    wire encoder0_position_scaled_14;
    wire encoder0_position_scaled_16;
    wire encoder0_position_scaled_18;
    wire commutation_state_prev_2;
    wire bfn_11_29_0_;
    wire \PWM.n12686 ;
    wire \PWM.n12687 ;
    wire \PWM.n12688 ;
    wire pwm_counter_4;
    wire \PWM.n12689 ;
    wire \PWM.n12690 ;
    wire \PWM.n12691 ;
    wire \PWM.n12692 ;
    wire \PWM.n12693 ;
    wire bfn_11_30_0_;
    wire \PWM.n12694 ;
    wire \PWM.n12695 ;
    wire pwm_counter_11;
    wire \PWM.n12696 ;
    wire \PWM.n12697 ;
    wire \PWM.n12698 ;
    wire \PWM.n12699 ;
    wire \PWM.n12700 ;
    wire \PWM.n12701 ;
    wire bfn_11_31_0_;
    wire \PWM.n12702 ;
    wire \PWM.n12703 ;
    wire \PWM.n12704 ;
    wire pwm_counter_20;
    wire \PWM.n12705 ;
    wire pwm_counter_21;
    wire \PWM.n12706 ;
    wire pwm_counter_22;
    wire \PWM.n12707 ;
    wire \PWM.n12708 ;
    wire \PWM.n12709 ;
    wire pwm_counter_24;
    wire bfn_11_32_0_;
    wire pwm_counter_25;
    wire \PWM.n12710 ;
    wire pwm_counter_26;
    wire \PWM.n12711 ;
    wire pwm_counter_27;
    wire \PWM.n12712 ;
    wire pwm_counter_28;
    wire \PWM.n12713 ;
    wire pwm_counter_29;
    wire \PWM.n12714 ;
    wire pwm_counter_30;
    wire \PWM.n12715 ;
    wire \PWM.n12716 ;
    wire bfn_12_17_0_;
    wire n12386;
    wire n12387;
    wire n12388;
    wire n12389;
    wire n12390;
    wire n12391;
    wire n12392;
    wire n12393;
    wire bfn_12_18_0_;
    wire n12394;
    wire n12395;
    wire n12396;
    wire n12397;
    wire n2721;
    wire n2788;
    wire n12398;
    wire n12399;
    wire n12400;
    wire n12401;
    wire n2718;
    wire n2785;
    wire bfn_12_19_0_;
    wire n2717;
    wire n2784;
    wire n12402;
    wire n12403;
    wire n12404;
    wire n2781;
    wire n12405;
    wire n12406;
    wire n12407;
    wire n12408;
    wire n12409;
    wire n2777;
    wire bfn_12_20_0_;
    wire n12410;
    wire n2985;
    wire n3017_cascade_;
    wire n2977;
    wire n2993;
    wire n2911;
    wire n2912;
    wire n13948_cascade_;
    wire n13954_cascade_;
    wire n2999;
    wire n2940_cascade_;
    wire n2996;
    wire n14340_cascade_;
    wire n2908;
    wire n14344;
    wire n3039_cascade_;
    wire n13466;
    wire n14334;
    wire n3121_cascade_;
    wire n3112_cascade_;
    wire n23_adj_707_cascade_;
    wire n25_adj_708_cascade_;
    wire n13832_cascade_;
    wire n13828;
    wire n13826;
    wire n13840_cascade_;
    wire n13846;
    wire n13848_cascade_;
    wire n5_adj_713;
    wire n13850_cascade_;
    wire n11656;
    wire n13852_cascade_;
    wire n13854;
    wire n37_adj_710;
    wire n7_adj_703;
    wire n14_adj_679_cascade_;
    wire n4781_cascade_;
    wire n14700;
    wire n1259;
    wire dti_counter_0;
    wire bfn_12_27_0_;
    wire n14693;
    wire n12742;
    wire n14692;
    wire n12743;
    wire n14691;
    wire dti_counter_3;
    wire n12744;
    wire n14690;
    wire dti_counter_4;
    wire n12745;
    wire n12746;
    wire n14688;
    wire dti_counter_6;
    wire n12747;
    wire n14687;
    wire n11202;
    wire n12748;
    wire dti_counter_7;
    wire pwm_setpoint_4;
    wire pwm_counter_2;
    wire pwm_counter_3;
    wire pwm_setpoint_3;
    wire n4_adj_698;
    wire dti_counter_5;
    wire commutation_state_prev_0;
    wire n14689;
    wire pwm_setpoint_2;
    wire pwm_setpoint_11;
    wire pwm_setpoint_8;
    wire pwm_counter_10;
    wire n21_adj_617_cascade_;
    wire n6_adj_606;
    wire n14842;
    wire pwm_setpoint_10;
    wire n11_adj_610_cascade_;
    wire pwm_setpoint_5;
    wire pwm_setpoint_6;
    wire n4825;
    wire n13_adj_612;
    wire n11_adj_610;
    wire n14745;
    wire pwm_setpoint_20;
    wire pwm_counter_5;
    wire pwm_counter_6;
    wire \PWM.n13596_cascade_ ;
    wire pwm_counter_8;
    wire \PWM.n26 ;
    wire n4823;
    wire \PWM.n17_cascade_ ;
    wire pwm_counter_31;
    wire \PWM.n29_cascade_ ;
    wire \PWM.n27 ;
    wire \PWM.pwm_counter_31__N_401 ;
    wire pwm_counter_19;
    wire n39;
    wire pwm_setpoint_19;
    wire n39_cascade_;
    wire n14883;
    wire pwm_counter_9;
    wire n14804;
    wire n19_adj_616_cascade_;
    wire n15_adj_613;
    wire n23_adj_618;
    wire n14800_cascade_;
    wire n19_adj_616;
    wire n17_adj_615;
    wire n9_adj_608;
    wire n21_adj_617;
    wire n14734;
    wire n14874;
    wire pwm_setpoint_12;
    wire pwm_counter_12;
    wire n25_adj_620;
    wire n2723;
    wire n2790;
    wire n2725;
    wire n2792;
    wire n13403;
    wire n14048;
    wire n2714;
    wire n14054_cascade_;
    wire n2710;
    wire n14060_cascade_;
    wire n2709;
    wire n2798;
    wire n2742_cascade_;
    wire n2731;
    wire n2728;
    wire n2795;
    wire n14238_cascade_;
    wire n14240_cascade_;
    wire n2720;
    wire n2787;
    wire n2789;
    wire n2722;
    wire n2797;
    wire n2730;
    wire n2724;
    wire n2791;
    wire n2786;
    wire n2719;
    wire n2921;
    wire n2921_cascade_;
    wire n2778;
    wire n2917;
    wire n2918;
    wire n13926;
    wire n2917_cascade_;
    wire n2916;
    wire n13934_cascade_;
    wire n13942;
    wire n2679;
    wire n2612;
    wire n2643;
    wire n2711;
    wire n15467;
    wire n2909;
    wire n2713;
    wire n2780;
    wire n14322_cascade_;
    wire n14328;
    wire n2992;
    wire n2991;
    wire n3023_cascade_;
    wire n14320;
    wire n2995;
    wire n2994;
    wire n2913;
    wire n2990;
    wire n2982;
    wire n2915;
    wire n3014_cascade_;
    wire n14408;
    wire n2940;
    wire n2989;
    wire n3021_cascade_;
    wire n319;
    wire bfn_13_23_0_;
    wire n318;
    wire n3301;
    wire n12521;
    wire n3233;
    wire n3300;
    wire n12522;
    wire n3232;
    wire n3299;
    wire n12523;
    wire n3231;
    wire n12524;
    wire n3298;
    wire n3230;
    wire n14697;
    wire n12525;
    wire n12526;
    wire n12527;
    wire n12528;
    wire bfn_13_24_0_;
    wire n3293;
    wire n12529;
    wire n12530;
    wire n3291;
    wire n12531;
    wire n3290;
    wire n12532;
    wire n12533;
    wire n3288;
    wire n12534;
    wire n12535;
    wire n12536;
    wire bfn_13_25_0_;
    wire n3285;
    wire n12537;
    wire n3217;
    wire n3284;
    wire n12538;
    wire n3216;
    wire n3283;
    wire n12539;
    wire n3215;
    wire n3282;
    wire n12540;
    wire n3214;
    wire n3281;
    wire n12541;
    wire n3280;
    wire n12542;
    wire n3212;
    wire n3279;
    wire n12543;
    wire n12544;
    wire n3211;
    wire n3278;
    wire bfn_13_26_0_;
    wire n3210;
    wire n3277;
    wire n12545;
    wire n3276;
    wire n12546;
    wire n3208;
    wire n3275;
    wire n12547;
    wire n3207;
    wire n3274;
    wire n12548;
    wire n3206;
    wire n3273;
    wire n12549;
    wire n3205;
    wire n3272;
    wire n12550;
    wire n15163;
    wire n12551;
    wire n14461;
    wire encoder0_position_scaled_3;
    wire dti_counter_2;
    wire dti_counter_1;
    wire n10_adj_680;
    wire n25_adj_591;
    wire bfn_13_28_0_;
    wire n12050;
    wire n23_adj_589;
    wire pwm_setpoint_23_N_171_2;
    wire n12051;
    wire pwm_setpoint_23_N_171_3;
    wire n12052;
    wire n21_adj_587;
    wire pwm_setpoint_23_N_171_4;
    wire n12053;
    wire n20_adj_586;
    wire pwm_setpoint_23_N_171_5;
    wire n12054;
    wire n19_adj_585;
    wire pwm_setpoint_23_N_171_6;
    wire n12055;
    wire n18_adj_584;
    wire n12056;
    wire n12057;
    wire pwm_setpoint_23_N_171_8;
    wire bfn_13_29_0_;
    wire n12058;
    wire n15_adj_581;
    wire pwm_setpoint_23_N_171_10;
    wire n12059;
    wire n14_adj_580;
    wire pwm_setpoint_23_N_171_11;
    wire n12060;
    wire pwm_setpoint_23_N_171_12;
    wire n12061;
    wire n12062;
    wire n11_adj_577;
    wire n12063;
    wire n12064;
    wire n12065;
    wire bfn_13_30_0_;
    wire n12066;
    wire n12067;
    wire pwm_setpoint_23_N_171_19;
    wire n12068;
    wire pwm_setpoint_23_N_171_20;
    wire n12069;
    wire n4_adj_570;
    wire pwm_setpoint_23_N_171_21;
    wire n12070;
    wire n12071;
    wire n12072;
    wire pwm_setpoint_23;
    wire pwm_setpoint_23_N_171_15;
    wire pwm_setpoint_23_N_171_18;
    wire pwm_counter_23;
    wire \PWM.n28 ;
    wire pwm_counter_15;
    wire pwm_counter_18;
    wire n37;
    wire pwm_setpoint_18;
    wire n37_cascade_;
    wire n14887;
    wire pwm_setpoint_23_N_171_22;
    wire pwm_setpoint_22;
    wire pwm_setpoint_23_N_171_17;
    wire n14870;
    wire n14832;
    wire pwm_counter_17;
    wire n2712;
    wire n2779;
    wire n2811_cascade_;
    wire n2794;
    wire n2727;
    wire n2716;
    wire n2783;
    wire n2782;
    wire n2715;
    wire n2814_cascade_;
    wire n14260;
    wire n2796;
    wire n2729;
    wire n2800;
    wire n2733;
    wire n2799;
    wire n2732;
    wire n14246;
    wire n14248_cascade_;
    wire n14254_cascade_;
    wire n14266;
    wire n2841_cascade_;
    wire n2923;
    wire n13932_cascade_;
    wire n13936;
    wire n2926;
    wire n2920;
    wire n2927;
    wire n2919;
    wire n2928;
    wire n2922;
    wire n2793;
    wire n2726;
    wire n2825_cascade_;
    wire n2924;
    wire n2925;
    wire n3122_cascade_;
    wire n2914;
    wire n316;
    wire n3101;
    wire bfn_14_21_0_;
    wire n3033;
    wire n3100;
    wire n12464;
    wire n3032;
    wire n3099;
    wire n12465;
    wire n3031;
    wire n3098;
    wire n12466;
    wire n3030;
    wire n3097;
    wire n12467;
    wire n3029;
    wire n3096;
    wire n12468;
    wire n3028;
    wire n3095;
    wire n12469;
    wire n3027;
    wire n3094;
    wire n12470;
    wire n12471;
    wire n3026;
    wire n3093;
    wire bfn_14_22_0_;
    wire n3025;
    wire n3092;
    wire n12472;
    wire n3024;
    wire n3091;
    wire n12473;
    wire n3023;
    wire n3090;
    wire n12474;
    wire n3022;
    wire n3089;
    wire n12475;
    wire n3021;
    wire n3088;
    wire n12476;
    wire n3020;
    wire n3087;
    wire n12477;
    wire n3019;
    wire n3086;
    wire n12478;
    wire n12479;
    wire n3018;
    wire n3085;
    wire bfn_14_23_0_;
    wire n3017;
    wire n3084;
    wire n12480;
    wire n3016;
    wire n3083;
    wire n12481;
    wire n12482;
    wire n3014;
    wire n3081;
    wire n12483;
    wire n3013;
    wire n3080;
    wire n12484;
    wire n3012;
    wire n3079;
    wire n12485;
    wire n12486;
    wire n12487;
    wire n3010;
    wire n3077;
    wire bfn_14_24_0_;
    wire n12488;
    wire n3008;
    wire n3075;
    wire n12489;
    wire n3007;
    wire n3074;
    wire n12490;
    wire n3006;
    wire n15123;
    wire n12491;
    wire n3295;
    wire n3294;
    wire n3221;
    wire n3218;
    wire n14368_cascade_;
    wire n14374;
    wire n3228;
    wire n3228_cascade_;
    wire n3224;
    wire n14362;
    wire n3223;
    wire n14366;
    wire n3227;
    wire n25_adj_545;
    wire bfn_14_26_0_;
    wire n24_adj_546;
    wire n12073;
    wire n23_adj_547;
    wire duty_2;
    wire n12074;
    wire n22_adj_548;
    wire n12075;
    wire n21_adj_549;
    wire duty_4;
    wire n12076;
    wire n20_adj_550;
    wire duty_5;
    wire n12077;
    wire duty_6;
    wire n12078;
    wire n18_adj_552;
    wire n12079;
    wire n12080;
    wire n17_adj_553;
    wire bfn_14_27_0_;
    wire n16_adj_554;
    wire n12081;
    wire n15_adj_555;
    wire duty_10;
    wire n12082;
    wire n14_adj_556;
    wire duty_11;
    wire n12083;
    wire n13_adj_557;
    wire n12084;
    wire n12_adj_558;
    wire n12085;
    wire n11_adj_559;
    wire n12086;
    wire n10_adj_560;
    wire n12087;
    wire n12088;
    wire n9_adj_561;
    wire bfn_14_28_0_;
    wire n8_adj_562;
    wire n12089;
    wire n7_adj_563;
    wire n12090;
    wire n6_adj_564;
    wire n12091;
    wire n5_adj_565;
    wire n12092;
    wire n4_adj_566;
    wire duty_21;
    wire n12093;
    wire n3;
    wire n12094;
    wire n2;
    wire n12095;
    wire pwm_setpoint_23_N_171_13;
    wire duty_15;
    wire n10_adj_576;
    wire duty_14;
    wire pwm_setpoint_23_N_171_14;
    wire pwm_counter_1;
    wire pwm_counter_0;
    wire n16_adj_582;
    wire duty_13;
    wire n12_adj_578;
    wire pwm_setpoint_23_N_171_0;
    wire duty_0;
    wire pwm_setpoint_0;
    wire duty_12;
    wire n13_adj_579;
    wire pwm_counter_14;
    wire pwm_counter_13;
    wire n27_adj_621;
    wire pwm_setpoint_13;
    wire n27_adj_621_cascade_;
    wire n4_adj_605;
    wire pwm_setpoint_14;
    wire n14840_cascade_;
    wire duty_22;
    wire n3_adj_569;
    wire n9_adj_575;
    wire duty_16;
    wire pwm_setpoint_23_N_171_16;
    wire duty_20;
    wire n5_adj_571;
    wire pwm_counter_7;
    wire n10_adj_609;
    wire n14722_cascade_;
    wire n14876_cascade_;
    wire n14886;
    wire pwm_setpoint_15;
    wire n14841;
    wire n14781;
    wire pwm_setpoint_23_N_171_7;
    wire duty_7;
    wire pwm_setpoint_7;
    wire pwm_setpoint_17;
    wire n12_adj_611_cascade_;
    wire n35;
    wire n30_adj_623;
    wire pwm_setpoint_16;
    wire pwm_counter_16;
    wire n33_adj_625;
    wire n31_adj_624;
    wire n14728;
    wire n33_adj_625_cascade_;
    wire n29_adj_622;
    wire n14724;
    wire duty_17;
    wire n8_adj_574;
    wire n28_adj_597;
    wire n31_adj_594;
    wire n32_adj_593_cascade_;
    wire n2910;
    wire n30_adj_595;
    wire n29_adj_596;
    wire n2801;
    wire n313;
    wire n2742;
    wire n2833_cascade_;
    wire n11756;
    wire n2932;
    wire n315;
    wire n2932_cascade_;
    wire n2933;
    wire n2930;
    wire n2931;
    wire n2929;
    wire n2930_cascade_;
    wire n11662;
    wire n13417;
    wire n314;
    wire n2901;
    wire bfn_15_20_0_;
    wire n2833;
    wire n2900;
    wire n12411;
    wire n2832;
    wire n2899;
    wire n12412;
    wire n2831;
    wire n2898;
    wire n12413;
    wire n2830;
    wire n2897;
    wire n12414;
    wire n2829;
    wire n2896;
    wire n12415;
    wire n2828;
    wire n2895;
    wire n12416;
    wire n2827;
    wire n2894;
    wire n12417;
    wire n12418;
    wire n2826;
    wire n2893;
    wire bfn_15_21_0_;
    wire n2825;
    wire n2892;
    wire n12419;
    wire n2824;
    wire n2891;
    wire n12420;
    wire n2823;
    wire n2890;
    wire n12421;
    wire n2822;
    wire n2889;
    wire n12422;
    wire n2821;
    wire n2888;
    wire n12423;
    wire n2820;
    wire n2887;
    wire n12424;
    wire n2819;
    wire n2886;
    wire n12425;
    wire n12426;
    wire n2818;
    wire n2885;
    wire bfn_15_22_0_;
    wire n2817;
    wire n2884;
    wire n12427;
    wire n2816;
    wire n2883;
    wire n12428;
    wire n2815;
    wire n2882;
    wire n12429;
    wire n2814;
    wire n2881;
    wire n12430;
    wire n2813;
    wire n2880;
    wire n12431;
    wire n2812;
    wire n2879;
    wire n12432;
    wire n2811;
    wire n2878;
    wire n12433;
    wire n12434;
    wire n2810;
    wire n2877;
    wire bfn_15_23_0_;
    wire n2809;
    wire n2876;
    wire n12435;
    wire n12436;
    wire n2808;
    wire n2875;
    wire n2907;
    wire n3220;
    wire n3287;
    wire n17_adj_705;
    wire n3296;
    wire n13822_cascade_;
    wire n3229;
    wire n15_adj_704;
    wire n13834_cascade_;
    wire n13842;
    wire n3222;
    wire n3289;
    wire n3286;
    wire n27_adj_709_cascade_;
    wire n3219;
    wire n13830;
    wire n3292;
    wire n3225;
    wire n3237;
    wire n21_adj_706;
    wire n3011;
    wire n3078;
    wire n3110_cascade_;
    wire n3209;
    wire n3226;
    wire n2841;
    wire n14921;
    wire n3009;
    wire n3076;
    wire ENCODER0_B_N;
    wire n3015;
    wire n3082;
    wire n3039;
    wire n3138;
    wire n3114_cascade_;
    wire n3213;
    wire n7_adj_712_cascade_;
    wire n8_adj_711;
    wire \quad_counter0.direction_N_530 ;
    wire n13676;
    wire n10_adj_714_cascade_;
    wire n16_adj_702_cascade_;
    wire n19_adj_701;
    wire n24_adj_590;
    wire duty_3;
    wire n22_adj_588;
    wire n21_adj_700_cascade_;
    wire n22_adj_699;
    wire duty_1;
    wire pwm_setpoint_23_N_171_1;
    wire pwm_setpoint_1;
    wire \quad_counter0.a_prev_N_537_cascade_ ;
    wire \quad_counter0.direction_N_534_cascade_ ;
    wire \quad_counter0.a_prev_N_537 ;
    wire \quad_counter0.a_prev ;
    wire \quad_counter0.b_new_1 ;
    wire \quad_counter0.b_new_0 ;
    wire \quad_counter0.debounce_cnt ;
    wire direction_N_531;
    wire b_prev;
    wire n1185;
    wire \quad_counter0.a_new_0 ;
    wire a_new_1;
    wire duty_19;
    wire n6_adj_572;
    wire duty_18;
    wire n7_adj_573;
    wire sweep_counter_0;
    wire bfn_16_17_0_;
    wire sweep_counter_1;
    wire n12606;
    wire sweep_counter_2;
    wire n12607;
    wire sweep_counter_3;
    wire n12608;
    wire sweep_counter_4;
    wire n12609;
    wire sweep_counter_5;
    wire n12610;
    wire sweep_counter_6;
    wire n12611;
    wire sweep_counter_7;
    wire n12612;
    wire n12613;
    wire sweep_counter_8;
    wire bfn_16_18_0_;
    wire sweep_counter_9;
    wire n12614;
    wire sweep_counter_10;
    wire n12615;
    wire sweep_counter_11;
    wire n12616;
    wire sweep_counter_12;
    wire n12617;
    wire sweep_counter_13;
    wire n12618;
    wire sweep_counter_14;
    wire n12619;
    wire sweep_counter_15;
    wire n12620;
    wire n12621;
    wire sweep_counter_16;
    wire bfn_16_19_0_;
    wire n12622;
    wire sweep_counter_17;
    wire n317;
    wire n3201;
    wire bfn_16_22_0_;
    wire n3133;
    wire n3200;
    wire n12492;
    wire n3132;
    wire n3199;
    wire n12493;
    wire n3131;
    wire n3198;
    wire n12494;
    wire n3130;
    wire n3197;
    wire n12495;
    wire n3129;
    wire n3196;
    wire n12496;
    wire n3128;
    wire n3195;
    wire n12497;
    wire n3127;
    wire n3194;
    wire n12498;
    wire n12499;
    wire n3126;
    wire n3193;
    wire bfn_16_23_0_;
    wire n3125;
    wire n3192;
    wire n12500;
    wire n3124;
    wire n3191;
    wire n12501;
    wire n3123;
    wire n3190;
    wire n12502;
    wire n3122;
    wire n3189;
    wire n12503;
    wire n3121;
    wire n3188;
    wire n12504;
    wire n3120;
    wire n3187;
    wire n12505;
    wire n3119;
    wire n3186;
    wire n12506;
    wire n12507;
    wire n3118;
    wire n3185;
    wire bfn_16_24_0_;
    wire n3117;
    wire n3184;
    wire n12508;
    wire n3116;
    wire n3183;
    wire n12509;
    wire n3115;
    wire n3182;
    wire n12510;
    wire n3114;
    wire n3181;
    wire n12511;
    wire n3113;
    wire n3180;
    wire n12512;
    wire n3112;
    wire n3179;
    wire n12513;
    wire n3111;
    wire n3178;
    wire n12514;
    wire n12515;
    wire n3110;
    wire n3177;
    wire bfn_16_25_0_;
    wire n3109;
    wire n3176;
    wire n12516;
    wire n3108;
    wire n3175;
    wire n12517;
    wire n3107;
    wire n3174;
    wire n12518;
    wire n3106;
    wire n3173;
    wire n12519;
    wire n15158;
    wire n3105;
    wire n12520;
    wire n3204;
    wire encoder0_position_target_0;
    wire bfn_16_26_0_;
    wire encoder0_position_target_1;
    wire n12663;
    wire encoder0_position_target_2;
    wire n12664;
    wire encoder0_position_target_3;
    wire n12665;
    wire encoder0_position_target_4;
    wire n12666;
    wire encoder0_position_target_5;
    wire n12667;
    wire encoder0_position_target_6;
    wire n12668;
    wire encoder0_position_target_7;
    wire n12669;
    wire n12670;
    wire encoder0_position_target_8;
    wire bfn_16_27_0_;
    wire encoder0_position_target_9;
    wire n12671;
    wire encoder0_position_target_10;
    wire n12672;
    wire encoder0_position_target_11;
    wire n12673;
    wire encoder0_position_target_12;
    wire n12674;
    wire encoder0_position_target_13;
    wire n12675;
    wire encoder0_position_target_14;
    wire n12676;
    wire encoder0_position_target_15;
    wire n12677;
    wire n12678;
    wire encoder0_position_target_16;
    wire bfn_16_28_0_;
    wire encoder0_position_target_17;
    wire n12679;
    wire encoder0_position_target_18;
    wire n12680;
    wire encoder0_position_target_19;
    wire n12681;
    wire encoder0_position_target_20;
    wire n12682;
    wire encoder0_position_target_21;
    wire n12683;
    wire encoder0_position_target_22;
    wire n12684;
    wire CONSTANT_ONE_NET;
    wire n12685;
    wire encoder0_position_target_23;
    wire n4856;
    wire n4890;
    wire pwm_setpoint_23_N_171_9;
    wire duty_9;
    wire pwm_setpoint_9;
    wire duty_8;
    wire n17_adj_583;
    wire commutation_state_prev_1;
    wire duty_23;
    wire pwm_setpoint_23__N_195;
    wire encoder0_position_scaled_6;
    wire n19_adj_551;
    wire dti;
    wire n4781;
    wire INLC_c_0;
    wire INLA_c_0;
    wire INLB_c_0;
    wire dir;
    wire commutation_state_1;
    wire commutation_state_0;
    wire commutation_state_2;
    wire CLK_N;
    wire n4842;
    wire n4886;
    wire GHA;
    wire INHA_c_0;
    wire GHC;
    wire INHC_c_0;
    wire GHB;
    wire pwm_out;
    wire INHB_c_0;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__56636),
            .DIN(N__56635),
            .DOUT(N__56634),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__56636),
            .PADOUT(N__56635),
            .PADIN(N__56634),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__56627),
            .DIN(N__56626),
            .DOUT(N__56625),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__56627),
            .PADOUT(N__56626),
            .PADIN(N__56625),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__56618),
            .DIN(N__56617),
            .DOUT(N__56616),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__56618),
            .PADOUT(N__56617),
            .PADIN(N__56616),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_A_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_A_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_A_pad_iopad (
            .OE(N__56609),
            .DIN(N__56608),
            .DOUT(N__56607),
            .PACKAGEPIN(ENCODER0_A));
    defparam ENCODER0_A_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_A_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_A_pad_preio (
            .PADOEN(N__56609),
            .PADOUT(N__56608),
            .PADIN(N__56607),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_A_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_B_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_B_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_B_pad_iopad (
            .OE(N__56600),
            .DIN(N__56599),
            .DOUT(N__56598),
            .PACKAGEPIN(ENCODER0_B));
    defparam ENCODER0_B_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_B_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_B_pad_preio (
            .PADOEN(N__56600),
            .PADOUT(N__56599),
            .PADIN(N__56598),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_B_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__56591),
            .DIN(N__56590),
            .DOUT(N__56589),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__56591),
            .PADOUT(N__56590),
            .PADIN(N__56589),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55810),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__56582),
            .DIN(N__56581),
            .DOUT(N__56580),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__56582),
            .PADOUT(N__56581),
            .PADIN(N__56580),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55744),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__56573),
            .DIN(N__56572),
            .DOUT(N__56571),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__56573),
            .PADOUT(N__56572),
            .PADIN(N__56571),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55789),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__56564),
            .DIN(N__56563),
            .DOUT(N__56562),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__56564),
            .PADOUT(N__56563),
            .PADIN(N__56562),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55411),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__56555),
            .DIN(N__56554),
            .DOUT(N__56553),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__56555),
            .PADOUT(N__56554),
            .PADIN(N__56553),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56455),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__56546),
            .DIN(N__56545),
            .DOUT(N__56544),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__56546),
            .PADOUT(N__56545),
            .PADIN(N__56544),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55426),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__56537),
            .DIN(N__56536),
            .DOUT(N__56535),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__56537),
            .PADOUT(N__56536),
            .PADIN(N__56535),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36871),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__56528),
            .DIN(N__56527),
            .DOUT(N__56526),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__56528),
            .PADOUT(N__56527),
            .PADIN(N__56526),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__56519),
            .DIN(N__56518),
            .DOUT(N__56517),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__56519),
            .PADOUT(N__56518),
            .PADIN(N__56517),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__56510),
            .DIN(N__56509),
            .DOUT(N__56508),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__56510),
            .PADOUT(N__56509),
            .PADIN(N__56508),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__56501),
            .DIN(N__56500),
            .DOUT(N__56499),
            .PACKAGEPIN(HALL1));
    defparam hall1_input_preio.PIN_TYPE=6'b000000;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__56501),
            .PADOUT(N__56500),
            .PADIN(N__56499),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_2 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56041),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__56492),
            .DIN(N__56491),
            .DOUT(N__56490),
            .PACKAGEPIN(HALL2));
    defparam hall2_input_preio.PIN_TYPE=6'b000000;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__56492),
            .PADOUT(N__56491),
            .PADIN(N__56490),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_1 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56039),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__56483),
            .DIN(N__56482),
            .DOUT(N__56481),
            .PACKAGEPIN(HALL3));
    defparam hall3_input_preio.PIN_TYPE=6'b000000;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__56483),
            .PADOUT(N__56482),
            .PADIN(N__56481),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_0 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56039),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__56474),
            .DIN(N__56473),
            .DOUT(N__56472),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__56474),
            .PADOUT(N__56473),
            .PADIN(N__56472),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__13460 (
            .O(N__56455),
            .I(N__56452));
    LocalMux I__13459 (
            .O(N__56452),
            .I(N__56449));
    IoSpan4Mux I__13458 (
            .O(N__56449),
            .I(N__56446));
    Span4Mux_s1_v I__13457 (
            .O(N__56446),
            .I(N__56443));
    Span4Mux_h I__13456 (
            .O(N__56443),
            .I(N__56440));
    Odrv4 I__13455 (
            .O(N__56440),
            .I(INLB_c_0));
    InMux I__13454 (
            .O(N__56437),
            .I(N__56431));
    InMux I__13453 (
            .O(N__56436),
            .I(N__56424));
    InMux I__13452 (
            .O(N__56435),
            .I(N__56424));
    CascadeMux I__13451 (
            .O(N__56434),
            .I(N__56421));
    LocalMux I__13450 (
            .O(N__56431),
            .I(N__56418));
    InMux I__13449 (
            .O(N__56430),
            .I(N__56413));
    InMux I__13448 (
            .O(N__56429),
            .I(N__56413));
    LocalMux I__13447 (
            .O(N__56424),
            .I(N__56410));
    InMux I__13446 (
            .O(N__56421),
            .I(N__56407));
    Span4Mux_s2_v I__13445 (
            .O(N__56418),
            .I(N__56404));
    LocalMux I__13444 (
            .O(N__56413),
            .I(N__56399));
    Span4Mux_s2_v I__13443 (
            .O(N__56410),
            .I(N__56399));
    LocalMux I__13442 (
            .O(N__56407),
            .I(dir));
    Odrv4 I__13441 (
            .O(N__56404),
            .I(dir));
    Odrv4 I__13440 (
            .O(N__56399),
            .I(dir));
    InMux I__13439 (
            .O(N__56392),
            .I(N__56383));
    InMux I__13438 (
            .O(N__56391),
            .I(N__56383));
    InMux I__13437 (
            .O(N__56390),
            .I(N__56377));
    InMux I__13436 (
            .O(N__56389),
            .I(N__56377));
    InMux I__13435 (
            .O(N__56388),
            .I(N__56371));
    LocalMux I__13434 (
            .O(N__56383),
            .I(N__56368));
    InMux I__13433 (
            .O(N__56382),
            .I(N__56365));
    LocalMux I__13432 (
            .O(N__56377),
            .I(N__56362));
    InMux I__13431 (
            .O(N__56376),
            .I(N__56359));
    InMux I__13430 (
            .O(N__56375),
            .I(N__56354));
    InMux I__13429 (
            .O(N__56374),
            .I(N__56354));
    LocalMux I__13428 (
            .O(N__56371),
            .I(N__56350));
    Span4Mux_v I__13427 (
            .O(N__56368),
            .I(N__56347));
    LocalMux I__13426 (
            .O(N__56365),
            .I(N__56344));
    Span4Mux_v I__13425 (
            .O(N__56362),
            .I(N__56341));
    LocalMux I__13424 (
            .O(N__56359),
            .I(N__56336));
    LocalMux I__13423 (
            .O(N__56354),
            .I(N__56336));
    CascadeMux I__13422 (
            .O(N__56353),
            .I(N__56333));
    Span4Mux_h I__13421 (
            .O(N__56350),
            .I(N__56330));
    Span4Mux_h I__13420 (
            .O(N__56347),
            .I(N__56323));
    Span4Mux_v I__13419 (
            .O(N__56344),
            .I(N__56323));
    Span4Mux_h I__13418 (
            .O(N__56341),
            .I(N__56323));
    Span4Mux_v I__13417 (
            .O(N__56336),
            .I(N__56320));
    InMux I__13416 (
            .O(N__56333),
            .I(N__56317));
    Span4Mux_v I__13415 (
            .O(N__56330),
            .I(N__56314));
    Sp12to4 I__13414 (
            .O(N__56323),
            .I(N__56309));
    Sp12to4 I__13413 (
            .O(N__56320),
            .I(N__56309));
    LocalMux I__13412 (
            .O(N__56317),
            .I(commutation_state_1));
    Odrv4 I__13411 (
            .O(N__56314),
            .I(commutation_state_1));
    Odrv12 I__13410 (
            .O(N__56309),
            .I(commutation_state_1));
    CascadeMux I__13409 (
            .O(N__56302),
            .I(N__56297));
    InMux I__13408 (
            .O(N__56301),
            .I(N__56291));
    InMux I__13407 (
            .O(N__56300),
            .I(N__56286));
    InMux I__13406 (
            .O(N__56297),
            .I(N__56286));
    InMux I__13405 (
            .O(N__56296),
            .I(N__56283));
    InMux I__13404 (
            .O(N__56295),
            .I(N__56278));
    InMux I__13403 (
            .O(N__56294),
            .I(N__56278));
    LocalMux I__13402 (
            .O(N__56291),
            .I(N__56272));
    LocalMux I__13401 (
            .O(N__56286),
            .I(N__56265));
    LocalMux I__13400 (
            .O(N__56283),
            .I(N__56265));
    LocalMux I__13399 (
            .O(N__56278),
            .I(N__56265));
    InMux I__13398 (
            .O(N__56277),
            .I(N__56260));
    InMux I__13397 (
            .O(N__56276),
            .I(N__56260));
    InMux I__13396 (
            .O(N__56275),
            .I(N__56257));
    Sp12to4 I__13395 (
            .O(N__56272),
            .I(N__56247));
    Span4Mux_s3_v I__13394 (
            .O(N__56265),
            .I(N__56244));
    LocalMux I__13393 (
            .O(N__56260),
            .I(N__56241));
    LocalMux I__13392 (
            .O(N__56257),
            .I(N__56238));
    InMux I__13391 (
            .O(N__56256),
            .I(N__56227));
    InMux I__13390 (
            .O(N__56255),
            .I(N__56227));
    InMux I__13389 (
            .O(N__56254),
            .I(N__56227));
    InMux I__13388 (
            .O(N__56253),
            .I(N__56227));
    InMux I__13387 (
            .O(N__56252),
            .I(N__56227));
    InMux I__13386 (
            .O(N__56251),
            .I(N__56224));
    InMux I__13385 (
            .O(N__56250),
            .I(N__56221));
    Span12Mux_s3_v I__13384 (
            .O(N__56247),
            .I(N__56216));
    Sp12to4 I__13383 (
            .O(N__56244),
            .I(N__56216));
    Span4Mux_v I__13382 (
            .O(N__56241),
            .I(N__56211));
    Span4Mux_v I__13381 (
            .O(N__56238),
            .I(N__56211));
    LocalMux I__13380 (
            .O(N__56227),
            .I(N__56206));
    LocalMux I__13379 (
            .O(N__56224),
            .I(N__56206));
    LocalMux I__13378 (
            .O(N__56221),
            .I(commutation_state_0));
    Odrv12 I__13377 (
            .O(N__56216),
            .I(commutation_state_0));
    Odrv4 I__13376 (
            .O(N__56211),
            .I(commutation_state_0));
    Odrv4 I__13375 (
            .O(N__56206),
            .I(commutation_state_0));
    CascadeMux I__13374 (
            .O(N__56197),
            .I(N__56191));
    CascadeMux I__13373 (
            .O(N__56196),
            .I(N__56188));
    CascadeMux I__13372 (
            .O(N__56195),
            .I(N__56184));
    CascadeMux I__13371 (
            .O(N__56194),
            .I(N__56181));
    InMux I__13370 (
            .O(N__56191),
            .I(N__56175));
    InMux I__13369 (
            .O(N__56188),
            .I(N__56175));
    InMux I__13368 (
            .O(N__56187),
            .I(N__56169));
    InMux I__13367 (
            .O(N__56184),
            .I(N__56169));
    InMux I__13366 (
            .O(N__56181),
            .I(N__56166));
    CascadeMux I__13365 (
            .O(N__56180),
            .I(N__56162));
    LocalMux I__13364 (
            .O(N__56175),
            .I(N__56159));
    CascadeMux I__13363 (
            .O(N__56174),
            .I(N__56156));
    LocalMux I__13362 (
            .O(N__56169),
            .I(N__56151));
    LocalMux I__13361 (
            .O(N__56166),
            .I(N__56151));
    InMux I__13360 (
            .O(N__56165),
            .I(N__56146));
    InMux I__13359 (
            .O(N__56162),
            .I(N__56146));
    Span4Mux_h I__13358 (
            .O(N__56159),
            .I(N__56142));
    InMux I__13357 (
            .O(N__56156),
            .I(N__56139));
    Span4Mux_h I__13356 (
            .O(N__56151),
            .I(N__56134));
    LocalMux I__13355 (
            .O(N__56146),
            .I(N__56134));
    InMux I__13354 (
            .O(N__56145),
            .I(N__56130));
    Span4Mux_h I__13353 (
            .O(N__56142),
            .I(N__56127));
    LocalMux I__13352 (
            .O(N__56139),
            .I(N__56124));
    Span4Mux_h I__13351 (
            .O(N__56134),
            .I(N__56121));
    InMux I__13350 (
            .O(N__56133),
            .I(N__56118));
    LocalMux I__13349 (
            .O(N__56130),
            .I(N__56115));
    Span4Mux_h I__13348 (
            .O(N__56127),
            .I(N__56112));
    Span4Mux_h I__13347 (
            .O(N__56124),
            .I(N__56107));
    Span4Mux_h I__13346 (
            .O(N__56121),
            .I(N__56107));
    LocalMux I__13345 (
            .O(N__56118),
            .I(commutation_state_2));
    Odrv4 I__13344 (
            .O(N__56115),
            .I(commutation_state_2));
    Odrv4 I__13343 (
            .O(N__56112),
            .I(commutation_state_2));
    Odrv4 I__13342 (
            .O(N__56107),
            .I(commutation_state_2));
    ClkMux I__13341 (
            .O(N__56098),
            .I(N__55918));
    ClkMux I__13340 (
            .O(N__56097),
            .I(N__55918));
    ClkMux I__13339 (
            .O(N__56096),
            .I(N__55918));
    ClkMux I__13338 (
            .O(N__56095),
            .I(N__55918));
    ClkMux I__13337 (
            .O(N__56094),
            .I(N__55918));
    ClkMux I__13336 (
            .O(N__56093),
            .I(N__55918));
    ClkMux I__13335 (
            .O(N__56092),
            .I(N__55918));
    ClkMux I__13334 (
            .O(N__56091),
            .I(N__55918));
    ClkMux I__13333 (
            .O(N__56090),
            .I(N__55918));
    ClkMux I__13332 (
            .O(N__56089),
            .I(N__55918));
    ClkMux I__13331 (
            .O(N__56088),
            .I(N__55918));
    ClkMux I__13330 (
            .O(N__56087),
            .I(N__55918));
    ClkMux I__13329 (
            .O(N__56086),
            .I(N__55918));
    ClkMux I__13328 (
            .O(N__56085),
            .I(N__55918));
    ClkMux I__13327 (
            .O(N__56084),
            .I(N__55918));
    ClkMux I__13326 (
            .O(N__56083),
            .I(N__55918));
    ClkMux I__13325 (
            .O(N__56082),
            .I(N__55918));
    ClkMux I__13324 (
            .O(N__56081),
            .I(N__55918));
    ClkMux I__13323 (
            .O(N__56080),
            .I(N__55918));
    ClkMux I__13322 (
            .O(N__56079),
            .I(N__55918));
    ClkMux I__13321 (
            .O(N__56078),
            .I(N__55918));
    ClkMux I__13320 (
            .O(N__56077),
            .I(N__55918));
    ClkMux I__13319 (
            .O(N__56076),
            .I(N__55918));
    ClkMux I__13318 (
            .O(N__56075),
            .I(N__55918));
    ClkMux I__13317 (
            .O(N__56074),
            .I(N__55918));
    ClkMux I__13316 (
            .O(N__56073),
            .I(N__55918));
    ClkMux I__13315 (
            .O(N__56072),
            .I(N__55918));
    ClkMux I__13314 (
            .O(N__56071),
            .I(N__55918));
    ClkMux I__13313 (
            .O(N__56070),
            .I(N__55918));
    ClkMux I__13312 (
            .O(N__56069),
            .I(N__55918));
    ClkMux I__13311 (
            .O(N__56068),
            .I(N__55918));
    ClkMux I__13310 (
            .O(N__56067),
            .I(N__55918));
    ClkMux I__13309 (
            .O(N__56066),
            .I(N__55918));
    ClkMux I__13308 (
            .O(N__56065),
            .I(N__55918));
    ClkMux I__13307 (
            .O(N__56064),
            .I(N__55918));
    ClkMux I__13306 (
            .O(N__56063),
            .I(N__55918));
    ClkMux I__13305 (
            .O(N__56062),
            .I(N__55918));
    ClkMux I__13304 (
            .O(N__56061),
            .I(N__55918));
    ClkMux I__13303 (
            .O(N__56060),
            .I(N__55918));
    ClkMux I__13302 (
            .O(N__56059),
            .I(N__55918));
    ClkMux I__13301 (
            .O(N__56058),
            .I(N__55918));
    ClkMux I__13300 (
            .O(N__56057),
            .I(N__55918));
    ClkMux I__13299 (
            .O(N__56056),
            .I(N__55918));
    ClkMux I__13298 (
            .O(N__56055),
            .I(N__55918));
    ClkMux I__13297 (
            .O(N__56054),
            .I(N__55918));
    ClkMux I__13296 (
            .O(N__56053),
            .I(N__55918));
    ClkMux I__13295 (
            .O(N__56052),
            .I(N__55918));
    ClkMux I__13294 (
            .O(N__56051),
            .I(N__55918));
    ClkMux I__13293 (
            .O(N__56050),
            .I(N__55918));
    ClkMux I__13292 (
            .O(N__56049),
            .I(N__55918));
    ClkMux I__13291 (
            .O(N__56048),
            .I(N__55918));
    ClkMux I__13290 (
            .O(N__56047),
            .I(N__55918));
    ClkMux I__13289 (
            .O(N__56046),
            .I(N__55918));
    ClkMux I__13288 (
            .O(N__56045),
            .I(N__55918));
    ClkMux I__13287 (
            .O(N__56044),
            .I(N__55918));
    ClkMux I__13286 (
            .O(N__56043),
            .I(N__55918));
    ClkMux I__13285 (
            .O(N__56042),
            .I(N__55918));
    ClkMux I__13284 (
            .O(N__56041),
            .I(N__55918));
    ClkMux I__13283 (
            .O(N__56040),
            .I(N__55918));
    ClkMux I__13282 (
            .O(N__56039),
            .I(N__55918));
    GlobalMux I__13281 (
            .O(N__55918),
            .I(N__55915));
    gio2CtrlBuf I__13280 (
            .O(N__55915),
            .I(CLK_N));
    CEMux I__13279 (
            .O(N__55912),
            .I(N__55909));
    LocalMux I__13278 (
            .O(N__55909),
            .I(N__55905));
    CEMux I__13277 (
            .O(N__55908),
            .I(N__55902));
    Span4Mux_v I__13276 (
            .O(N__55905),
            .I(N__55897));
    LocalMux I__13275 (
            .O(N__55902),
            .I(N__55894));
    CEMux I__13274 (
            .O(N__55901),
            .I(N__55891));
    CEMux I__13273 (
            .O(N__55900),
            .I(N__55888));
    Span4Mux_s1_v I__13272 (
            .O(N__55897),
            .I(N__55884));
    Sp12to4 I__13271 (
            .O(N__55894),
            .I(N__55879));
    LocalMux I__13270 (
            .O(N__55891),
            .I(N__55879));
    LocalMux I__13269 (
            .O(N__55888),
            .I(N__55876));
    InMux I__13268 (
            .O(N__55887),
            .I(N__55873));
    Odrv4 I__13267 (
            .O(N__55884),
            .I(n4842));
    Odrv12 I__13266 (
            .O(N__55879),
            .I(n4842));
    Odrv4 I__13265 (
            .O(N__55876),
            .I(n4842));
    LocalMux I__13264 (
            .O(N__55873),
            .I(n4842));
    SRMux I__13263 (
            .O(N__55864),
            .I(N__55861));
    LocalMux I__13262 (
            .O(N__55861),
            .I(N__55856));
    SRMux I__13261 (
            .O(N__55860),
            .I(N__55852));
    SRMux I__13260 (
            .O(N__55859),
            .I(N__55849));
    Span4Mux_h I__13259 (
            .O(N__55856),
            .I(N__55846));
    SRMux I__13258 (
            .O(N__55855),
            .I(N__55843));
    LocalMux I__13257 (
            .O(N__55852),
            .I(N__55840));
    LocalMux I__13256 (
            .O(N__55849),
            .I(N__55837));
    Span4Mux_h I__13255 (
            .O(N__55846),
            .I(N__55832));
    LocalMux I__13254 (
            .O(N__55843),
            .I(N__55832));
    Span4Mux_h I__13253 (
            .O(N__55840),
            .I(N__55829));
    Span4Mux_h I__13252 (
            .O(N__55837),
            .I(N__55826));
    Span4Mux_s2_v I__13251 (
            .O(N__55832),
            .I(N__55823));
    Odrv4 I__13250 (
            .O(N__55829),
            .I(n4886));
    Odrv4 I__13249 (
            .O(N__55826),
            .I(n4886));
    Odrv4 I__13248 (
            .O(N__55823),
            .I(n4886));
    InMux I__13247 (
            .O(N__55816),
            .I(N__55813));
    LocalMux I__13246 (
            .O(N__55813),
            .I(GHA));
    IoInMux I__13245 (
            .O(N__55810),
            .I(N__55807));
    LocalMux I__13244 (
            .O(N__55807),
            .I(N__55804));
    IoSpan4Mux I__13243 (
            .O(N__55804),
            .I(N__55801));
    Span4Mux_s0_v I__13242 (
            .O(N__55801),
            .I(N__55798));
    Odrv4 I__13241 (
            .O(N__55798),
            .I(INHA_c_0));
    InMux I__13240 (
            .O(N__55795),
            .I(N__55792));
    LocalMux I__13239 (
            .O(N__55792),
            .I(GHC));
    IoInMux I__13238 (
            .O(N__55789),
            .I(N__55786));
    LocalMux I__13237 (
            .O(N__55786),
            .I(N__55783));
    Span12Mux_s2_v I__13236 (
            .O(N__55783),
            .I(N__55780));
    Odrv12 I__13235 (
            .O(N__55780),
            .I(INHC_c_0));
    InMux I__13234 (
            .O(N__55777),
            .I(N__55774));
    LocalMux I__13233 (
            .O(N__55774),
            .I(GHB));
    InMux I__13232 (
            .O(N__55771),
            .I(N__55768));
    LocalMux I__13231 (
            .O(N__55768),
            .I(N__55763));
    InMux I__13230 (
            .O(N__55767),
            .I(N__55758));
    InMux I__13229 (
            .O(N__55766),
            .I(N__55758));
    Span4Mux_s2_v I__13228 (
            .O(N__55763),
            .I(N__55755));
    LocalMux I__13227 (
            .O(N__55758),
            .I(N__55752));
    Sp12to4 I__13226 (
            .O(N__55755),
            .I(N__55747));
    Sp12to4 I__13225 (
            .O(N__55752),
            .I(N__55747));
    Odrv12 I__13224 (
            .O(N__55747),
            .I(pwm_out));
    IoInMux I__13223 (
            .O(N__55744),
            .I(N__55741));
    LocalMux I__13222 (
            .O(N__55741),
            .I(N__55738));
    Span4Mux_s2_v I__13221 (
            .O(N__55738),
            .I(N__55735));
    Span4Mux_h I__13220 (
            .O(N__55735),
            .I(N__55732));
    Odrv4 I__13219 (
            .O(N__55732),
            .I(INHB_c_0));
    InMux I__13218 (
            .O(N__55729),
            .I(N__55726));
    LocalMux I__13217 (
            .O(N__55726),
            .I(N__55723));
    Span4Mux_h I__13216 (
            .O(N__55723),
            .I(N__55720));
    Span4Mux_h I__13215 (
            .O(N__55720),
            .I(N__55717));
    Odrv4 I__13214 (
            .O(N__55717),
            .I(commutation_state_prev_1));
    CascadeMux I__13213 (
            .O(N__55714),
            .I(N__55703));
    InMux I__13212 (
            .O(N__55713),
            .I(N__55685));
    InMux I__13211 (
            .O(N__55712),
            .I(N__55685));
    InMux I__13210 (
            .O(N__55711),
            .I(N__55685));
    InMux I__13209 (
            .O(N__55710),
            .I(N__55685));
    InMux I__13208 (
            .O(N__55709),
            .I(N__55682));
    InMux I__13207 (
            .O(N__55708),
            .I(N__55679));
    InMux I__13206 (
            .O(N__55707),
            .I(N__55676));
    InMux I__13205 (
            .O(N__55706),
            .I(N__55673));
    InMux I__13204 (
            .O(N__55703),
            .I(N__55668));
    InMux I__13203 (
            .O(N__55702),
            .I(N__55668));
    InMux I__13202 (
            .O(N__55701),
            .I(N__55657));
    InMux I__13201 (
            .O(N__55700),
            .I(N__55657));
    InMux I__13200 (
            .O(N__55699),
            .I(N__55657));
    InMux I__13199 (
            .O(N__55698),
            .I(N__55657));
    InMux I__13198 (
            .O(N__55697),
            .I(N__55657));
    InMux I__13197 (
            .O(N__55696),
            .I(N__55648));
    InMux I__13196 (
            .O(N__55695),
            .I(N__55645));
    InMux I__13195 (
            .O(N__55694),
            .I(N__55641));
    LocalMux I__13194 (
            .O(N__55685),
            .I(N__55638));
    LocalMux I__13193 (
            .O(N__55682),
            .I(N__55633));
    LocalMux I__13192 (
            .O(N__55679),
            .I(N__55633));
    LocalMux I__13191 (
            .O(N__55676),
            .I(N__55628));
    LocalMux I__13190 (
            .O(N__55673),
            .I(N__55628));
    LocalMux I__13189 (
            .O(N__55668),
            .I(N__55623));
    LocalMux I__13188 (
            .O(N__55657),
            .I(N__55623));
    InMux I__13187 (
            .O(N__55656),
            .I(N__55618));
    InMux I__13186 (
            .O(N__55655),
            .I(N__55618));
    InMux I__13185 (
            .O(N__55654),
            .I(N__55615));
    InMux I__13184 (
            .O(N__55653),
            .I(N__55608));
    InMux I__13183 (
            .O(N__55652),
            .I(N__55608));
    InMux I__13182 (
            .O(N__55651),
            .I(N__55608));
    LocalMux I__13181 (
            .O(N__55648),
            .I(N__55605));
    LocalMux I__13180 (
            .O(N__55645),
            .I(N__55602));
    InMux I__13179 (
            .O(N__55644),
            .I(N__55599));
    LocalMux I__13178 (
            .O(N__55641),
            .I(N__55596));
    Span4Mux_h I__13177 (
            .O(N__55638),
            .I(N__55587));
    Span4Mux_v I__13176 (
            .O(N__55633),
            .I(N__55587));
    Span4Mux_v I__13175 (
            .O(N__55628),
            .I(N__55587));
    Span4Mux_v I__13174 (
            .O(N__55623),
            .I(N__55587));
    LocalMux I__13173 (
            .O(N__55618),
            .I(N__55576));
    LocalMux I__13172 (
            .O(N__55615),
            .I(N__55576));
    LocalMux I__13171 (
            .O(N__55608),
            .I(N__55576));
    Span4Mux_h I__13170 (
            .O(N__55605),
            .I(N__55576));
    Span4Mux_h I__13169 (
            .O(N__55602),
            .I(N__55576));
    LocalMux I__13168 (
            .O(N__55599),
            .I(duty_23));
    Odrv12 I__13167 (
            .O(N__55596),
            .I(duty_23));
    Odrv4 I__13166 (
            .O(N__55587),
            .I(duty_23));
    Odrv4 I__13165 (
            .O(N__55576),
            .I(duty_23));
    SRMux I__13164 (
            .O(N__55567),
            .I(N__55564));
    LocalMux I__13163 (
            .O(N__55564),
            .I(N__55560));
    InMux I__13162 (
            .O(N__55563),
            .I(N__55557));
    Sp12to4 I__13161 (
            .O(N__55560),
            .I(N__55552));
    LocalMux I__13160 (
            .O(N__55557),
            .I(N__55552));
    Span12Mux_s5_v I__13159 (
            .O(N__55552),
            .I(N__55549));
    Odrv12 I__13158 (
            .O(N__55549),
            .I(pwm_setpoint_23__N_195));
    InMux I__13157 (
            .O(N__55546),
            .I(N__55543));
    LocalMux I__13156 (
            .O(N__55543),
            .I(N__55540));
    Span4Mux_v I__13155 (
            .O(N__55540),
            .I(N__55537));
    Sp12to4 I__13154 (
            .O(N__55537),
            .I(N__55534));
    Odrv12 I__13153 (
            .O(N__55534),
            .I(encoder0_position_scaled_6));
    CascadeMux I__13152 (
            .O(N__55531),
            .I(N__55528));
    InMux I__13151 (
            .O(N__55528),
            .I(N__55525));
    LocalMux I__13150 (
            .O(N__55525),
            .I(N__55522));
    Span4Mux_v I__13149 (
            .O(N__55522),
            .I(N__55519));
    Odrv4 I__13148 (
            .O(N__55519),
            .I(n19_adj_551));
    InMux I__13147 (
            .O(N__55516),
            .I(N__55512));
    InMux I__13146 (
            .O(N__55515),
            .I(N__55509));
    LocalMux I__13145 (
            .O(N__55512),
            .I(N__55501));
    LocalMux I__13144 (
            .O(N__55509),
            .I(N__55501));
    InMux I__13143 (
            .O(N__55508),
            .I(N__55496));
    InMux I__13142 (
            .O(N__55507),
            .I(N__55496));
    InMux I__13141 (
            .O(N__55506),
            .I(N__55492));
    Span4Mux_v I__13140 (
            .O(N__55501),
            .I(N__55489));
    LocalMux I__13139 (
            .O(N__55496),
            .I(N__55486));
    InMux I__13138 (
            .O(N__55495),
            .I(N__55483));
    LocalMux I__13137 (
            .O(N__55492),
            .I(N__55476));
    Span4Mux_h I__13136 (
            .O(N__55489),
            .I(N__55476));
    Span4Mux_v I__13135 (
            .O(N__55486),
            .I(N__55476));
    LocalMux I__13134 (
            .O(N__55483),
            .I(dti));
    Odrv4 I__13133 (
            .O(N__55476),
            .I(dti));
    InMux I__13132 (
            .O(N__55471),
            .I(N__55466));
    InMux I__13131 (
            .O(N__55470),
            .I(N__55463));
    InMux I__13130 (
            .O(N__55469),
            .I(N__55460));
    LocalMux I__13129 (
            .O(N__55466),
            .I(N__55457));
    LocalMux I__13128 (
            .O(N__55463),
            .I(N__55454));
    LocalMux I__13127 (
            .O(N__55460),
            .I(N__55451));
    Span4Mux_s3_v I__13126 (
            .O(N__55457),
            .I(N__55448));
    Span4Mux_h I__13125 (
            .O(N__55454),
            .I(N__55444));
    Span4Mux_h I__13124 (
            .O(N__55451),
            .I(N__55441));
    Span4Mux_h I__13123 (
            .O(N__55448),
            .I(N__55438));
    InMux I__13122 (
            .O(N__55447),
            .I(N__55435));
    Odrv4 I__13121 (
            .O(N__55444),
            .I(n4781));
    Odrv4 I__13120 (
            .O(N__55441),
            .I(n4781));
    Odrv4 I__13119 (
            .O(N__55438),
            .I(n4781));
    LocalMux I__13118 (
            .O(N__55435),
            .I(n4781));
    IoInMux I__13117 (
            .O(N__55426),
            .I(N__55423));
    LocalMux I__13116 (
            .O(N__55423),
            .I(N__55420));
    Span12Mux_s1_v I__13115 (
            .O(N__55420),
            .I(N__55417));
    Span12Mux_h I__13114 (
            .O(N__55417),
            .I(N__55414));
    Odrv12 I__13113 (
            .O(N__55414),
            .I(INLC_c_0));
    IoInMux I__13112 (
            .O(N__55411),
            .I(N__55408));
    LocalMux I__13111 (
            .O(N__55408),
            .I(N__55405));
    Span4Mux_s1_v I__13110 (
            .O(N__55405),
            .I(N__55402));
    Span4Mux_h I__13109 (
            .O(N__55402),
            .I(N__55399));
    Odrv4 I__13108 (
            .O(N__55399),
            .I(INLA_c_0));
    CascadeMux I__13107 (
            .O(N__55396),
            .I(N__55393));
    InMux I__13106 (
            .O(N__55393),
            .I(N__55389));
    InMux I__13105 (
            .O(N__55392),
            .I(N__55386));
    LocalMux I__13104 (
            .O(N__55389),
            .I(N__55383));
    LocalMux I__13103 (
            .O(N__55386),
            .I(N__55377));
    Span4Mux_h I__13102 (
            .O(N__55383),
            .I(N__55377));
    InMux I__13101 (
            .O(N__55382),
            .I(N__55374));
    Odrv4 I__13100 (
            .O(N__55377),
            .I(encoder0_position_target_18));
    LocalMux I__13099 (
            .O(N__55374),
            .I(encoder0_position_target_18));
    InMux I__13098 (
            .O(N__55369),
            .I(n12680));
    CascadeMux I__13097 (
            .O(N__55366),
            .I(N__55363));
    InMux I__13096 (
            .O(N__55363),
            .I(N__55359));
    CascadeMux I__13095 (
            .O(N__55362),
            .I(N__55356));
    LocalMux I__13094 (
            .O(N__55359),
            .I(N__55353));
    InMux I__13093 (
            .O(N__55356),
            .I(N__55349));
    Span4Mux_h I__13092 (
            .O(N__55353),
            .I(N__55346));
    InMux I__13091 (
            .O(N__55352),
            .I(N__55343));
    LocalMux I__13090 (
            .O(N__55349),
            .I(encoder0_position_target_19));
    Odrv4 I__13089 (
            .O(N__55346),
            .I(encoder0_position_target_19));
    LocalMux I__13088 (
            .O(N__55343),
            .I(encoder0_position_target_19));
    InMux I__13087 (
            .O(N__55336),
            .I(n12681));
    CascadeMux I__13086 (
            .O(N__55333),
            .I(N__55330));
    InMux I__13085 (
            .O(N__55330),
            .I(N__55326));
    InMux I__13084 (
            .O(N__55329),
            .I(N__55322));
    LocalMux I__13083 (
            .O(N__55326),
            .I(N__55319));
    InMux I__13082 (
            .O(N__55325),
            .I(N__55316));
    LocalMux I__13081 (
            .O(N__55322),
            .I(encoder0_position_target_20));
    Odrv4 I__13080 (
            .O(N__55319),
            .I(encoder0_position_target_20));
    LocalMux I__13079 (
            .O(N__55316),
            .I(encoder0_position_target_20));
    InMux I__13078 (
            .O(N__55309),
            .I(n12682));
    CascadeMux I__13077 (
            .O(N__55306),
            .I(N__55302));
    CascadeMux I__13076 (
            .O(N__55305),
            .I(N__55299));
    InMux I__13075 (
            .O(N__55302),
            .I(N__55296));
    InMux I__13074 (
            .O(N__55299),
            .I(N__55292));
    LocalMux I__13073 (
            .O(N__55296),
            .I(N__55289));
    InMux I__13072 (
            .O(N__55295),
            .I(N__55286));
    LocalMux I__13071 (
            .O(N__55292),
            .I(encoder0_position_target_21));
    Odrv4 I__13070 (
            .O(N__55289),
            .I(encoder0_position_target_21));
    LocalMux I__13069 (
            .O(N__55286),
            .I(encoder0_position_target_21));
    InMux I__13068 (
            .O(N__55279),
            .I(n12683));
    CascadeMux I__13067 (
            .O(N__55276),
            .I(N__55273));
    InMux I__13066 (
            .O(N__55273),
            .I(N__55269));
    InMux I__13065 (
            .O(N__55272),
            .I(N__55265));
    LocalMux I__13064 (
            .O(N__55269),
            .I(N__55262));
    InMux I__13063 (
            .O(N__55268),
            .I(N__55259));
    LocalMux I__13062 (
            .O(N__55265),
            .I(encoder0_position_target_22));
    Odrv4 I__13061 (
            .O(N__55262),
            .I(encoder0_position_target_22));
    LocalMux I__13060 (
            .O(N__55259),
            .I(encoder0_position_target_22));
    InMux I__13059 (
            .O(N__55252),
            .I(n12684));
    CascadeMux I__13058 (
            .O(N__55249),
            .I(N__55243));
    CascadeMux I__13057 (
            .O(N__55248),
            .I(N__55240));
    CascadeMux I__13056 (
            .O(N__55247),
            .I(N__55237));
    CascadeMux I__13055 (
            .O(N__55246),
            .I(N__55230));
    InMux I__13054 (
            .O(N__55243),
            .I(N__55202));
    InMux I__13053 (
            .O(N__55240),
            .I(N__55202));
    InMux I__13052 (
            .O(N__55237),
            .I(N__55202));
    InMux I__13051 (
            .O(N__55236),
            .I(N__55193));
    InMux I__13050 (
            .O(N__55235),
            .I(N__55193));
    InMux I__13049 (
            .O(N__55234),
            .I(N__55193));
    InMux I__13048 (
            .O(N__55233),
            .I(N__55193));
    InMux I__13047 (
            .O(N__55230),
            .I(N__55180));
    InMux I__13046 (
            .O(N__55229),
            .I(N__55180));
    InMux I__13045 (
            .O(N__55228),
            .I(N__55175));
    InMux I__13044 (
            .O(N__55227),
            .I(N__55175));
    CascadeMux I__13043 (
            .O(N__55226),
            .I(N__55169));
    InMux I__13042 (
            .O(N__55225),
            .I(N__55156));
    InMux I__13041 (
            .O(N__55224),
            .I(N__55156));
    InMux I__13040 (
            .O(N__55223),
            .I(N__55153));
    InMux I__13039 (
            .O(N__55222),
            .I(N__55146));
    InMux I__13038 (
            .O(N__55221),
            .I(N__55146));
    InMux I__13037 (
            .O(N__55220),
            .I(N__55146));
    CascadeMux I__13036 (
            .O(N__55219),
            .I(N__55142));
    CascadeMux I__13035 (
            .O(N__55218),
            .I(N__55137));
    CascadeMux I__13034 (
            .O(N__55217),
            .I(N__55118));
    CascadeMux I__13033 (
            .O(N__55216),
            .I(N__55114));
    CascadeMux I__13032 (
            .O(N__55215),
            .I(N__55110));
    CascadeMux I__13031 (
            .O(N__55214),
            .I(N__55106));
    CascadeMux I__13030 (
            .O(N__55213),
            .I(N__55103));
    CascadeMux I__13029 (
            .O(N__55212),
            .I(N__55099));
    CascadeMux I__13028 (
            .O(N__55211),
            .I(N__55095));
    CascadeMux I__13027 (
            .O(N__55210),
            .I(N__55091));
    CascadeMux I__13026 (
            .O(N__55209),
            .I(N__55073));
    LocalMux I__13025 (
            .O(N__55202),
            .I(N__55057));
    LocalMux I__13024 (
            .O(N__55193),
            .I(N__55054));
    InMux I__13023 (
            .O(N__55192),
            .I(N__55047));
    InMux I__13022 (
            .O(N__55191),
            .I(N__55047));
    InMux I__13021 (
            .O(N__55190),
            .I(N__55047));
    CascadeMux I__13020 (
            .O(N__55189),
            .I(N__55044));
    CascadeMux I__13019 (
            .O(N__55188),
            .I(N__55041));
    CascadeMux I__13018 (
            .O(N__55187),
            .I(N__55038));
    CascadeMux I__13017 (
            .O(N__55186),
            .I(N__55035));
    CascadeMux I__13016 (
            .O(N__55185),
            .I(N__55031));
    LocalMux I__13015 (
            .O(N__55180),
            .I(N__55026));
    LocalMux I__13014 (
            .O(N__55175),
            .I(N__55026));
    InMux I__13013 (
            .O(N__55174),
            .I(N__55019));
    InMux I__13012 (
            .O(N__55173),
            .I(N__55019));
    InMux I__13011 (
            .O(N__55172),
            .I(N__55019));
    InMux I__13010 (
            .O(N__55169),
            .I(N__55010));
    InMux I__13009 (
            .O(N__55168),
            .I(N__55010));
    InMux I__13008 (
            .O(N__55167),
            .I(N__55010));
    InMux I__13007 (
            .O(N__55166),
            .I(N__55010));
    InMux I__13006 (
            .O(N__55165),
            .I(N__55001));
    InMux I__13005 (
            .O(N__55164),
            .I(N__55001));
    InMux I__13004 (
            .O(N__55163),
            .I(N__55001));
    InMux I__13003 (
            .O(N__55162),
            .I(N__55001));
    CascadeMux I__13002 (
            .O(N__55161),
            .I(N__54998));
    LocalMux I__13001 (
            .O(N__55156),
            .I(N__54968));
    LocalMux I__13000 (
            .O(N__55153),
            .I(N__54968));
    LocalMux I__12999 (
            .O(N__55146),
            .I(N__54968));
    InMux I__12998 (
            .O(N__55145),
            .I(N__54959));
    InMux I__12997 (
            .O(N__55142),
            .I(N__54959));
    InMux I__12996 (
            .O(N__55141),
            .I(N__54959));
    InMux I__12995 (
            .O(N__55140),
            .I(N__54959));
    InMux I__12994 (
            .O(N__55137),
            .I(N__54952));
    InMux I__12993 (
            .O(N__55136),
            .I(N__54952));
    InMux I__12992 (
            .O(N__55135),
            .I(N__54952));
    CascadeMux I__12991 (
            .O(N__55134),
            .I(N__54942));
    CascadeMux I__12990 (
            .O(N__55133),
            .I(N__54931));
    CascadeMux I__12989 (
            .O(N__55132),
            .I(N__54928));
    CascadeMux I__12988 (
            .O(N__55131),
            .I(N__54917));
    CascadeMux I__12987 (
            .O(N__55130),
            .I(N__54914));
    CascadeMux I__12986 (
            .O(N__55129),
            .I(N__54911));
    CascadeMux I__12985 (
            .O(N__55128),
            .I(N__54908));
    CascadeMux I__12984 (
            .O(N__55127),
            .I(N__54905));
    CascadeMux I__12983 (
            .O(N__55126),
            .I(N__54902));
    CascadeMux I__12982 (
            .O(N__55125),
            .I(N__54899));
    CascadeMux I__12981 (
            .O(N__55124),
            .I(N__54896));
    CascadeMux I__12980 (
            .O(N__55123),
            .I(N__54893));
    CascadeMux I__12979 (
            .O(N__55122),
            .I(N__54890));
    InMux I__12978 (
            .O(N__55121),
            .I(N__54848));
    InMux I__12977 (
            .O(N__55118),
            .I(N__54848));
    InMux I__12976 (
            .O(N__55117),
            .I(N__54848));
    InMux I__12975 (
            .O(N__55114),
            .I(N__54848));
    InMux I__12974 (
            .O(N__55113),
            .I(N__54848));
    InMux I__12973 (
            .O(N__55110),
            .I(N__54848));
    InMux I__12972 (
            .O(N__55109),
            .I(N__54848));
    InMux I__12971 (
            .O(N__55106),
            .I(N__54848));
    InMux I__12970 (
            .O(N__55103),
            .I(N__54831));
    InMux I__12969 (
            .O(N__55102),
            .I(N__54831));
    InMux I__12968 (
            .O(N__55099),
            .I(N__54831));
    InMux I__12967 (
            .O(N__55098),
            .I(N__54831));
    InMux I__12966 (
            .O(N__55095),
            .I(N__54831));
    InMux I__12965 (
            .O(N__55094),
            .I(N__54831));
    InMux I__12964 (
            .O(N__55091),
            .I(N__54831));
    InMux I__12963 (
            .O(N__55090),
            .I(N__54831));
    CascadeMux I__12962 (
            .O(N__55089),
            .I(N__54828));
    CascadeMux I__12961 (
            .O(N__55088),
            .I(N__54824));
    CascadeMux I__12960 (
            .O(N__55087),
            .I(N__54820));
    CascadeMux I__12959 (
            .O(N__55086),
            .I(N__54816));
    CascadeMux I__12958 (
            .O(N__55085),
            .I(N__54812));
    CascadeMux I__12957 (
            .O(N__55084),
            .I(N__54809));
    CascadeMux I__12956 (
            .O(N__55083),
            .I(N__54806));
    CascadeMux I__12955 (
            .O(N__55082),
            .I(N__54803));
    CascadeMux I__12954 (
            .O(N__55081),
            .I(N__54800));
    CascadeMux I__12953 (
            .O(N__55080),
            .I(N__54797));
    CascadeMux I__12952 (
            .O(N__55079),
            .I(N__54794));
    CascadeMux I__12951 (
            .O(N__55078),
            .I(N__54791));
    CascadeMux I__12950 (
            .O(N__55077),
            .I(N__54788));
    CascadeMux I__12949 (
            .O(N__55076),
            .I(N__54785));
    InMux I__12948 (
            .O(N__55073),
            .I(N__54779));
    InMux I__12947 (
            .O(N__55072),
            .I(N__54779));
    InMux I__12946 (
            .O(N__55071),
            .I(N__54774));
    InMux I__12945 (
            .O(N__55070),
            .I(N__54774));
    InMux I__12944 (
            .O(N__55069),
            .I(N__54762));
    InMux I__12943 (
            .O(N__55068),
            .I(N__54762));
    InMux I__12942 (
            .O(N__55067),
            .I(N__54759));
    InMux I__12941 (
            .O(N__55066),
            .I(N__54756));
    InMux I__12940 (
            .O(N__55065),
            .I(N__54749));
    InMux I__12939 (
            .O(N__55064),
            .I(N__54749));
    InMux I__12938 (
            .O(N__55063),
            .I(N__54749));
    CascadeMux I__12937 (
            .O(N__55062),
            .I(N__54745));
    CascadeMux I__12936 (
            .O(N__55061),
            .I(N__54735));
    InMux I__12935 (
            .O(N__55060),
            .I(N__54724));
    Span4Mux_v I__12934 (
            .O(N__55057),
            .I(N__54717));
    Span4Mux_h I__12933 (
            .O(N__55054),
            .I(N__54717));
    LocalMux I__12932 (
            .O(N__55047),
            .I(N__54717));
    InMux I__12931 (
            .O(N__55044),
            .I(N__54712));
    InMux I__12930 (
            .O(N__55041),
            .I(N__54712));
    InMux I__12929 (
            .O(N__55038),
            .I(N__54703));
    InMux I__12928 (
            .O(N__55035),
            .I(N__54703));
    InMux I__12927 (
            .O(N__55034),
            .I(N__54703));
    InMux I__12926 (
            .O(N__55031),
            .I(N__54703));
    Span4Mux_s3_v I__12925 (
            .O(N__55026),
            .I(N__54694));
    LocalMux I__12924 (
            .O(N__55019),
            .I(N__54694));
    LocalMux I__12923 (
            .O(N__55010),
            .I(N__54689));
    LocalMux I__12922 (
            .O(N__55001),
            .I(N__54689));
    InMux I__12921 (
            .O(N__54998),
            .I(N__54686));
    CascadeMux I__12920 (
            .O(N__54997),
            .I(N__54683));
    CascadeMux I__12919 (
            .O(N__54996),
            .I(N__54680));
    CascadeMux I__12918 (
            .O(N__54995),
            .I(N__54673));
    CascadeMux I__12917 (
            .O(N__54994),
            .I(N__54670));
    CascadeMux I__12916 (
            .O(N__54993),
            .I(N__54665));
    CascadeMux I__12915 (
            .O(N__54992),
            .I(N__54662));
    CascadeMux I__12914 (
            .O(N__54991),
            .I(N__54659));
    CascadeMux I__12913 (
            .O(N__54990),
            .I(N__54656));
    CascadeMux I__12912 (
            .O(N__54989),
            .I(N__54653));
    CascadeMux I__12911 (
            .O(N__54988),
            .I(N__54650));
    CascadeMux I__12910 (
            .O(N__54987),
            .I(N__54646));
    CascadeMux I__12909 (
            .O(N__54986),
            .I(N__54643));
    CascadeMux I__12908 (
            .O(N__54985),
            .I(N__54640));
    CascadeMux I__12907 (
            .O(N__54984),
            .I(N__54637));
    CascadeMux I__12906 (
            .O(N__54983),
            .I(N__54634));
    CascadeMux I__12905 (
            .O(N__54982),
            .I(N__54631));
    CascadeMux I__12904 (
            .O(N__54981),
            .I(N__54628));
    CascadeMux I__12903 (
            .O(N__54980),
            .I(N__54625));
    CascadeMux I__12902 (
            .O(N__54979),
            .I(N__54622));
    CascadeMux I__12901 (
            .O(N__54978),
            .I(N__54606));
    CascadeMux I__12900 (
            .O(N__54977),
            .I(N__54600));
    CascadeMux I__12899 (
            .O(N__54976),
            .I(N__54590));
    CascadeMux I__12898 (
            .O(N__54975),
            .I(N__54586));
    Span4Mux_s2_v I__12897 (
            .O(N__54968),
            .I(N__54573));
    LocalMux I__12896 (
            .O(N__54959),
            .I(N__54573));
    LocalMux I__12895 (
            .O(N__54952),
            .I(N__54573));
    InMux I__12894 (
            .O(N__54951),
            .I(N__54570));
    InMux I__12893 (
            .O(N__54950),
            .I(N__54567));
    InMux I__12892 (
            .O(N__54949),
            .I(N__54560));
    InMux I__12891 (
            .O(N__54948),
            .I(N__54560));
    InMux I__12890 (
            .O(N__54947),
            .I(N__54560));
    InMux I__12889 (
            .O(N__54946),
            .I(N__54549));
    InMux I__12888 (
            .O(N__54945),
            .I(N__54549));
    InMux I__12887 (
            .O(N__54942),
            .I(N__54549));
    InMux I__12886 (
            .O(N__54941),
            .I(N__54549));
    InMux I__12885 (
            .O(N__54940),
            .I(N__54549));
    InMux I__12884 (
            .O(N__54939),
            .I(N__54546));
    InMux I__12883 (
            .O(N__54938),
            .I(N__54539));
    InMux I__12882 (
            .O(N__54937),
            .I(N__54539));
    InMux I__12881 (
            .O(N__54936),
            .I(N__54539));
    CascadeMux I__12880 (
            .O(N__54935),
            .I(N__54536));
    CascadeMux I__12879 (
            .O(N__54934),
            .I(N__54532));
    InMux I__12878 (
            .O(N__54931),
            .I(N__54522));
    InMux I__12877 (
            .O(N__54928),
            .I(N__54522));
    InMux I__12876 (
            .O(N__54927),
            .I(N__54522));
    InMux I__12875 (
            .O(N__54926),
            .I(N__54522));
    CascadeMux I__12874 (
            .O(N__54925),
            .I(N__54514));
    CascadeMux I__12873 (
            .O(N__54924),
            .I(N__54511));
    CascadeMux I__12872 (
            .O(N__54923),
            .I(N__54506));
    CascadeMux I__12871 (
            .O(N__54922),
            .I(N__54502));
    CascadeMux I__12870 (
            .O(N__54921),
            .I(N__54498));
    CascadeMux I__12869 (
            .O(N__54920),
            .I(N__54495));
    InMux I__12868 (
            .O(N__54917),
            .I(N__54488));
    InMux I__12867 (
            .O(N__54914),
            .I(N__54488));
    InMux I__12866 (
            .O(N__54911),
            .I(N__54488));
    InMux I__12865 (
            .O(N__54908),
            .I(N__54479));
    InMux I__12864 (
            .O(N__54905),
            .I(N__54479));
    InMux I__12863 (
            .O(N__54902),
            .I(N__54479));
    InMux I__12862 (
            .O(N__54899),
            .I(N__54479));
    InMux I__12861 (
            .O(N__54896),
            .I(N__54472));
    InMux I__12860 (
            .O(N__54893),
            .I(N__54472));
    InMux I__12859 (
            .O(N__54890),
            .I(N__54472));
    CascadeMux I__12858 (
            .O(N__54889),
            .I(N__54468));
    CascadeMux I__12857 (
            .O(N__54888),
            .I(N__54465));
    CascadeMux I__12856 (
            .O(N__54887),
            .I(N__54462));
    CascadeMux I__12855 (
            .O(N__54886),
            .I(N__54459));
    CascadeMux I__12854 (
            .O(N__54885),
            .I(N__54456));
    CascadeMux I__12853 (
            .O(N__54884),
            .I(N__54453));
    CascadeMux I__12852 (
            .O(N__54883),
            .I(N__54450));
    CascadeMux I__12851 (
            .O(N__54882),
            .I(N__54447));
    CascadeMux I__12850 (
            .O(N__54881),
            .I(N__54444));
    CascadeMux I__12849 (
            .O(N__54880),
            .I(N__54441));
    CascadeMux I__12848 (
            .O(N__54879),
            .I(N__54438));
    CascadeMux I__12847 (
            .O(N__54878),
            .I(N__54435));
    CascadeMux I__12846 (
            .O(N__54877),
            .I(N__54432));
    CascadeMux I__12845 (
            .O(N__54876),
            .I(N__54428));
    CascadeMux I__12844 (
            .O(N__54875),
            .I(N__54425));
    CascadeMux I__12843 (
            .O(N__54874),
            .I(N__54422));
    CascadeMux I__12842 (
            .O(N__54873),
            .I(N__54419));
    CascadeMux I__12841 (
            .O(N__54872),
            .I(N__54416));
    CascadeMux I__12840 (
            .O(N__54871),
            .I(N__54413));
    CascadeMux I__12839 (
            .O(N__54870),
            .I(N__54410));
    CascadeMux I__12838 (
            .O(N__54869),
            .I(N__54407));
    CascadeMux I__12837 (
            .O(N__54868),
            .I(N__54404));
    CascadeMux I__12836 (
            .O(N__54867),
            .I(N__54400));
    CascadeMux I__12835 (
            .O(N__54866),
            .I(N__54397));
    CascadeMux I__12834 (
            .O(N__54865),
            .I(N__54394));
    LocalMux I__12833 (
            .O(N__54848),
            .I(N__54389));
    LocalMux I__12832 (
            .O(N__54831),
            .I(N__54389));
    InMux I__12831 (
            .O(N__54828),
            .I(N__54374));
    InMux I__12830 (
            .O(N__54827),
            .I(N__54374));
    InMux I__12829 (
            .O(N__54824),
            .I(N__54374));
    InMux I__12828 (
            .O(N__54823),
            .I(N__54374));
    InMux I__12827 (
            .O(N__54820),
            .I(N__54374));
    InMux I__12826 (
            .O(N__54819),
            .I(N__54374));
    InMux I__12825 (
            .O(N__54816),
            .I(N__54374));
    InMux I__12824 (
            .O(N__54815),
            .I(N__54367));
    InMux I__12823 (
            .O(N__54812),
            .I(N__54367));
    InMux I__12822 (
            .O(N__54809),
            .I(N__54367));
    InMux I__12821 (
            .O(N__54806),
            .I(N__54358));
    InMux I__12820 (
            .O(N__54803),
            .I(N__54358));
    InMux I__12819 (
            .O(N__54800),
            .I(N__54358));
    InMux I__12818 (
            .O(N__54797),
            .I(N__54358));
    InMux I__12817 (
            .O(N__54794),
            .I(N__54347));
    InMux I__12816 (
            .O(N__54791),
            .I(N__54347));
    InMux I__12815 (
            .O(N__54788),
            .I(N__54347));
    InMux I__12814 (
            .O(N__54785),
            .I(N__54347));
    InMux I__12813 (
            .O(N__54784),
            .I(N__54347));
    LocalMux I__12812 (
            .O(N__54779),
            .I(N__54331));
    LocalMux I__12811 (
            .O(N__54774),
            .I(N__54331));
    InMux I__12810 (
            .O(N__54773),
            .I(N__54324));
    InMux I__12809 (
            .O(N__54772),
            .I(N__54324));
    InMux I__12808 (
            .O(N__54771),
            .I(N__54324));
    CascadeMux I__12807 (
            .O(N__54770),
            .I(N__54318));
    CascadeMux I__12806 (
            .O(N__54769),
            .I(N__54315));
    CascadeMux I__12805 (
            .O(N__54768),
            .I(N__54312));
    CascadeMux I__12804 (
            .O(N__54767),
            .I(N__54309));
    LocalMux I__12803 (
            .O(N__54762),
            .I(N__54299));
    LocalMux I__12802 (
            .O(N__54759),
            .I(N__54299));
    LocalMux I__12801 (
            .O(N__54756),
            .I(N__54299));
    LocalMux I__12800 (
            .O(N__54749),
            .I(N__54299));
    InMux I__12799 (
            .O(N__54748),
            .I(N__54292));
    InMux I__12798 (
            .O(N__54745),
            .I(N__54292));
    InMux I__12797 (
            .O(N__54744),
            .I(N__54292));
    InMux I__12796 (
            .O(N__54743),
            .I(N__54287));
    InMux I__12795 (
            .O(N__54742),
            .I(N__54287));
    InMux I__12794 (
            .O(N__54741),
            .I(N__54284));
    InMux I__12793 (
            .O(N__54740),
            .I(N__54277));
    InMux I__12792 (
            .O(N__54739),
            .I(N__54277));
    InMux I__12791 (
            .O(N__54738),
            .I(N__54277));
    InMux I__12790 (
            .O(N__54735),
            .I(N__54272));
    InMux I__12789 (
            .O(N__54734),
            .I(N__54272));
    InMux I__12788 (
            .O(N__54733),
            .I(N__54267));
    InMux I__12787 (
            .O(N__54732),
            .I(N__54267));
    CascadeMux I__12786 (
            .O(N__54731),
            .I(N__54263));
    CascadeMux I__12785 (
            .O(N__54730),
            .I(N__54260));
    CascadeMux I__12784 (
            .O(N__54729),
            .I(N__54257));
    CascadeMux I__12783 (
            .O(N__54728),
            .I(N__54245));
    CascadeMux I__12782 (
            .O(N__54727),
            .I(N__54242));
    LocalMux I__12781 (
            .O(N__54724),
            .I(N__54235));
    Span4Mux_v I__12780 (
            .O(N__54717),
            .I(N__54235));
    LocalMux I__12779 (
            .O(N__54712),
            .I(N__54230));
    LocalMux I__12778 (
            .O(N__54703),
            .I(N__54230));
    InMux I__12777 (
            .O(N__54702),
            .I(N__54227));
    InMux I__12776 (
            .O(N__54701),
            .I(N__54220));
    InMux I__12775 (
            .O(N__54700),
            .I(N__54220));
    InMux I__12774 (
            .O(N__54699),
            .I(N__54220));
    Span4Mux_v I__12773 (
            .O(N__54694),
            .I(N__54213));
    Span4Mux_h I__12772 (
            .O(N__54689),
            .I(N__54213));
    LocalMux I__12771 (
            .O(N__54686),
            .I(N__54213));
    InMux I__12770 (
            .O(N__54683),
            .I(N__54204));
    InMux I__12769 (
            .O(N__54680),
            .I(N__54204));
    InMux I__12768 (
            .O(N__54679),
            .I(N__54204));
    InMux I__12767 (
            .O(N__54678),
            .I(N__54204));
    CascadeMux I__12766 (
            .O(N__54677),
            .I(N__54201));
    CascadeMux I__12765 (
            .O(N__54676),
            .I(N__54198));
    InMux I__12764 (
            .O(N__54673),
            .I(N__54191));
    InMux I__12763 (
            .O(N__54670),
            .I(N__54191));
    InMux I__12762 (
            .O(N__54669),
            .I(N__54191));
    InMux I__12761 (
            .O(N__54668),
            .I(N__54186));
    InMux I__12760 (
            .O(N__54665),
            .I(N__54186));
    InMux I__12759 (
            .O(N__54662),
            .I(N__54183));
    InMux I__12758 (
            .O(N__54659),
            .I(N__54172));
    InMux I__12757 (
            .O(N__54656),
            .I(N__54172));
    InMux I__12756 (
            .O(N__54653),
            .I(N__54172));
    InMux I__12755 (
            .O(N__54650),
            .I(N__54172));
    InMux I__12754 (
            .O(N__54649),
            .I(N__54172));
    InMux I__12753 (
            .O(N__54646),
            .I(N__54163));
    InMux I__12752 (
            .O(N__54643),
            .I(N__54163));
    InMux I__12751 (
            .O(N__54640),
            .I(N__54163));
    InMux I__12750 (
            .O(N__54637),
            .I(N__54163));
    InMux I__12749 (
            .O(N__54634),
            .I(N__54154));
    InMux I__12748 (
            .O(N__54631),
            .I(N__54154));
    InMux I__12747 (
            .O(N__54628),
            .I(N__54154));
    InMux I__12746 (
            .O(N__54625),
            .I(N__54154));
    InMux I__12745 (
            .O(N__54622),
            .I(N__54143));
    InMux I__12744 (
            .O(N__54621),
            .I(N__54143));
    InMux I__12743 (
            .O(N__54620),
            .I(N__54143));
    InMux I__12742 (
            .O(N__54619),
            .I(N__54143));
    InMux I__12741 (
            .O(N__54618),
            .I(N__54143));
    InMux I__12740 (
            .O(N__54617),
            .I(N__54134));
    InMux I__12739 (
            .O(N__54616),
            .I(N__54134));
    InMux I__12738 (
            .O(N__54615),
            .I(N__54134));
    InMux I__12737 (
            .O(N__54614),
            .I(N__54134));
    InMux I__12736 (
            .O(N__54613),
            .I(N__54131));
    InMux I__12735 (
            .O(N__54612),
            .I(N__54124));
    InMux I__12734 (
            .O(N__54611),
            .I(N__54124));
    InMux I__12733 (
            .O(N__54610),
            .I(N__54124));
    InMux I__12732 (
            .O(N__54609),
            .I(N__54119));
    InMux I__12731 (
            .O(N__54606),
            .I(N__54119));
    CascadeMux I__12730 (
            .O(N__54605),
            .I(N__54116));
    CascadeMux I__12729 (
            .O(N__54604),
            .I(N__54112));
    CascadeMux I__12728 (
            .O(N__54603),
            .I(N__54109));
    InMux I__12727 (
            .O(N__54600),
            .I(N__54106));
    InMux I__12726 (
            .O(N__54599),
            .I(N__54103));
    InMux I__12725 (
            .O(N__54598),
            .I(N__54100));
    InMux I__12724 (
            .O(N__54597),
            .I(N__54095));
    InMux I__12723 (
            .O(N__54596),
            .I(N__54095));
    InMux I__12722 (
            .O(N__54595),
            .I(N__54090));
    InMux I__12721 (
            .O(N__54594),
            .I(N__54090));
    InMux I__12720 (
            .O(N__54593),
            .I(N__54085));
    InMux I__12719 (
            .O(N__54590),
            .I(N__54085));
    CascadeMux I__12718 (
            .O(N__54589),
            .I(N__54079));
    InMux I__12717 (
            .O(N__54586),
            .I(N__54070));
    InMux I__12716 (
            .O(N__54585),
            .I(N__54070));
    InMux I__12715 (
            .O(N__54584),
            .I(N__54070));
    InMux I__12714 (
            .O(N__54583),
            .I(N__54063));
    InMux I__12713 (
            .O(N__54582),
            .I(N__54063));
    InMux I__12712 (
            .O(N__54581),
            .I(N__54063));
    InMux I__12711 (
            .O(N__54580),
            .I(N__54060));
    Span4Mux_v I__12710 (
            .O(N__54573),
            .I(N__54042));
    LocalMux I__12709 (
            .O(N__54570),
            .I(N__54042));
    LocalMux I__12708 (
            .O(N__54567),
            .I(N__54042));
    LocalMux I__12707 (
            .O(N__54560),
            .I(N__54042));
    LocalMux I__12706 (
            .O(N__54549),
            .I(N__54042));
    LocalMux I__12705 (
            .O(N__54546),
            .I(N__54042));
    LocalMux I__12704 (
            .O(N__54539),
            .I(N__54042));
    InMux I__12703 (
            .O(N__54536),
            .I(N__54039));
    InMux I__12702 (
            .O(N__54535),
            .I(N__54034));
    InMux I__12701 (
            .O(N__54532),
            .I(N__54034));
    InMux I__12700 (
            .O(N__54531),
            .I(N__54031));
    LocalMux I__12699 (
            .O(N__54522),
            .I(N__54028));
    InMux I__12698 (
            .O(N__54521),
            .I(N__54025));
    InMux I__12697 (
            .O(N__54520),
            .I(N__54018));
    InMux I__12696 (
            .O(N__54519),
            .I(N__54018));
    InMux I__12695 (
            .O(N__54518),
            .I(N__54018));
    InMux I__12694 (
            .O(N__54517),
            .I(N__54013));
    InMux I__12693 (
            .O(N__54514),
            .I(N__54013));
    InMux I__12692 (
            .O(N__54511),
            .I(N__53998));
    InMux I__12691 (
            .O(N__54510),
            .I(N__53998));
    InMux I__12690 (
            .O(N__54509),
            .I(N__53998));
    InMux I__12689 (
            .O(N__54506),
            .I(N__53998));
    InMux I__12688 (
            .O(N__54505),
            .I(N__53998));
    InMux I__12687 (
            .O(N__54502),
            .I(N__53998));
    InMux I__12686 (
            .O(N__54501),
            .I(N__53998));
    InMux I__12685 (
            .O(N__54498),
            .I(N__53993));
    InMux I__12684 (
            .O(N__54495),
            .I(N__53993));
    LocalMux I__12683 (
            .O(N__54488),
            .I(N__53983));
    LocalMux I__12682 (
            .O(N__54479),
            .I(N__53983));
    LocalMux I__12681 (
            .O(N__54472),
            .I(N__53983));
    InMux I__12680 (
            .O(N__54471),
            .I(N__53974));
    InMux I__12679 (
            .O(N__54468),
            .I(N__53974));
    InMux I__12678 (
            .O(N__54465),
            .I(N__53974));
    InMux I__12677 (
            .O(N__54462),
            .I(N__53974));
    InMux I__12676 (
            .O(N__54459),
            .I(N__53965));
    InMux I__12675 (
            .O(N__54456),
            .I(N__53965));
    InMux I__12674 (
            .O(N__54453),
            .I(N__53965));
    InMux I__12673 (
            .O(N__54450),
            .I(N__53965));
    InMux I__12672 (
            .O(N__54447),
            .I(N__53958));
    InMux I__12671 (
            .O(N__54444),
            .I(N__53958));
    InMux I__12670 (
            .O(N__54441),
            .I(N__53958));
    InMux I__12669 (
            .O(N__54438),
            .I(N__53947));
    InMux I__12668 (
            .O(N__54435),
            .I(N__53947));
    InMux I__12667 (
            .O(N__54432),
            .I(N__53947));
    InMux I__12666 (
            .O(N__54431),
            .I(N__53947));
    InMux I__12665 (
            .O(N__54428),
            .I(N__53947));
    InMux I__12664 (
            .O(N__54425),
            .I(N__53938));
    InMux I__12663 (
            .O(N__54422),
            .I(N__53938));
    InMux I__12662 (
            .O(N__54419),
            .I(N__53938));
    InMux I__12661 (
            .O(N__54416),
            .I(N__53938));
    InMux I__12660 (
            .O(N__54413),
            .I(N__53929));
    InMux I__12659 (
            .O(N__54410),
            .I(N__53929));
    InMux I__12658 (
            .O(N__54407),
            .I(N__53929));
    InMux I__12657 (
            .O(N__54404),
            .I(N__53929));
    InMux I__12656 (
            .O(N__54403),
            .I(N__53920));
    InMux I__12655 (
            .O(N__54400),
            .I(N__53920));
    InMux I__12654 (
            .O(N__54397),
            .I(N__53920));
    InMux I__12653 (
            .O(N__54394),
            .I(N__53920));
    Span4Mux_v I__12652 (
            .O(N__54389),
            .I(N__53909));
    LocalMux I__12651 (
            .O(N__54374),
            .I(N__53909));
    LocalMux I__12650 (
            .O(N__54367),
            .I(N__53909));
    LocalMux I__12649 (
            .O(N__54358),
            .I(N__53909));
    LocalMux I__12648 (
            .O(N__54347),
            .I(N__53909));
    InMux I__12647 (
            .O(N__54346),
            .I(N__53906));
    InMux I__12646 (
            .O(N__54345),
            .I(N__53899));
    InMux I__12645 (
            .O(N__54344),
            .I(N__53899));
    InMux I__12644 (
            .O(N__54343),
            .I(N__53899));
    InMux I__12643 (
            .O(N__54342),
            .I(N__53892));
    InMux I__12642 (
            .O(N__54341),
            .I(N__53892));
    InMux I__12641 (
            .O(N__54340),
            .I(N__53892));
    CascadeMux I__12640 (
            .O(N__54339),
            .I(N__53887));
    CascadeMux I__12639 (
            .O(N__54338),
            .I(N__53884));
    CascadeMux I__12638 (
            .O(N__54337),
            .I(N__53881));
    CascadeMux I__12637 (
            .O(N__54336),
            .I(N__53878));
    Span4Mux_h I__12636 (
            .O(N__54331),
            .I(N__53872));
    LocalMux I__12635 (
            .O(N__54324),
            .I(N__53872));
    CascadeMux I__12634 (
            .O(N__54323),
            .I(N__53866));
    CascadeMux I__12633 (
            .O(N__54322),
            .I(N__53862));
    CascadeMux I__12632 (
            .O(N__54321),
            .I(N__53855));
    InMux I__12631 (
            .O(N__54318),
            .I(N__53852));
    InMux I__12630 (
            .O(N__54315),
            .I(N__53845));
    InMux I__12629 (
            .O(N__54312),
            .I(N__53845));
    InMux I__12628 (
            .O(N__54309),
            .I(N__53845));
    CascadeMux I__12627 (
            .O(N__54308),
            .I(N__53842));
    Span4Mux_s3_v I__12626 (
            .O(N__54299),
            .I(N__53822));
    LocalMux I__12625 (
            .O(N__54292),
            .I(N__53822));
    LocalMux I__12624 (
            .O(N__54287),
            .I(N__53811));
    LocalMux I__12623 (
            .O(N__54284),
            .I(N__53811));
    LocalMux I__12622 (
            .O(N__54277),
            .I(N__53811));
    LocalMux I__12621 (
            .O(N__54272),
            .I(N__53811));
    LocalMux I__12620 (
            .O(N__54267),
            .I(N__53811));
    InMux I__12619 (
            .O(N__54266),
            .I(N__53808));
    InMux I__12618 (
            .O(N__54263),
            .I(N__53805));
    InMux I__12617 (
            .O(N__54260),
            .I(N__53796));
    InMux I__12616 (
            .O(N__54257),
            .I(N__53796));
    InMux I__12615 (
            .O(N__54256),
            .I(N__53796));
    InMux I__12614 (
            .O(N__54255),
            .I(N__53796));
    InMux I__12613 (
            .O(N__54254),
            .I(N__53793));
    CascadeMux I__12612 (
            .O(N__54253),
            .I(N__53786));
    CascadeMux I__12611 (
            .O(N__54252),
            .I(N__53783));
    CascadeMux I__12610 (
            .O(N__54251),
            .I(N__53780));
    CascadeMux I__12609 (
            .O(N__54250),
            .I(N__53777));
    CascadeMux I__12608 (
            .O(N__54249),
            .I(N__53774));
    CascadeMux I__12607 (
            .O(N__54248),
            .I(N__53770));
    InMux I__12606 (
            .O(N__54245),
            .I(N__53755));
    InMux I__12605 (
            .O(N__54242),
            .I(N__53755));
    InMux I__12604 (
            .O(N__54241),
            .I(N__53755));
    InMux I__12603 (
            .O(N__54240),
            .I(N__53755));
    Span4Mux_h I__12602 (
            .O(N__54235),
            .I(N__53742));
    Span4Mux_v I__12601 (
            .O(N__54230),
            .I(N__53742));
    LocalMux I__12600 (
            .O(N__54227),
            .I(N__53742));
    LocalMux I__12599 (
            .O(N__54220),
            .I(N__53742));
    Span4Mux_v I__12598 (
            .O(N__54213),
            .I(N__53742));
    LocalMux I__12597 (
            .O(N__54204),
            .I(N__53742));
    InMux I__12596 (
            .O(N__54201),
            .I(N__53737));
    InMux I__12595 (
            .O(N__54198),
            .I(N__53737));
    LocalMux I__12594 (
            .O(N__54191),
            .I(N__53719));
    LocalMux I__12593 (
            .O(N__54186),
            .I(N__53719));
    LocalMux I__12592 (
            .O(N__54183),
            .I(N__53719));
    LocalMux I__12591 (
            .O(N__54172),
            .I(N__53719));
    LocalMux I__12590 (
            .O(N__54163),
            .I(N__53719));
    LocalMux I__12589 (
            .O(N__54154),
            .I(N__53719));
    LocalMux I__12588 (
            .O(N__54143),
            .I(N__53719));
    LocalMux I__12587 (
            .O(N__54134),
            .I(N__53719));
    LocalMux I__12586 (
            .O(N__54131),
            .I(N__53714));
    LocalMux I__12585 (
            .O(N__54124),
            .I(N__53714));
    LocalMux I__12584 (
            .O(N__54119),
            .I(N__53711));
    InMux I__12583 (
            .O(N__54116),
            .I(N__53702));
    InMux I__12582 (
            .O(N__54115),
            .I(N__53702));
    InMux I__12581 (
            .O(N__54112),
            .I(N__53702));
    InMux I__12580 (
            .O(N__54109),
            .I(N__53702));
    LocalMux I__12579 (
            .O(N__54106),
            .I(N__53697));
    LocalMux I__12578 (
            .O(N__54103),
            .I(N__53697));
    LocalMux I__12577 (
            .O(N__54100),
            .I(N__53690));
    LocalMux I__12576 (
            .O(N__54095),
            .I(N__53690));
    LocalMux I__12575 (
            .O(N__54090),
            .I(N__53690));
    LocalMux I__12574 (
            .O(N__54085),
            .I(N__53687));
    InMux I__12573 (
            .O(N__54084),
            .I(N__53682));
    InMux I__12572 (
            .O(N__54083),
            .I(N__53682));
    InMux I__12571 (
            .O(N__54082),
            .I(N__53677));
    InMux I__12570 (
            .O(N__54079),
            .I(N__53677));
    CascadeMux I__12569 (
            .O(N__54078),
            .I(N__53673));
    CascadeMux I__12568 (
            .O(N__54077),
            .I(N__53669));
    LocalMux I__12567 (
            .O(N__54070),
            .I(N__53659));
    LocalMux I__12566 (
            .O(N__54063),
            .I(N__53654));
    LocalMux I__12565 (
            .O(N__54060),
            .I(N__53654));
    InMux I__12564 (
            .O(N__54059),
            .I(N__53647));
    InMux I__12563 (
            .O(N__54058),
            .I(N__53647));
    InMux I__12562 (
            .O(N__54057),
            .I(N__53647));
    Span4Mux_v I__12561 (
            .O(N__54042),
            .I(N__53630));
    LocalMux I__12560 (
            .O(N__54039),
            .I(N__53630));
    LocalMux I__12559 (
            .O(N__54034),
            .I(N__53630));
    LocalMux I__12558 (
            .O(N__54031),
            .I(N__53630));
    Span4Mux_h I__12557 (
            .O(N__54028),
            .I(N__53630));
    LocalMux I__12556 (
            .O(N__54025),
            .I(N__53630));
    LocalMux I__12555 (
            .O(N__54018),
            .I(N__53630));
    LocalMux I__12554 (
            .O(N__54013),
            .I(N__53630));
    LocalMux I__12553 (
            .O(N__53998),
            .I(N__53625));
    LocalMux I__12552 (
            .O(N__53993),
            .I(N__53625));
    CascadeMux I__12551 (
            .O(N__53992),
            .I(N__53622));
    CascadeMux I__12550 (
            .O(N__53991),
            .I(N__53617));
    CascadeMux I__12549 (
            .O(N__53990),
            .I(N__53612));
    Span4Mux_v I__12548 (
            .O(N__53983),
            .I(N__53608));
    LocalMux I__12547 (
            .O(N__53974),
            .I(N__53593));
    LocalMux I__12546 (
            .O(N__53965),
            .I(N__53593));
    LocalMux I__12545 (
            .O(N__53958),
            .I(N__53593));
    LocalMux I__12544 (
            .O(N__53947),
            .I(N__53593));
    LocalMux I__12543 (
            .O(N__53938),
            .I(N__53593));
    LocalMux I__12542 (
            .O(N__53929),
            .I(N__53593));
    LocalMux I__12541 (
            .O(N__53920),
            .I(N__53593));
    Span4Mux_v I__12540 (
            .O(N__53909),
            .I(N__53584));
    LocalMux I__12539 (
            .O(N__53906),
            .I(N__53584));
    LocalMux I__12538 (
            .O(N__53899),
            .I(N__53584));
    LocalMux I__12537 (
            .O(N__53892),
            .I(N__53584));
    InMux I__12536 (
            .O(N__53891),
            .I(N__53581));
    InMux I__12535 (
            .O(N__53890),
            .I(N__53570));
    InMux I__12534 (
            .O(N__53887),
            .I(N__53570));
    InMux I__12533 (
            .O(N__53884),
            .I(N__53570));
    InMux I__12532 (
            .O(N__53881),
            .I(N__53570));
    InMux I__12531 (
            .O(N__53878),
            .I(N__53570));
    CascadeMux I__12530 (
            .O(N__53877),
            .I(N__53566));
    Span4Mux_v I__12529 (
            .O(N__53872),
            .I(N__53557));
    CascadeMux I__12528 (
            .O(N__53871),
            .I(N__53554));
    CascadeMux I__12527 (
            .O(N__53870),
            .I(N__53551));
    CascadeMux I__12526 (
            .O(N__53869),
            .I(N__53547));
    InMux I__12525 (
            .O(N__53866),
            .I(N__53536));
    InMux I__12524 (
            .O(N__53865),
            .I(N__53536));
    InMux I__12523 (
            .O(N__53862),
            .I(N__53536));
    InMux I__12522 (
            .O(N__53861),
            .I(N__53536));
    InMux I__12521 (
            .O(N__53860),
            .I(N__53536));
    InMux I__12520 (
            .O(N__53859),
            .I(N__53529));
    InMux I__12519 (
            .O(N__53858),
            .I(N__53529));
    InMux I__12518 (
            .O(N__53855),
            .I(N__53529));
    LocalMux I__12517 (
            .O(N__53852),
            .I(N__53524));
    LocalMux I__12516 (
            .O(N__53845),
            .I(N__53524));
    InMux I__12515 (
            .O(N__53842),
            .I(N__53514));
    InMux I__12514 (
            .O(N__53841),
            .I(N__53514));
    InMux I__12513 (
            .O(N__53840),
            .I(N__53514));
    InMux I__12512 (
            .O(N__53839),
            .I(N__53514));
    CascadeMux I__12511 (
            .O(N__53838),
            .I(N__53511));
    CascadeMux I__12510 (
            .O(N__53837),
            .I(N__53507));
    CascadeMux I__12509 (
            .O(N__53836),
            .I(N__53504));
    CascadeMux I__12508 (
            .O(N__53835),
            .I(N__53501));
    CascadeMux I__12507 (
            .O(N__53834),
            .I(N__53497));
    CascadeMux I__12506 (
            .O(N__53833),
            .I(N__53493));
    CascadeMux I__12505 (
            .O(N__53832),
            .I(N__53490));
    CascadeMux I__12504 (
            .O(N__53831),
            .I(N__53486));
    InMux I__12503 (
            .O(N__53830),
            .I(N__53479));
    InMux I__12502 (
            .O(N__53829),
            .I(N__53472));
    InMux I__12501 (
            .O(N__53828),
            .I(N__53472));
    InMux I__12500 (
            .O(N__53827),
            .I(N__53472));
    Span4Mux_v I__12499 (
            .O(N__53822),
            .I(N__53461));
    Span4Mux_v I__12498 (
            .O(N__53811),
            .I(N__53461));
    LocalMux I__12497 (
            .O(N__53808),
            .I(N__53461));
    LocalMux I__12496 (
            .O(N__53805),
            .I(N__53461));
    LocalMux I__12495 (
            .O(N__53796),
            .I(N__53461));
    LocalMux I__12494 (
            .O(N__53793),
            .I(N__53458));
    InMux I__12493 (
            .O(N__53792),
            .I(N__53451));
    InMux I__12492 (
            .O(N__53791),
            .I(N__53451));
    InMux I__12491 (
            .O(N__53790),
            .I(N__53451));
    InMux I__12490 (
            .O(N__53789),
            .I(N__53444));
    InMux I__12489 (
            .O(N__53786),
            .I(N__53444));
    InMux I__12488 (
            .O(N__53783),
            .I(N__53444));
    InMux I__12487 (
            .O(N__53780),
            .I(N__53437));
    InMux I__12486 (
            .O(N__53777),
            .I(N__53437));
    InMux I__12485 (
            .O(N__53774),
            .I(N__53437));
    InMux I__12484 (
            .O(N__53773),
            .I(N__53426));
    InMux I__12483 (
            .O(N__53770),
            .I(N__53426));
    InMux I__12482 (
            .O(N__53769),
            .I(N__53426));
    InMux I__12481 (
            .O(N__53768),
            .I(N__53426));
    InMux I__12480 (
            .O(N__53767),
            .I(N__53426));
    InMux I__12479 (
            .O(N__53766),
            .I(N__53419));
    InMux I__12478 (
            .O(N__53765),
            .I(N__53419));
    InMux I__12477 (
            .O(N__53764),
            .I(N__53419));
    LocalMux I__12476 (
            .O(N__53755),
            .I(N__53408));
    Span4Mux_h I__12475 (
            .O(N__53742),
            .I(N__53408));
    LocalMux I__12474 (
            .O(N__53737),
            .I(N__53408));
    InMux I__12473 (
            .O(N__53736),
            .I(N__53405));
    Span4Mux_v I__12472 (
            .O(N__53719),
            .I(N__53400));
    Span4Mux_h I__12471 (
            .O(N__53714),
            .I(N__53400));
    Span4Mux_h I__12470 (
            .O(N__53711),
            .I(N__53395));
    LocalMux I__12469 (
            .O(N__53702),
            .I(N__53395));
    Span4Mux_h I__12468 (
            .O(N__53697),
            .I(N__53388));
    Span4Mux_v I__12467 (
            .O(N__53690),
            .I(N__53388));
    Span4Mux_h I__12466 (
            .O(N__53687),
            .I(N__53388));
    LocalMux I__12465 (
            .O(N__53682),
            .I(N__53383));
    LocalMux I__12464 (
            .O(N__53677),
            .I(N__53383));
    InMux I__12463 (
            .O(N__53676),
            .I(N__53374));
    InMux I__12462 (
            .O(N__53673),
            .I(N__53374));
    InMux I__12461 (
            .O(N__53672),
            .I(N__53374));
    InMux I__12460 (
            .O(N__53669),
            .I(N__53374));
    CascadeMux I__12459 (
            .O(N__53668),
            .I(N__53370));
    CascadeMux I__12458 (
            .O(N__53667),
            .I(N__53367));
    CascadeMux I__12457 (
            .O(N__53666),
            .I(N__53363));
    CascadeMux I__12456 (
            .O(N__53665),
            .I(N__53353));
    CascadeMux I__12455 (
            .O(N__53664),
            .I(N__53344));
    CascadeMux I__12454 (
            .O(N__53663),
            .I(N__53341));
    CascadeMux I__12453 (
            .O(N__53662),
            .I(N__53337));
    Span4Mux_v I__12452 (
            .O(N__53659),
            .I(N__53330));
    Span4Mux_h I__12451 (
            .O(N__53654),
            .I(N__53330));
    LocalMux I__12450 (
            .O(N__53647),
            .I(N__53330));
    Span4Mux_v I__12449 (
            .O(N__53630),
            .I(N__53325));
    Span4Mux_v I__12448 (
            .O(N__53625),
            .I(N__53325));
    InMux I__12447 (
            .O(N__53622),
            .I(N__53318));
    InMux I__12446 (
            .O(N__53621),
            .I(N__53318));
    InMux I__12445 (
            .O(N__53620),
            .I(N__53318));
    InMux I__12444 (
            .O(N__53617),
            .I(N__53307));
    InMux I__12443 (
            .O(N__53616),
            .I(N__53307));
    InMux I__12442 (
            .O(N__53615),
            .I(N__53307));
    InMux I__12441 (
            .O(N__53612),
            .I(N__53307));
    InMux I__12440 (
            .O(N__53611),
            .I(N__53307));
    Span4Mux_h I__12439 (
            .O(N__53608),
            .I(N__53296));
    Span4Mux_v I__12438 (
            .O(N__53593),
            .I(N__53296));
    Span4Mux_h I__12437 (
            .O(N__53584),
            .I(N__53296));
    LocalMux I__12436 (
            .O(N__53581),
            .I(N__53296));
    LocalMux I__12435 (
            .O(N__53570),
            .I(N__53296));
    InMux I__12434 (
            .O(N__53569),
            .I(N__53293));
    InMux I__12433 (
            .O(N__53566),
            .I(N__53284));
    InMux I__12432 (
            .O(N__53565),
            .I(N__53284));
    InMux I__12431 (
            .O(N__53564),
            .I(N__53284));
    InMux I__12430 (
            .O(N__53563),
            .I(N__53284));
    InMux I__12429 (
            .O(N__53562),
            .I(N__53277));
    InMux I__12428 (
            .O(N__53561),
            .I(N__53277));
    InMux I__12427 (
            .O(N__53560),
            .I(N__53277));
    Span4Mux_v I__12426 (
            .O(N__53557),
            .I(N__53274));
    InMux I__12425 (
            .O(N__53554),
            .I(N__53265));
    InMux I__12424 (
            .O(N__53551),
            .I(N__53265));
    InMux I__12423 (
            .O(N__53550),
            .I(N__53265));
    InMux I__12422 (
            .O(N__53547),
            .I(N__53265));
    LocalMux I__12421 (
            .O(N__53536),
            .I(N__53258));
    LocalMux I__12420 (
            .O(N__53529),
            .I(N__53258));
    Span4Mux_v I__12419 (
            .O(N__53524),
            .I(N__53258));
    InMux I__12418 (
            .O(N__53523),
            .I(N__53255));
    LocalMux I__12417 (
            .O(N__53514),
            .I(N__53252));
    InMux I__12416 (
            .O(N__53511),
            .I(N__53243));
    InMux I__12415 (
            .O(N__53510),
            .I(N__53243));
    InMux I__12414 (
            .O(N__53507),
            .I(N__53243));
    InMux I__12413 (
            .O(N__53504),
            .I(N__53243));
    InMux I__12412 (
            .O(N__53501),
            .I(N__53232));
    InMux I__12411 (
            .O(N__53500),
            .I(N__53232));
    InMux I__12410 (
            .O(N__53497),
            .I(N__53232));
    InMux I__12409 (
            .O(N__53496),
            .I(N__53232));
    InMux I__12408 (
            .O(N__53493),
            .I(N__53232));
    InMux I__12407 (
            .O(N__53490),
            .I(N__53225));
    InMux I__12406 (
            .O(N__53489),
            .I(N__53225));
    InMux I__12405 (
            .O(N__53486),
            .I(N__53225));
    InMux I__12404 (
            .O(N__53485),
            .I(N__53222));
    InMux I__12403 (
            .O(N__53484),
            .I(N__53215));
    InMux I__12402 (
            .O(N__53483),
            .I(N__53215));
    InMux I__12401 (
            .O(N__53482),
            .I(N__53215));
    LocalMux I__12400 (
            .O(N__53479),
            .I(N__53210));
    LocalMux I__12399 (
            .O(N__53472),
            .I(N__53210));
    Span4Mux_v I__12398 (
            .O(N__53461),
            .I(N__53195));
    Span4Mux_s2_h I__12397 (
            .O(N__53458),
            .I(N__53195));
    LocalMux I__12396 (
            .O(N__53451),
            .I(N__53195));
    LocalMux I__12395 (
            .O(N__53444),
            .I(N__53195));
    LocalMux I__12394 (
            .O(N__53437),
            .I(N__53195));
    LocalMux I__12393 (
            .O(N__53426),
            .I(N__53195));
    LocalMux I__12392 (
            .O(N__53419),
            .I(N__53195));
    InMux I__12391 (
            .O(N__53418),
            .I(N__53192));
    InMux I__12390 (
            .O(N__53417),
            .I(N__53185));
    InMux I__12389 (
            .O(N__53416),
            .I(N__53185));
    InMux I__12388 (
            .O(N__53415),
            .I(N__53185));
    Span4Mux_v I__12387 (
            .O(N__53408),
            .I(N__53180));
    LocalMux I__12386 (
            .O(N__53405),
            .I(N__53180));
    Span4Mux_h I__12385 (
            .O(N__53400),
            .I(N__53172));
    Span4Mux_v I__12384 (
            .O(N__53395),
            .I(N__53172));
    Span4Mux_v I__12383 (
            .O(N__53388),
            .I(N__53165));
    Span4Mux_h I__12382 (
            .O(N__53383),
            .I(N__53165));
    LocalMux I__12381 (
            .O(N__53374),
            .I(N__53165));
    InMux I__12380 (
            .O(N__53373),
            .I(N__53154));
    InMux I__12379 (
            .O(N__53370),
            .I(N__53154));
    InMux I__12378 (
            .O(N__53367),
            .I(N__53154));
    InMux I__12377 (
            .O(N__53366),
            .I(N__53154));
    InMux I__12376 (
            .O(N__53363),
            .I(N__53154));
    InMux I__12375 (
            .O(N__53362),
            .I(N__53151));
    InMux I__12374 (
            .O(N__53361),
            .I(N__53144));
    InMux I__12373 (
            .O(N__53360),
            .I(N__53144));
    InMux I__12372 (
            .O(N__53359),
            .I(N__53144));
    InMux I__12371 (
            .O(N__53358),
            .I(N__53137));
    InMux I__12370 (
            .O(N__53357),
            .I(N__53137));
    InMux I__12369 (
            .O(N__53356),
            .I(N__53137));
    InMux I__12368 (
            .O(N__53353),
            .I(N__53126));
    InMux I__12367 (
            .O(N__53352),
            .I(N__53126));
    InMux I__12366 (
            .O(N__53351),
            .I(N__53126));
    InMux I__12365 (
            .O(N__53350),
            .I(N__53126));
    InMux I__12364 (
            .O(N__53349),
            .I(N__53126));
    CascadeMux I__12363 (
            .O(N__53348),
            .I(N__53121));
    CascadeMux I__12362 (
            .O(N__53347),
            .I(N__53118));
    InMux I__12361 (
            .O(N__53344),
            .I(N__53109));
    InMux I__12360 (
            .O(N__53341),
            .I(N__53109));
    InMux I__12359 (
            .O(N__53340),
            .I(N__53109));
    InMux I__12358 (
            .O(N__53337),
            .I(N__53109));
    Span4Mux_v I__12357 (
            .O(N__53330),
            .I(N__53105));
    Span4Mux_v I__12356 (
            .O(N__53325),
            .I(N__53098));
    LocalMux I__12355 (
            .O(N__53318),
            .I(N__53098));
    LocalMux I__12354 (
            .O(N__53307),
            .I(N__53098));
    Span4Mux_v I__12353 (
            .O(N__53296),
            .I(N__53093));
    LocalMux I__12352 (
            .O(N__53293),
            .I(N__53093));
    LocalMux I__12351 (
            .O(N__53284),
            .I(N__53088));
    LocalMux I__12350 (
            .O(N__53277),
            .I(N__53088));
    Span4Mux_h I__12349 (
            .O(N__53274),
            .I(N__53083));
    LocalMux I__12348 (
            .O(N__53265),
            .I(N__53083));
    Span4Mux_h I__12347 (
            .O(N__53258),
            .I(N__53066));
    LocalMux I__12346 (
            .O(N__53255),
            .I(N__53066));
    Span4Mux_h I__12345 (
            .O(N__53252),
            .I(N__53066));
    LocalMux I__12344 (
            .O(N__53243),
            .I(N__53066));
    LocalMux I__12343 (
            .O(N__53232),
            .I(N__53066));
    LocalMux I__12342 (
            .O(N__53225),
            .I(N__53066));
    LocalMux I__12341 (
            .O(N__53222),
            .I(N__53066));
    LocalMux I__12340 (
            .O(N__53215),
            .I(N__53066));
    Span4Mux_s2_h I__12339 (
            .O(N__53210),
            .I(N__53054));
    Span4Mux_v I__12338 (
            .O(N__53195),
            .I(N__53054));
    LocalMux I__12337 (
            .O(N__53192),
            .I(N__53054));
    LocalMux I__12336 (
            .O(N__53185),
            .I(N__53054));
    Span4Mux_v I__12335 (
            .O(N__53180),
            .I(N__53051));
    InMux I__12334 (
            .O(N__53179),
            .I(N__53044));
    InMux I__12333 (
            .O(N__53178),
            .I(N__53044));
    InMux I__12332 (
            .O(N__53177),
            .I(N__53044));
    Span4Mux_h I__12331 (
            .O(N__53172),
            .I(N__53029));
    Span4Mux_v I__12330 (
            .O(N__53165),
            .I(N__53029));
    LocalMux I__12329 (
            .O(N__53154),
            .I(N__53029));
    LocalMux I__12328 (
            .O(N__53151),
            .I(N__53029));
    LocalMux I__12327 (
            .O(N__53144),
            .I(N__53029));
    LocalMux I__12326 (
            .O(N__53137),
            .I(N__53029));
    LocalMux I__12325 (
            .O(N__53126),
            .I(N__53029));
    InMux I__12324 (
            .O(N__53125),
            .I(N__53020));
    InMux I__12323 (
            .O(N__53124),
            .I(N__53020));
    InMux I__12322 (
            .O(N__53121),
            .I(N__53020));
    InMux I__12321 (
            .O(N__53118),
            .I(N__53020));
    LocalMux I__12320 (
            .O(N__53109),
            .I(N__53017));
    CascadeMux I__12319 (
            .O(N__53108),
            .I(N__53011));
    Span4Mux_v I__12318 (
            .O(N__53105),
            .I(N__53002));
    Span4Mux_h I__12317 (
            .O(N__53098),
            .I(N__53002));
    Span4Mux_v I__12316 (
            .O(N__53093),
            .I(N__52999));
    Span4Mux_v I__12315 (
            .O(N__53088),
            .I(N__52996));
    Span4Mux_v I__12314 (
            .O(N__53083),
            .I(N__52991));
    Span4Mux_v I__12313 (
            .O(N__53066),
            .I(N__52991));
    InMux I__12312 (
            .O(N__53065),
            .I(N__52986));
    InMux I__12311 (
            .O(N__53064),
            .I(N__52986));
    CascadeMux I__12310 (
            .O(N__53063),
            .I(N__52982));
    Span4Mux_h I__12309 (
            .O(N__53054),
            .I(N__52975));
    Span4Mux_h I__12308 (
            .O(N__53051),
            .I(N__52975));
    LocalMux I__12307 (
            .O(N__53044),
            .I(N__52975));
    Span4Mux_v I__12306 (
            .O(N__53029),
            .I(N__52968));
    LocalMux I__12305 (
            .O(N__53020),
            .I(N__52968));
    Span4Mux_h I__12304 (
            .O(N__53017),
            .I(N__52968));
    InMux I__12303 (
            .O(N__53016),
            .I(N__52961));
    InMux I__12302 (
            .O(N__53015),
            .I(N__52961));
    InMux I__12301 (
            .O(N__53014),
            .I(N__52961));
    InMux I__12300 (
            .O(N__53011),
            .I(N__52950));
    InMux I__12299 (
            .O(N__53010),
            .I(N__52950));
    InMux I__12298 (
            .O(N__53009),
            .I(N__52950));
    InMux I__12297 (
            .O(N__53008),
            .I(N__52950));
    InMux I__12296 (
            .O(N__53007),
            .I(N__52950));
    Span4Mux_v I__12295 (
            .O(N__53002),
            .I(N__52939));
    Span4Mux_h I__12294 (
            .O(N__52999),
            .I(N__52939));
    Span4Mux_h I__12293 (
            .O(N__52996),
            .I(N__52939));
    Span4Mux_v I__12292 (
            .O(N__52991),
            .I(N__52939));
    LocalMux I__12291 (
            .O(N__52986),
            .I(N__52939));
    InMux I__12290 (
            .O(N__52985),
            .I(N__52934));
    InMux I__12289 (
            .O(N__52982),
            .I(N__52934));
    Odrv4 I__12288 (
            .O(N__52975),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12287 (
            .O(N__52968),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12286 (
            .O(N__52961),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12285 (
            .O(N__52950),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12284 (
            .O(N__52939),
            .I(CONSTANT_ONE_NET));
    LocalMux I__12283 (
            .O(N__52934),
            .I(CONSTANT_ONE_NET));
    InMux I__12282 (
            .O(N__52921),
            .I(n12685));
    InMux I__12281 (
            .O(N__52918),
            .I(N__52914));
    InMux I__12280 (
            .O(N__52917),
            .I(N__52910));
    LocalMux I__12279 (
            .O(N__52914),
            .I(N__52907));
    InMux I__12278 (
            .O(N__52913),
            .I(N__52904));
    LocalMux I__12277 (
            .O(N__52910),
            .I(encoder0_position_target_23));
    Odrv4 I__12276 (
            .O(N__52907),
            .I(encoder0_position_target_23));
    LocalMux I__12275 (
            .O(N__52904),
            .I(encoder0_position_target_23));
    CEMux I__12274 (
            .O(N__52897),
            .I(N__52893));
    CEMux I__12273 (
            .O(N__52896),
            .I(N__52890));
    LocalMux I__12272 (
            .O(N__52893),
            .I(N__52887));
    LocalMux I__12271 (
            .O(N__52890),
            .I(N__52884));
    Span4Mux_v I__12270 (
            .O(N__52887),
            .I(N__52876));
    Span4Mux_h I__12269 (
            .O(N__52884),
            .I(N__52876));
    SRMux I__12268 (
            .O(N__52883),
            .I(N__52873));
    SRMux I__12267 (
            .O(N__52882),
            .I(N__52870));
    CEMux I__12266 (
            .O(N__52881),
            .I(N__52866));
    Span4Mux_v I__12265 (
            .O(N__52876),
            .I(N__52860));
    LocalMux I__12264 (
            .O(N__52873),
            .I(N__52860));
    LocalMux I__12263 (
            .O(N__52870),
            .I(N__52857));
    SRMux I__12262 (
            .O(N__52869),
            .I(N__52854));
    LocalMux I__12261 (
            .O(N__52866),
            .I(N__52851));
    InMux I__12260 (
            .O(N__52865),
            .I(N__52848));
    Span4Mux_v I__12259 (
            .O(N__52860),
            .I(N__52845));
    Span4Mux_h I__12258 (
            .O(N__52857),
            .I(N__52840));
    LocalMux I__12257 (
            .O(N__52854),
            .I(N__52840));
    Span12Mux_h I__12256 (
            .O(N__52851),
            .I(N__52835));
    LocalMux I__12255 (
            .O(N__52848),
            .I(N__52835));
    Odrv4 I__12254 (
            .O(N__52845),
            .I(n4856));
    Odrv4 I__12253 (
            .O(N__52840),
            .I(n4856));
    Odrv12 I__12252 (
            .O(N__52835),
            .I(n4856));
    SRMux I__12251 (
            .O(N__52828),
            .I(N__52824));
    SRMux I__12250 (
            .O(N__52827),
            .I(N__52820));
    LocalMux I__12249 (
            .O(N__52824),
            .I(N__52817));
    SRMux I__12248 (
            .O(N__52823),
            .I(N__52814));
    LocalMux I__12247 (
            .O(N__52820),
            .I(N__52811));
    Span4Mux_v I__12246 (
            .O(N__52817),
            .I(N__52806));
    LocalMux I__12245 (
            .O(N__52814),
            .I(N__52806));
    Odrv4 I__12244 (
            .O(N__52811),
            .I(n4890));
    Odrv4 I__12243 (
            .O(N__52806),
            .I(n4890));
    InMux I__12242 (
            .O(N__52801),
            .I(N__52798));
    LocalMux I__12241 (
            .O(N__52798),
            .I(N__52795));
    Odrv12 I__12240 (
            .O(N__52795),
            .I(pwm_setpoint_23_N_171_9));
    InMux I__12239 (
            .O(N__52792),
            .I(N__52789));
    LocalMux I__12238 (
            .O(N__52789),
            .I(N__52785));
    InMux I__12237 (
            .O(N__52788),
            .I(N__52782));
    Span4Mux_h I__12236 (
            .O(N__52785),
            .I(N__52779));
    LocalMux I__12235 (
            .O(N__52782),
            .I(N__52776));
    Odrv4 I__12234 (
            .O(N__52779),
            .I(duty_9));
    Odrv12 I__12233 (
            .O(N__52776),
            .I(duty_9));
    InMux I__12232 (
            .O(N__52771),
            .I(N__52767));
    InMux I__12231 (
            .O(N__52770),
            .I(N__52764));
    LocalMux I__12230 (
            .O(N__52767),
            .I(N__52760));
    LocalMux I__12229 (
            .O(N__52764),
            .I(N__52757));
    InMux I__12228 (
            .O(N__52763),
            .I(N__52754));
    Span4Mux_h I__12227 (
            .O(N__52760),
            .I(N__52751));
    Span4Mux_s3_v I__12226 (
            .O(N__52757),
            .I(N__52748));
    LocalMux I__12225 (
            .O(N__52754),
            .I(N__52745));
    Span4Mux_h I__12224 (
            .O(N__52751),
            .I(N__52742));
    Sp12to4 I__12223 (
            .O(N__52748),
            .I(N__52737));
    Span12Mux_s3_v I__12222 (
            .O(N__52745),
            .I(N__52737));
    Odrv4 I__12221 (
            .O(N__52742),
            .I(pwm_setpoint_9));
    Odrv12 I__12220 (
            .O(N__52737),
            .I(pwm_setpoint_9));
    InMux I__12219 (
            .O(N__52732),
            .I(N__52728));
    InMux I__12218 (
            .O(N__52731),
            .I(N__52725));
    LocalMux I__12217 (
            .O(N__52728),
            .I(N__52722));
    LocalMux I__12216 (
            .O(N__52725),
            .I(N__52719));
    Span4Mux_h I__12215 (
            .O(N__52722),
            .I(N__52714));
    Span4Mux_h I__12214 (
            .O(N__52719),
            .I(N__52714));
    Odrv4 I__12213 (
            .O(N__52714),
            .I(duty_8));
    InMux I__12212 (
            .O(N__52711),
            .I(N__52708));
    LocalMux I__12211 (
            .O(N__52708),
            .I(N__52705));
    Odrv4 I__12210 (
            .O(N__52705),
            .I(n17_adj_583));
    CascadeMux I__12209 (
            .O(N__52702),
            .I(N__52698));
    InMux I__12208 (
            .O(N__52701),
            .I(N__52695));
    InMux I__12207 (
            .O(N__52698),
            .I(N__52691));
    LocalMux I__12206 (
            .O(N__52695),
            .I(N__52688));
    InMux I__12205 (
            .O(N__52694),
            .I(N__52685));
    LocalMux I__12204 (
            .O(N__52691),
            .I(encoder0_position_target_10));
    Odrv4 I__12203 (
            .O(N__52688),
            .I(encoder0_position_target_10));
    LocalMux I__12202 (
            .O(N__52685),
            .I(encoder0_position_target_10));
    InMux I__12201 (
            .O(N__52678),
            .I(n12672));
    InMux I__12200 (
            .O(N__52675),
            .I(N__52671));
    InMux I__12199 (
            .O(N__52674),
            .I(N__52667));
    LocalMux I__12198 (
            .O(N__52671),
            .I(N__52664));
    InMux I__12197 (
            .O(N__52670),
            .I(N__52661));
    LocalMux I__12196 (
            .O(N__52667),
            .I(encoder0_position_target_11));
    Odrv4 I__12195 (
            .O(N__52664),
            .I(encoder0_position_target_11));
    LocalMux I__12194 (
            .O(N__52661),
            .I(encoder0_position_target_11));
    InMux I__12193 (
            .O(N__52654),
            .I(n12673));
    CascadeMux I__12192 (
            .O(N__52651),
            .I(N__52647));
    CascadeMux I__12191 (
            .O(N__52650),
            .I(N__52644));
    InMux I__12190 (
            .O(N__52647),
            .I(N__52641));
    InMux I__12189 (
            .O(N__52644),
            .I(N__52637));
    LocalMux I__12188 (
            .O(N__52641),
            .I(N__52634));
    InMux I__12187 (
            .O(N__52640),
            .I(N__52631));
    LocalMux I__12186 (
            .O(N__52637),
            .I(encoder0_position_target_12));
    Odrv4 I__12185 (
            .O(N__52634),
            .I(encoder0_position_target_12));
    LocalMux I__12184 (
            .O(N__52631),
            .I(encoder0_position_target_12));
    InMux I__12183 (
            .O(N__52624),
            .I(n12674));
    CascadeMux I__12182 (
            .O(N__52621),
            .I(N__52618));
    InMux I__12181 (
            .O(N__52618),
            .I(N__52613));
    InMux I__12180 (
            .O(N__52617),
            .I(N__52610));
    InMux I__12179 (
            .O(N__52616),
            .I(N__52607));
    LocalMux I__12178 (
            .O(N__52613),
            .I(N__52604));
    LocalMux I__12177 (
            .O(N__52610),
            .I(N__52601));
    LocalMux I__12176 (
            .O(N__52607),
            .I(encoder0_position_target_13));
    Odrv4 I__12175 (
            .O(N__52604),
            .I(encoder0_position_target_13));
    Odrv4 I__12174 (
            .O(N__52601),
            .I(encoder0_position_target_13));
    InMux I__12173 (
            .O(N__52594),
            .I(n12675));
    InMux I__12172 (
            .O(N__52591),
            .I(N__52587));
    CascadeMux I__12171 (
            .O(N__52590),
            .I(N__52583));
    LocalMux I__12170 (
            .O(N__52587),
            .I(N__52580));
    CascadeMux I__12169 (
            .O(N__52586),
            .I(N__52577));
    InMux I__12168 (
            .O(N__52583),
            .I(N__52574));
    Span4Mux_h I__12167 (
            .O(N__52580),
            .I(N__52571));
    InMux I__12166 (
            .O(N__52577),
            .I(N__52568));
    LocalMux I__12165 (
            .O(N__52574),
            .I(encoder0_position_target_14));
    Odrv4 I__12164 (
            .O(N__52571),
            .I(encoder0_position_target_14));
    LocalMux I__12163 (
            .O(N__52568),
            .I(encoder0_position_target_14));
    InMux I__12162 (
            .O(N__52561),
            .I(n12676));
    CascadeMux I__12161 (
            .O(N__52558),
            .I(N__52555));
    InMux I__12160 (
            .O(N__52555),
            .I(N__52551));
    InMux I__12159 (
            .O(N__52554),
            .I(N__52547));
    LocalMux I__12158 (
            .O(N__52551),
            .I(N__52544));
    InMux I__12157 (
            .O(N__52550),
            .I(N__52541));
    LocalMux I__12156 (
            .O(N__52547),
            .I(encoder0_position_target_15));
    Odrv12 I__12155 (
            .O(N__52544),
            .I(encoder0_position_target_15));
    LocalMux I__12154 (
            .O(N__52541),
            .I(encoder0_position_target_15));
    InMux I__12153 (
            .O(N__52534),
            .I(n12677));
    InMux I__12152 (
            .O(N__52531),
            .I(N__52527));
    InMux I__12151 (
            .O(N__52530),
            .I(N__52523));
    LocalMux I__12150 (
            .O(N__52527),
            .I(N__52520));
    InMux I__12149 (
            .O(N__52526),
            .I(N__52517));
    LocalMux I__12148 (
            .O(N__52523),
            .I(encoder0_position_target_16));
    Odrv4 I__12147 (
            .O(N__52520),
            .I(encoder0_position_target_16));
    LocalMux I__12146 (
            .O(N__52517),
            .I(encoder0_position_target_16));
    InMux I__12145 (
            .O(N__52510),
            .I(bfn_16_28_0_));
    CascadeMux I__12144 (
            .O(N__52507),
            .I(N__52504));
    InMux I__12143 (
            .O(N__52504),
            .I(N__52500));
    CascadeMux I__12142 (
            .O(N__52503),
            .I(N__52497));
    LocalMux I__12141 (
            .O(N__52500),
            .I(N__52494));
    InMux I__12140 (
            .O(N__52497),
            .I(N__52490));
    Span4Mux_h I__12139 (
            .O(N__52494),
            .I(N__52487));
    InMux I__12138 (
            .O(N__52493),
            .I(N__52484));
    LocalMux I__12137 (
            .O(N__52490),
            .I(encoder0_position_target_17));
    Odrv4 I__12136 (
            .O(N__52487),
            .I(encoder0_position_target_17));
    LocalMux I__12135 (
            .O(N__52484),
            .I(encoder0_position_target_17));
    InMux I__12134 (
            .O(N__52477),
            .I(n12679));
    InMux I__12133 (
            .O(N__52474),
            .I(N__52471));
    LocalMux I__12132 (
            .O(N__52471),
            .I(N__52467));
    InMux I__12131 (
            .O(N__52470),
            .I(N__52463));
    Span4Mux_h I__12130 (
            .O(N__52467),
            .I(N__52460));
    InMux I__12129 (
            .O(N__52466),
            .I(N__52457));
    LocalMux I__12128 (
            .O(N__52463),
            .I(encoder0_position_target_1));
    Odrv4 I__12127 (
            .O(N__52460),
            .I(encoder0_position_target_1));
    LocalMux I__12126 (
            .O(N__52457),
            .I(encoder0_position_target_1));
    InMux I__12125 (
            .O(N__52450),
            .I(n12663));
    CascadeMux I__12124 (
            .O(N__52447),
            .I(N__52444));
    InMux I__12123 (
            .O(N__52444),
            .I(N__52440));
    CascadeMux I__12122 (
            .O(N__52443),
            .I(N__52437));
    LocalMux I__12121 (
            .O(N__52440),
            .I(N__52434));
    InMux I__12120 (
            .O(N__52437),
            .I(N__52430));
    Span4Mux_h I__12119 (
            .O(N__52434),
            .I(N__52427));
    InMux I__12118 (
            .O(N__52433),
            .I(N__52424));
    LocalMux I__12117 (
            .O(N__52430),
            .I(encoder0_position_target_2));
    Odrv4 I__12116 (
            .O(N__52427),
            .I(encoder0_position_target_2));
    LocalMux I__12115 (
            .O(N__52424),
            .I(encoder0_position_target_2));
    InMux I__12114 (
            .O(N__52417),
            .I(n12664));
    InMux I__12113 (
            .O(N__52414),
            .I(N__52411));
    LocalMux I__12112 (
            .O(N__52411),
            .I(N__52407));
    InMux I__12111 (
            .O(N__52410),
            .I(N__52403));
    Span4Mux_h I__12110 (
            .O(N__52407),
            .I(N__52400));
    InMux I__12109 (
            .O(N__52406),
            .I(N__52397));
    LocalMux I__12108 (
            .O(N__52403),
            .I(encoder0_position_target_3));
    Odrv4 I__12107 (
            .O(N__52400),
            .I(encoder0_position_target_3));
    LocalMux I__12106 (
            .O(N__52397),
            .I(encoder0_position_target_3));
    InMux I__12105 (
            .O(N__52390),
            .I(n12665));
    InMux I__12104 (
            .O(N__52387),
            .I(N__52383));
    CascadeMux I__12103 (
            .O(N__52386),
            .I(N__52380));
    LocalMux I__12102 (
            .O(N__52383),
            .I(N__52377));
    InMux I__12101 (
            .O(N__52380),
            .I(N__52373));
    Span4Mux_h I__12100 (
            .O(N__52377),
            .I(N__52370));
    InMux I__12099 (
            .O(N__52376),
            .I(N__52367));
    LocalMux I__12098 (
            .O(N__52373),
            .I(encoder0_position_target_4));
    Odrv4 I__12097 (
            .O(N__52370),
            .I(encoder0_position_target_4));
    LocalMux I__12096 (
            .O(N__52367),
            .I(encoder0_position_target_4));
    InMux I__12095 (
            .O(N__52360),
            .I(n12666));
    InMux I__12094 (
            .O(N__52357),
            .I(N__52353));
    InMux I__12093 (
            .O(N__52356),
            .I(N__52349));
    LocalMux I__12092 (
            .O(N__52353),
            .I(N__52346));
    InMux I__12091 (
            .O(N__52352),
            .I(N__52343));
    LocalMux I__12090 (
            .O(N__52349),
            .I(encoder0_position_target_5));
    Odrv4 I__12089 (
            .O(N__52346),
            .I(encoder0_position_target_5));
    LocalMux I__12088 (
            .O(N__52343),
            .I(encoder0_position_target_5));
    InMux I__12087 (
            .O(N__52336),
            .I(n12667));
    CascadeMux I__12086 (
            .O(N__52333),
            .I(N__52329));
    InMux I__12085 (
            .O(N__52332),
            .I(N__52326));
    InMux I__12084 (
            .O(N__52329),
            .I(N__52322));
    LocalMux I__12083 (
            .O(N__52326),
            .I(N__52319));
    InMux I__12082 (
            .O(N__52325),
            .I(N__52316));
    LocalMux I__12081 (
            .O(N__52322),
            .I(encoder0_position_target_6));
    Odrv4 I__12080 (
            .O(N__52319),
            .I(encoder0_position_target_6));
    LocalMux I__12079 (
            .O(N__52316),
            .I(encoder0_position_target_6));
    InMux I__12078 (
            .O(N__52309),
            .I(n12668));
    InMux I__12077 (
            .O(N__52306),
            .I(N__52302));
    InMux I__12076 (
            .O(N__52305),
            .I(N__52298));
    LocalMux I__12075 (
            .O(N__52302),
            .I(N__52295));
    InMux I__12074 (
            .O(N__52301),
            .I(N__52292));
    LocalMux I__12073 (
            .O(N__52298),
            .I(encoder0_position_target_7));
    Odrv4 I__12072 (
            .O(N__52295),
            .I(encoder0_position_target_7));
    LocalMux I__12071 (
            .O(N__52292),
            .I(encoder0_position_target_7));
    InMux I__12070 (
            .O(N__52285),
            .I(n12669));
    CascadeMux I__12069 (
            .O(N__52282),
            .I(N__52277));
    InMux I__12068 (
            .O(N__52281),
            .I(N__52274));
    CascadeMux I__12067 (
            .O(N__52280),
            .I(N__52271));
    InMux I__12066 (
            .O(N__52277),
            .I(N__52268));
    LocalMux I__12065 (
            .O(N__52274),
            .I(N__52265));
    InMux I__12064 (
            .O(N__52271),
            .I(N__52262));
    LocalMux I__12063 (
            .O(N__52268),
            .I(encoder0_position_target_8));
    Odrv4 I__12062 (
            .O(N__52265),
            .I(encoder0_position_target_8));
    LocalMux I__12061 (
            .O(N__52262),
            .I(encoder0_position_target_8));
    InMux I__12060 (
            .O(N__52255),
            .I(bfn_16_27_0_));
    InMux I__12059 (
            .O(N__52252),
            .I(N__52249));
    LocalMux I__12058 (
            .O(N__52249),
            .I(N__52245));
    InMux I__12057 (
            .O(N__52248),
            .I(N__52241));
    Span4Mux_h I__12056 (
            .O(N__52245),
            .I(N__52238));
    InMux I__12055 (
            .O(N__52244),
            .I(N__52235));
    LocalMux I__12054 (
            .O(N__52241),
            .I(encoder0_position_target_9));
    Odrv4 I__12053 (
            .O(N__52238),
            .I(encoder0_position_target_9));
    LocalMux I__12052 (
            .O(N__52235),
            .I(encoder0_position_target_9));
    InMux I__12051 (
            .O(N__52228),
            .I(n12671));
    InMux I__12050 (
            .O(N__52225),
            .I(N__52221));
    InMux I__12049 (
            .O(N__52224),
            .I(N__52218));
    LocalMux I__12048 (
            .O(N__52221),
            .I(N__52215));
    LocalMux I__12047 (
            .O(N__52218),
            .I(N__52211));
    Span4Mux_v I__12046 (
            .O(N__52215),
            .I(N__52208));
    InMux I__12045 (
            .O(N__52214),
            .I(N__52205));
    Span4Mux_v I__12044 (
            .O(N__52211),
            .I(N__52202));
    Span4Mux_h I__12043 (
            .O(N__52208),
            .I(N__52199));
    LocalMux I__12042 (
            .O(N__52205),
            .I(N__52196));
    Odrv4 I__12041 (
            .O(N__52202),
            .I(n3111));
    Odrv4 I__12040 (
            .O(N__52199),
            .I(n3111));
    Odrv12 I__12039 (
            .O(N__52196),
            .I(n3111));
    CascadeMux I__12038 (
            .O(N__52189),
            .I(N__52186));
    InMux I__12037 (
            .O(N__52186),
            .I(N__52183));
    LocalMux I__12036 (
            .O(N__52183),
            .I(N__52180));
    Odrv12 I__12035 (
            .O(N__52180),
            .I(n3178));
    InMux I__12034 (
            .O(N__52177),
            .I(n12514));
    InMux I__12033 (
            .O(N__52174),
            .I(N__52171));
    LocalMux I__12032 (
            .O(N__52171),
            .I(N__52168));
    Span4Mux_v I__12031 (
            .O(N__52168),
            .I(N__52164));
    InMux I__12030 (
            .O(N__52167),
            .I(N__52161));
    Span4Mux_h I__12029 (
            .O(N__52164),
            .I(N__52158));
    LocalMux I__12028 (
            .O(N__52161),
            .I(n3110));
    Odrv4 I__12027 (
            .O(N__52158),
            .I(n3110));
    InMux I__12026 (
            .O(N__52153),
            .I(N__52150));
    LocalMux I__12025 (
            .O(N__52150),
            .I(n3177));
    InMux I__12024 (
            .O(N__52147),
            .I(bfn_16_25_0_));
    InMux I__12023 (
            .O(N__52144),
            .I(N__52141));
    LocalMux I__12022 (
            .O(N__52141),
            .I(N__52137));
    InMux I__12021 (
            .O(N__52140),
            .I(N__52134));
    Span4Mux_v I__12020 (
            .O(N__52137),
            .I(N__52130));
    LocalMux I__12019 (
            .O(N__52134),
            .I(N__52127));
    InMux I__12018 (
            .O(N__52133),
            .I(N__52124));
    Span4Mux_h I__12017 (
            .O(N__52130),
            .I(N__52119));
    Span4Mux_v I__12016 (
            .O(N__52127),
            .I(N__52119));
    LocalMux I__12015 (
            .O(N__52124),
            .I(n3109));
    Odrv4 I__12014 (
            .O(N__52119),
            .I(n3109));
    CascadeMux I__12013 (
            .O(N__52114),
            .I(N__52111));
    InMux I__12012 (
            .O(N__52111),
            .I(N__52108));
    LocalMux I__12011 (
            .O(N__52108),
            .I(N__52105));
    Span4Mux_v I__12010 (
            .O(N__52105),
            .I(N__52102));
    Span4Mux_h I__12009 (
            .O(N__52102),
            .I(N__52099));
    Odrv4 I__12008 (
            .O(N__52099),
            .I(n3176));
    InMux I__12007 (
            .O(N__52096),
            .I(n12516));
    CascadeMux I__12006 (
            .O(N__52093),
            .I(N__52089));
    InMux I__12005 (
            .O(N__52092),
            .I(N__52086));
    InMux I__12004 (
            .O(N__52089),
            .I(N__52083));
    LocalMux I__12003 (
            .O(N__52086),
            .I(N__52078));
    LocalMux I__12002 (
            .O(N__52083),
            .I(N__52078));
    Span4Mux_h I__12001 (
            .O(N__52078),
            .I(N__52074));
    InMux I__12000 (
            .O(N__52077),
            .I(N__52071));
    Span4Mux_h I__11999 (
            .O(N__52074),
            .I(N__52068));
    LocalMux I__11998 (
            .O(N__52071),
            .I(n3108));
    Odrv4 I__11997 (
            .O(N__52068),
            .I(n3108));
    InMux I__11996 (
            .O(N__52063),
            .I(N__52060));
    LocalMux I__11995 (
            .O(N__52060),
            .I(N__52057));
    Span4Mux_h I__11994 (
            .O(N__52057),
            .I(N__52054));
    Span4Mux_h I__11993 (
            .O(N__52054),
            .I(N__52051));
    Odrv4 I__11992 (
            .O(N__52051),
            .I(n3175));
    InMux I__11991 (
            .O(N__52048),
            .I(n12517));
    InMux I__11990 (
            .O(N__52045),
            .I(N__52042));
    LocalMux I__11989 (
            .O(N__52042),
            .I(N__52037));
    InMux I__11988 (
            .O(N__52041),
            .I(N__52032));
    InMux I__11987 (
            .O(N__52040),
            .I(N__52032));
    Span4Mux_v I__11986 (
            .O(N__52037),
            .I(N__52029));
    LocalMux I__11985 (
            .O(N__52032),
            .I(N__52026));
    Span4Mux_h I__11984 (
            .O(N__52029),
            .I(N__52023));
    Span4Mux_v I__11983 (
            .O(N__52026),
            .I(N__52020));
    Odrv4 I__11982 (
            .O(N__52023),
            .I(n3107));
    Odrv4 I__11981 (
            .O(N__52020),
            .I(n3107));
    InMux I__11980 (
            .O(N__52015),
            .I(N__52012));
    LocalMux I__11979 (
            .O(N__52012),
            .I(N__52009));
    Span12Mux_h I__11978 (
            .O(N__52009),
            .I(N__52006));
    Odrv12 I__11977 (
            .O(N__52006),
            .I(n3174));
    InMux I__11976 (
            .O(N__52003),
            .I(n12518));
    InMux I__11975 (
            .O(N__52000),
            .I(N__51997));
    LocalMux I__11974 (
            .O(N__51997),
            .I(N__51993));
    InMux I__11973 (
            .O(N__51996),
            .I(N__51989));
    Span4Mux_h I__11972 (
            .O(N__51993),
            .I(N__51986));
    InMux I__11971 (
            .O(N__51992),
            .I(N__51983));
    LocalMux I__11970 (
            .O(N__51989),
            .I(N__51980));
    Span4Mux_h I__11969 (
            .O(N__51986),
            .I(N__51975));
    LocalMux I__11968 (
            .O(N__51983),
            .I(N__51975));
    Odrv4 I__11967 (
            .O(N__51980),
            .I(n3106));
    Odrv4 I__11966 (
            .O(N__51975),
            .I(n3106));
    InMux I__11965 (
            .O(N__51970),
            .I(N__51967));
    LocalMux I__11964 (
            .O(N__51967),
            .I(N__51964));
    Span4Mux_h I__11963 (
            .O(N__51964),
            .I(N__51961));
    Span4Mux_h I__11962 (
            .O(N__51961),
            .I(N__51958));
    Odrv4 I__11961 (
            .O(N__51958),
            .I(n3173));
    InMux I__11960 (
            .O(N__51955),
            .I(n12519));
    InMux I__11959 (
            .O(N__51952),
            .I(N__51948));
    InMux I__11958 (
            .O(N__51951),
            .I(N__51945));
    LocalMux I__11957 (
            .O(N__51948),
            .I(N__51942));
    LocalMux I__11956 (
            .O(N__51945),
            .I(n15158));
    Odrv12 I__11955 (
            .O(N__51942),
            .I(n15158));
    CascadeMux I__11954 (
            .O(N__51937),
            .I(N__51934));
    InMux I__11953 (
            .O(N__51934),
            .I(N__51931));
    LocalMux I__11952 (
            .O(N__51931),
            .I(N__51927));
    InMux I__11951 (
            .O(N__51930),
            .I(N__51924));
    Span4Mux_v I__11950 (
            .O(N__51927),
            .I(N__51921));
    LocalMux I__11949 (
            .O(N__51924),
            .I(N__51918));
    Odrv4 I__11948 (
            .O(N__51921),
            .I(n3105));
    Odrv12 I__11947 (
            .O(N__51918),
            .I(n3105));
    InMux I__11946 (
            .O(N__51913),
            .I(n12520));
    CascadeMux I__11945 (
            .O(N__51910),
            .I(N__51906));
    InMux I__11944 (
            .O(N__51909),
            .I(N__51903));
    InMux I__11943 (
            .O(N__51906),
            .I(N__51900));
    LocalMux I__11942 (
            .O(N__51903),
            .I(N__51897));
    LocalMux I__11941 (
            .O(N__51900),
            .I(N__51894));
    Span4Mux_h I__11940 (
            .O(N__51897),
            .I(N__51891));
    Span4Mux_v I__11939 (
            .O(N__51894),
            .I(N__51888));
    Span4Mux_h I__11938 (
            .O(N__51891),
            .I(N__51885));
    Odrv4 I__11937 (
            .O(N__51888),
            .I(n3204));
    Odrv4 I__11936 (
            .O(N__51885),
            .I(n3204));
    InMux I__11935 (
            .O(N__51880),
            .I(N__51876));
    InMux I__11934 (
            .O(N__51879),
            .I(N__51872));
    LocalMux I__11933 (
            .O(N__51876),
            .I(N__51869));
    InMux I__11932 (
            .O(N__51875),
            .I(N__51866));
    LocalMux I__11931 (
            .O(N__51872),
            .I(encoder0_position_target_0));
    Odrv4 I__11930 (
            .O(N__51869),
            .I(encoder0_position_target_0));
    LocalMux I__11929 (
            .O(N__51866),
            .I(encoder0_position_target_0));
    InMux I__11928 (
            .O(N__51859),
            .I(bfn_16_26_0_));
    InMux I__11927 (
            .O(N__51856),
            .I(N__51853));
    LocalMux I__11926 (
            .O(N__51853),
            .I(N__51849));
    InMux I__11925 (
            .O(N__51852),
            .I(N__51846));
    Span4Mux_h I__11924 (
            .O(N__51849),
            .I(N__51843));
    LocalMux I__11923 (
            .O(N__51846),
            .I(N__51839));
    Span4Mux_h I__11922 (
            .O(N__51843),
            .I(N__51836));
    InMux I__11921 (
            .O(N__51842),
            .I(N__51833));
    Odrv4 I__11920 (
            .O(N__51839),
            .I(n3118));
    Odrv4 I__11919 (
            .O(N__51836),
            .I(n3118));
    LocalMux I__11918 (
            .O(N__51833),
            .I(n3118));
    CascadeMux I__11917 (
            .O(N__51826),
            .I(N__51823));
    InMux I__11916 (
            .O(N__51823),
            .I(N__51820));
    LocalMux I__11915 (
            .O(N__51820),
            .I(N__51817));
    Span4Mux_v I__11914 (
            .O(N__51817),
            .I(N__51814));
    Span4Mux_h I__11913 (
            .O(N__51814),
            .I(N__51811));
    Odrv4 I__11912 (
            .O(N__51811),
            .I(n3185));
    InMux I__11911 (
            .O(N__51808),
            .I(bfn_16_24_0_));
    CascadeMux I__11910 (
            .O(N__51805),
            .I(N__51801));
    InMux I__11909 (
            .O(N__51804),
            .I(N__51798));
    InMux I__11908 (
            .O(N__51801),
            .I(N__51795));
    LocalMux I__11907 (
            .O(N__51798),
            .I(N__51792));
    LocalMux I__11906 (
            .O(N__51795),
            .I(N__51789));
    Span4Mux_v I__11905 (
            .O(N__51792),
            .I(N__51786));
    Span4Mux_v I__11904 (
            .O(N__51789),
            .I(N__51783));
    Span4Mux_h I__11903 (
            .O(N__51786),
            .I(N__51780));
    Odrv4 I__11902 (
            .O(N__51783),
            .I(n3117));
    Odrv4 I__11901 (
            .O(N__51780),
            .I(n3117));
    InMux I__11900 (
            .O(N__51775),
            .I(N__51772));
    LocalMux I__11899 (
            .O(N__51772),
            .I(N__51769));
    Span4Mux_v I__11898 (
            .O(N__51769),
            .I(N__51766));
    Span4Mux_h I__11897 (
            .O(N__51766),
            .I(N__51763));
    Odrv4 I__11896 (
            .O(N__51763),
            .I(n3184));
    InMux I__11895 (
            .O(N__51760),
            .I(n12508));
    InMux I__11894 (
            .O(N__51757),
            .I(N__51754));
    LocalMux I__11893 (
            .O(N__51754),
            .I(N__51751));
    Span4Mux_h I__11892 (
            .O(N__51751),
            .I(N__51746));
    InMux I__11891 (
            .O(N__51750),
            .I(N__51743));
    InMux I__11890 (
            .O(N__51749),
            .I(N__51740));
    Span4Mux_v I__11889 (
            .O(N__51746),
            .I(N__51735));
    LocalMux I__11888 (
            .O(N__51743),
            .I(N__51735));
    LocalMux I__11887 (
            .O(N__51740),
            .I(n3116));
    Odrv4 I__11886 (
            .O(N__51735),
            .I(n3116));
    InMux I__11885 (
            .O(N__51730),
            .I(N__51727));
    LocalMux I__11884 (
            .O(N__51727),
            .I(N__51724));
    Span4Mux_h I__11883 (
            .O(N__51724),
            .I(N__51721));
    Odrv4 I__11882 (
            .O(N__51721),
            .I(n3183));
    InMux I__11881 (
            .O(N__51718),
            .I(n12509));
    CascadeMux I__11880 (
            .O(N__51715),
            .I(N__51712));
    InMux I__11879 (
            .O(N__51712),
            .I(N__51708));
    InMux I__11878 (
            .O(N__51711),
            .I(N__51705));
    LocalMux I__11877 (
            .O(N__51708),
            .I(N__51702));
    LocalMux I__11876 (
            .O(N__51705),
            .I(N__51699));
    Span4Mux_v I__11875 (
            .O(N__51702),
            .I(N__51696));
    Span4Mux_v I__11874 (
            .O(N__51699),
            .I(N__51693));
    Span4Mux_v I__11873 (
            .O(N__51696),
            .I(N__51688));
    Span4Mux_h I__11872 (
            .O(N__51693),
            .I(N__51688));
    Odrv4 I__11871 (
            .O(N__51688),
            .I(n3115));
    InMux I__11870 (
            .O(N__51685),
            .I(N__51682));
    LocalMux I__11869 (
            .O(N__51682),
            .I(N__51679));
    Span4Mux_v I__11868 (
            .O(N__51679),
            .I(N__51676));
    Odrv4 I__11867 (
            .O(N__51676),
            .I(n3182));
    InMux I__11866 (
            .O(N__51673),
            .I(n12510));
    InMux I__11865 (
            .O(N__51670),
            .I(N__51667));
    LocalMux I__11864 (
            .O(N__51667),
            .I(N__51664));
    Span4Mux_h I__11863 (
            .O(N__51664),
            .I(N__51660));
    InMux I__11862 (
            .O(N__51663),
            .I(N__51657));
    Span4Mux_v I__11861 (
            .O(N__51660),
            .I(N__51654));
    LocalMux I__11860 (
            .O(N__51657),
            .I(n3114));
    Odrv4 I__11859 (
            .O(N__51654),
            .I(n3114));
    InMux I__11858 (
            .O(N__51649),
            .I(N__51646));
    LocalMux I__11857 (
            .O(N__51646),
            .I(n3181));
    InMux I__11856 (
            .O(N__51643),
            .I(n12511));
    InMux I__11855 (
            .O(N__51640),
            .I(N__51636));
    InMux I__11854 (
            .O(N__51639),
            .I(N__51633));
    LocalMux I__11853 (
            .O(N__51636),
            .I(N__51629));
    LocalMux I__11852 (
            .O(N__51633),
            .I(N__51626));
    InMux I__11851 (
            .O(N__51632),
            .I(N__51623));
    Span4Mux_v I__11850 (
            .O(N__51629),
            .I(N__51618));
    Span4Mux_h I__11849 (
            .O(N__51626),
            .I(N__51618));
    LocalMux I__11848 (
            .O(N__51623),
            .I(n3113));
    Odrv4 I__11847 (
            .O(N__51618),
            .I(n3113));
    CascadeMux I__11846 (
            .O(N__51613),
            .I(N__51610));
    InMux I__11845 (
            .O(N__51610),
            .I(N__51607));
    LocalMux I__11844 (
            .O(N__51607),
            .I(N__51604));
    Span4Mux_h I__11843 (
            .O(N__51604),
            .I(N__51601));
    Span4Mux_h I__11842 (
            .O(N__51601),
            .I(N__51598));
    Odrv4 I__11841 (
            .O(N__51598),
            .I(n3180));
    InMux I__11840 (
            .O(N__51595),
            .I(n12512));
    InMux I__11839 (
            .O(N__51592),
            .I(N__51589));
    LocalMux I__11838 (
            .O(N__51589),
            .I(N__51585));
    InMux I__11837 (
            .O(N__51588),
            .I(N__51582));
    Span4Mux_h I__11836 (
            .O(N__51585),
            .I(N__51579));
    LocalMux I__11835 (
            .O(N__51582),
            .I(N__51576));
    Odrv4 I__11834 (
            .O(N__51579),
            .I(n3112));
    Odrv4 I__11833 (
            .O(N__51576),
            .I(n3112));
    InMux I__11832 (
            .O(N__51571),
            .I(N__51568));
    LocalMux I__11831 (
            .O(N__51568),
            .I(N__51565));
    Span4Mux_h I__11830 (
            .O(N__51565),
            .I(N__51562));
    Odrv4 I__11829 (
            .O(N__51562),
            .I(n3179));
    InMux I__11828 (
            .O(N__51559),
            .I(n12513));
    InMux I__11827 (
            .O(N__51556),
            .I(N__51552));
    CascadeMux I__11826 (
            .O(N__51555),
            .I(N__51549));
    LocalMux I__11825 (
            .O(N__51552),
            .I(N__51545));
    InMux I__11824 (
            .O(N__51549),
            .I(N__51542));
    InMux I__11823 (
            .O(N__51548),
            .I(N__51539));
    Span4Mux_h I__11822 (
            .O(N__51545),
            .I(N__51536));
    LocalMux I__11821 (
            .O(N__51542),
            .I(N__51533));
    LocalMux I__11820 (
            .O(N__51539),
            .I(N__51530));
    Span4Mux_v I__11819 (
            .O(N__51536),
            .I(N__51523));
    Span4Mux_v I__11818 (
            .O(N__51533),
            .I(N__51523));
    Span4Mux_h I__11817 (
            .O(N__51530),
            .I(N__51523));
    Odrv4 I__11816 (
            .O(N__51523),
            .I(n3126));
    CascadeMux I__11815 (
            .O(N__51520),
            .I(N__51517));
    InMux I__11814 (
            .O(N__51517),
            .I(N__51514));
    LocalMux I__11813 (
            .O(N__51514),
            .I(N__51511));
    Span4Mux_h I__11812 (
            .O(N__51511),
            .I(N__51508));
    Span4Mux_h I__11811 (
            .O(N__51508),
            .I(N__51505));
    Odrv4 I__11810 (
            .O(N__51505),
            .I(n3193));
    InMux I__11809 (
            .O(N__51502),
            .I(bfn_16_23_0_));
    InMux I__11808 (
            .O(N__51499),
            .I(N__51494));
    InMux I__11807 (
            .O(N__51498),
            .I(N__51491));
    InMux I__11806 (
            .O(N__51497),
            .I(N__51488));
    LocalMux I__11805 (
            .O(N__51494),
            .I(N__51485));
    LocalMux I__11804 (
            .O(N__51491),
            .I(N__51482));
    LocalMux I__11803 (
            .O(N__51488),
            .I(N__51479));
    Span4Mux_h I__11802 (
            .O(N__51485),
            .I(N__51476));
    Span4Mux_h I__11801 (
            .O(N__51482),
            .I(N__51473));
    Odrv4 I__11800 (
            .O(N__51479),
            .I(n3125));
    Odrv4 I__11799 (
            .O(N__51476),
            .I(n3125));
    Odrv4 I__11798 (
            .O(N__51473),
            .I(n3125));
    CascadeMux I__11797 (
            .O(N__51466),
            .I(N__51463));
    InMux I__11796 (
            .O(N__51463),
            .I(N__51460));
    LocalMux I__11795 (
            .O(N__51460),
            .I(N__51457));
    Span4Mux_v I__11794 (
            .O(N__51457),
            .I(N__51454));
    Odrv4 I__11793 (
            .O(N__51454),
            .I(n3192));
    InMux I__11792 (
            .O(N__51451),
            .I(n12500));
    InMux I__11791 (
            .O(N__51448),
            .I(N__51445));
    LocalMux I__11790 (
            .O(N__51445),
            .I(N__51441));
    InMux I__11789 (
            .O(N__51444),
            .I(N__51438));
    Span4Mux_v I__11788 (
            .O(N__51441),
            .I(N__51435));
    LocalMux I__11787 (
            .O(N__51438),
            .I(N__51431));
    Span4Mux_h I__11786 (
            .O(N__51435),
            .I(N__51428));
    InMux I__11785 (
            .O(N__51434),
            .I(N__51425));
    Odrv4 I__11784 (
            .O(N__51431),
            .I(n3124));
    Odrv4 I__11783 (
            .O(N__51428),
            .I(n3124));
    LocalMux I__11782 (
            .O(N__51425),
            .I(n3124));
    InMux I__11781 (
            .O(N__51418),
            .I(N__51415));
    LocalMux I__11780 (
            .O(N__51415),
            .I(N__51412));
    Odrv12 I__11779 (
            .O(N__51412),
            .I(n3191));
    InMux I__11778 (
            .O(N__51409),
            .I(n12501));
    CascadeMux I__11777 (
            .O(N__51406),
            .I(N__51402));
    InMux I__11776 (
            .O(N__51405),
            .I(N__51399));
    InMux I__11775 (
            .O(N__51402),
            .I(N__51396));
    LocalMux I__11774 (
            .O(N__51399),
            .I(N__51392));
    LocalMux I__11773 (
            .O(N__51396),
            .I(N__51389));
    InMux I__11772 (
            .O(N__51395),
            .I(N__51386));
    Span4Mux_v I__11771 (
            .O(N__51392),
            .I(N__51383));
    Span4Mux_h I__11770 (
            .O(N__51389),
            .I(N__51380));
    LocalMux I__11769 (
            .O(N__51386),
            .I(N__51377));
    Span4Mux_h I__11768 (
            .O(N__51383),
            .I(N__51372));
    Span4Mux_v I__11767 (
            .O(N__51380),
            .I(N__51372));
    Odrv4 I__11766 (
            .O(N__51377),
            .I(n3123));
    Odrv4 I__11765 (
            .O(N__51372),
            .I(n3123));
    CascadeMux I__11764 (
            .O(N__51367),
            .I(N__51364));
    InMux I__11763 (
            .O(N__51364),
            .I(N__51361));
    LocalMux I__11762 (
            .O(N__51361),
            .I(N__51358));
    Span4Mux_v I__11761 (
            .O(N__51358),
            .I(N__51355));
    Odrv4 I__11760 (
            .O(N__51355),
            .I(n3190));
    InMux I__11759 (
            .O(N__51352),
            .I(n12502));
    InMux I__11758 (
            .O(N__51349),
            .I(N__51345));
    CascadeMux I__11757 (
            .O(N__51348),
            .I(N__51342));
    LocalMux I__11756 (
            .O(N__51345),
            .I(N__51339));
    InMux I__11755 (
            .O(N__51342),
            .I(N__51336));
    Span4Mux_h I__11754 (
            .O(N__51339),
            .I(N__51333));
    LocalMux I__11753 (
            .O(N__51336),
            .I(N__51330));
    Odrv4 I__11752 (
            .O(N__51333),
            .I(n3122));
    Odrv12 I__11751 (
            .O(N__51330),
            .I(n3122));
    InMux I__11750 (
            .O(N__51325),
            .I(N__51322));
    LocalMux I__11749 (
            .O(N__51322),
            .I(N__51319));
    Span4Mux_v I__11748 (
            .O(N__51319),
            .I(N__51316));
    Odrv4 I__11747 (
            .O(N__51316),
            .I(n3189));
    InMux I__11746 (
            .O(N__51313),
            .I(n12503));
    InMux I__11745 (
            .O(N__51310),
            .I(N__51306));
    InMux I__11744 (
            .O(N__51309),
            .I(N__51303));
    LocalMux I__11743 (
            .O(N__51306),
            .I(N__51300));
    LocalMux I__11742 (
            .O(N__51303),
            .I(N__51297));
    Span4Mux_h I__11741 (
            .O(N__51300),
            .I(N__51294));
    Odrv12 I__11740 (
            .O(N__51297),
            .I(n3121));
    Odrv4 I__11739 (
            .O(N__51294),
            .I(n3121));
    InMux I__11738 (
            .O(N__51289),
            .I(N__51286));
    LocalMux I__11737 (
            .O(N__51286),
            .I(N__51283));
    Span4Mux_h I__11736 (
            .O(N__51283),
            .I(N__51280));
    Odrv4 I__11735 (
            .O(N__51280),
            .I(n3188));
    InMux I__11734 (
            .O(N__51277),
            .I(n12504));
    InMux I__11733 (
            .O(N__51274),
            .I(N__51269));
    InMux I__11732 (
            .O(N__51273),
            .I(N__51266));
    InMux I__11731 (
            .O(N__51272),
            .I(N__51263));
    LocalMux I__11730 (
            .O(N__51269),
            .I(N__51260));
    LocalMux I__11729 (
            .O(N__51266),
            .I(N__51257));
    LocalMux I__11728 (
            .O(N__51263),
            .I(N__51254));
    Span4Mux_h I__11727 (
            .O(N__51260),
            .I(N__51251));
    Span4Mux_h I__11726 (
            .O(N__51257),
            .I(N__51248));
    Odrv4 I__11725 (
            .O(N__51254),
            .I(n3120));
    Odrv4 I__11724 (
            .O(N__51251),
            .I(n3120));
    Odrv4 I__11723 (
            .O(N__51248),
            .I(n3120));
    CascadeMux I__11722 (
            .O(N__51241),
            .I(N__51238));
    InMux I__11721 (
            .O(N__51238),
            .I(N__51235));
    LocalMux I__11720 (
            .O(N__51235),
            .I(N__51232));
    Span4Mux_h I__11719 (
            .O(N__51232),
            .I(N__51229));
    Odrv4 I__11718 (
            .O(N__51229),
            .I(n3187));
    InMux I__11717 (
            .O(N__51226),
            .I(n12505));
    InMux I__11716 (
            .O(N__51223),
            .I(N__51219));
    InMux I__11715 (
            .O(N__51222),
            .I(N__51216));
    LocalMux I__11714 (
            .O(N__51219),
            .I(N__51213));
    LocalMux I__11713 (
            .O(N__51216),
            .I(N__51207));
    Span12Mux_v I__11712 (
            .O(N__51213),
            .I(N__51207));
    InMux I__11711 (
            .O(N__51212),
            .I(N__51204));
    Odrv12 I__11710 (
            .O(N__51207),
            .I(n3119));
    LocalMux I__11709 (
            .O(N__51204),
            .I(n3119));
    CascadeMux I__11708 (
            .O(N__51199),
            .I(N__51196));
    InMux I__11707 (
            .O(N__51196),
            .I(N__51193));
    LocalMux I__11706 (
            .O(N__51193),
            .I(N__51190));
    Span4Mux_h I__11705 (
            .O(N__51190),
            .I(N__51187));
    Odrv4 I__11704 (
            .O(N__51187),
            .I(n3186));
    InMux I__11703 (
            .O(N__51184),
            .I(n12506));
    InMux I__11702 (
            .O(N__51181),
            .I(N__51177));
    InMux I__11701 (
            .O(N__51180),
            .I(N__51173));
    LocalMux I__11700 (
            .O(N__51177),
            .I(N__51170));
    InMux I__11699 (
            .O(N__51176),
            .I(N__51167));
    LocalMux I__11698 (
            .O(N__51173),
            .I(N__51164));
    Span4Mux_v I__11697 (
            .O(N__51170),
            .I(N__51159));
    LocalMux I__11696 (
            .O(N__51167),
            .I(N__51159));
    Sp12to4 I__11695 (
            .O(N__51164),
            .I(N__51156));
    Span4Mux_h I__11694 (
            .O(N__51159),
            .I(N__51153));
    Span12Mux_v I__11693 (
            .O(N__51156),
            .I(N__51150));
    Span4Mux_v I__11692 (
            .O(N__51153),
            .I(N__51147));
    Span12Mux_h I__11691 (
            .O(N__51150),
            .I(N__51144));
    Odrv4 I__11690 (
            .O(N__51147),
            .I(n317));
    Odrv12 I__11689 (
            .O(N__51144),
            .I(n317));
    InMux I__11688 (
            .O(N__51139),
            .I(N__51136));
    LocalMux I__11687 (
            .O(N__51136),
            .I(N__51133));
    Span4Mux_h I__11686 (
            .O(N__51133),
            .I(N__51130));
    Span4Mux_h I__11685 (
            .O(N__51130),
            .I(N__51127));
    Span4Mux_h I__11684 (
            .O(N__51127),
            .I(N__51124));
    Odrv4 I__11683 (
            .O(N__51124),
            .I(n3201));
    InMux I__11682 (
            .O(N__51121),
            .I(bfn_16_22_0_));
    CascadeMux I__11681 (
            .O(N__51118),
            .I(N__51114));
    CascadeMux I__11680 (
            .O(N__51117),
            .I(N__51111));
    InMux I__11679 (
            .O(N__51114),
            .I(N__51107));
    InMux I__11678 (
            .O(N__51111),
            .I(N__51102));
    InMux I__11677 (
            .O(N__51110),
            .I(N__51102));
    LocalMux I__11676 (
            .O(N__51107),
            .I(N__51099));
    LocalMux I__11675 (
            .O(N__51102),
            .I(n3133));
    Odrv12 I__11674 (
            .O(N__51099),
            .I(n3133));
    InMux I__11673 (
            .O(N__51094),
            .I(N__51091));
    LocalMux I__11672 (
            .O(N__51091),
            .I(N__51088));
    Span4Mux_h I__11671 (
            .O(N__51088),
            .I(N__51085));
    Span4Mux_h I__11670 (
            .O(N__51085),
            .I(N__51082));
    Odrv4 I__11669 (
            .O(N__51082),
            .I(n3200));
    InMux I__11668 (
            .O(N__51079),
            .I(n12492));
    CascadeMux I__11667 (
            .O(N__51076),
            .I(N__51073));
    InMux I__11666 (
            .O(N__51073),
            .I(N__51070));
    LocalMux I__11665 (
            .O(N__51070),
            .I(N__51065));
    InMux I__11664 (
            .O(N__51069),
            .I(N__51062));
    CascadeMux I__11663 (
            .O(N__51068),
            .I(N__51059));
    Span4Mux_h I__11662 (
            .O(N__51065),
            .I(N__51056));
    LocalMux I__11661 (
            .O(N__51062),
            .I(N__51053));
    InMux I__11660 (
            .O(N__51059),
            .I(N__51050));
    Span4Mux_h I__11659 (
            .O(N__51056),
            .I(N__51047));
    Odrv4 I__11658 (
            .O(N__51053),
            .I(n3132));
    LocalMux I__11657 (
            .O(N__51050),
            .I(n3132));
    Odrv4 I__11656 (
            .O(N__51047),
            .I(n3132));
    CascadeMux I__11655 (
            .O(N__51040),
            .I(N__51037));
    InMux I__11654 (
            .O(N__51037),
            .I(N__51034));
    LocalMux I__11653 (
            .O(N__51034),
            .I(N__51031));
    Span4Mux_v I__11652 (
            .O(N__51031),
            .I(N__51028));
    Span4Mux_h I__11651 (
            .O(N__51028),
            .I(N__51025));
    Odrv4 I__11650 (
            .O(N__51025),
            .I(n3199));
    InMux I__11649 (
            .O(N__51022),
            .I(n12493));
    CascadeMux I__11648 (
            .O(N__51019),
            .I(N__51016));
    InMux I__11647 (
            .O(N__51016),
            .I(N__51013));
    LocalMux I__11646 (
            .O(N__51013),
            .I(N__51008));
    InMux I__11645 (
            .O(N__51012),
            .I(N__51003));
    InMux I__11644 (
            .O(N__51011),
            .I(N__51003));
    Odrv12 I__11643 (
            .O(N__51008),
            .I(n3131));
    LocalMux I__11642 (
            .O(N__51003),
            .I(n3131));
    InMux I__11641 (
            .O(N__50998),
            .I(N__50995));
    LocalMux I__11640 (
            .O(N__50995),
            .I(N__50992));
    Span12Mux_s10_v I__11639 (
            .O(N__50992),
            .I(N__50989));
    Odrv12 I__11638 (
            .O(N__50989),
            .I(n3198));
    InMux I__11637 (
            .O(N__50986),
            .I(n12494));
    CascadeMux I__11636 (
            .O(N__50983),
            .I(N__50979));
    InMux I__11635 (
            .O(N__50982),
            .I(N__50975));
    InMux I__11634 (
            .O(N__50979),
            .I(N__50972));
    InMux I__11633 (
            .O(N__50978),
            .I(N__50969));
    LocalMux I__11632 (
            .O(N__50975),
            .I(N__50966));
    LocalMux I__11631 (
            .O(N__50972),
            .I(N__50963));
    LocalMux I__11630 (
            .O(N__50969),
            .I(N__50960));
    Span4Mux_v I__11629 (
            .O(N__50966),
            .I(N__50953));
    Span4Mux_h I__11628 (
            .O(N__50963),
            .I(N__50953));
    Span4Mux_v I__11627 (
            .O(N__50960),
            .I(N__50953));
    Odrv4 I__11626 (
            .O(N__50953),
            .I(n3130));
    CascadeMux I__11625 (
            .O(N__50950),
            .I(N__50947));
    InMux I__11624 (
            .O(N__50947),
            .I(N__50944));
    LocalMux I__11623 (
            .O(N__50944),
            .I(N__50941));
    Span4Mux_h I__11622 (
            .O(N__50941),
            .I(N__50938));
    Span4Mux_h I__11621 (
            .O(N__50938),
            .I(N__50935));
    Odrv4 I__11620 (
            .O(N__50935),
            .I(n3197));
    InMux I__11619 (
            .O(N__50932),
            .I(n12495));
    InMux I__11618 (
            .O(N__50929),
            .I(N__50925));
    InMux I__11617 (
            .O(N__50928),
            .I(N__50921));
    LocalMux I__11616 (
            .O(N__50925),
            .I(N__50918));
    InMux I__11615 (
            .O(N__50924),
            .I(N__50915));
    LocalMux I__11614 (
            .O(N__50921),
            .I(N__50912));
    Span4Mux_h I__11613 (
            .O(N__50918),
            .I(N__50909));
    LocalMux I__11612 (
            .O(N__50915),
            .I(N__50906));
    Span4Mux_h I__11611 (
            .O(N__50912),
            .I(N__50903));
    Odrv4 I__11610 (
            .O(N__50909),
            .I(n3129));
    Odrv12 I__11609 (
            .O(N__50906),
            .I(n3129));
    Odrv4 I__11608 (
            .O(N__50903),
            .I(n3129));
    CascadeMux I__11607 (
            .O(N__50896),
            .I(N__50893));
    InMux I__11606 (
            .O(N__50893),
            .I(N__50890));
    LocalMux I__11605 (
            .O(N__50890),
            .I(N__50887));
    Span4Mux_h I__11604 (
            .O(N__50887),
            .I(N__50884));
    Odrv4 I__11603 (
            .O(N__50884),
            .I(n3196));
    InMux I__11602 (
            .O(N__50881),
            .I(n12496));
    CascadeMux I__11601 (
            .O(N__50878),
            .I(N__50874));
    InMux I__11600 (
            .O(N__50877),
            .I(N__50871));
    InMux I__11599 (
            .O(N__50874),
            .I(N__50868));
    LocalMux I__11598 (
            .O(N__50871),
            .I(N__50865));
    LocalMux I__11597 (
            .O(N__50868),
            .I(N__50862));
    Span4Mux_v I__11596 (
            .O(N__50865),
            .I(N__50859));
    Span4Mux_h I__11595 (
            .O(N__50862),
            .I(N__50856));
    Span4Mux_v I__11594 (
            .O(N__50859),
            .I(N__50852));
    Span4Mux_h I__11593 (
            .O(N__50856),
            .I(N__50849));
    InMux I__11592 (
            .O(N__50855),
            .I(N__50846));
    Odrv4 I__11591 (
            .O(N__50852),
            .I(n3128));
    Odrv4 I__11590 (
            .O(N__50849),
            .I(n3128));
    LocalMux I__11589 (
            .O(N__50846),
            .I(n3128));
    InMux I__11588 (
            .O(N__50839),
            .I(N__50836));
    LocalMux I__11587 (
            .O(N__50836),
            .I(N__50833));
    Span4Mux_v I__11586 (
            .O(N__50833),
            .I(N__50830));
    Odrv4 I__11585 (
            .O(N__50830),
            .I(n3195));
    InMux I__11584 (
            .O(N__50827),
            .I(n12497));
    CascadeMux I__11583 (
            .O(N__50824),
            .I(N__50821));
    InMux I__11582 (
            .O(N__50821),
            .I(N__50817));
    CascadeMux I__11581 (
            .O(N__50820),
            .I(N__50814));
    LocalMux I__11580 (
            .O(N__50817),
            .I(N__50811));
    InMux I__11579 (
            .O(N__50814),
            .I(N__50808));
    Span4Mux_v I__11578 (
            .O(N__50811),
            .I(N__50803));
    LocalMux I__11577 (
            .O(N__50808),
            .I(N__50803));
    Span4Mux_v I__11576 (
            .O(N__50803),
            .I(N__50800));
    Span4Mux_h I__11575 (
            .O(N__50800),
            .I(N__50796));
    InMux I__11574 (
            .O(N__50799),
            .I(N__50793));
    Odrv4 I__11573 (
            .O(N__50796),
            .I(n3127));
    LocalMux I__11572 (
            .O(N__50793),
            .I(n3127));
    InMux I__11571 (
            .O(N__50788),
            .I(N__50785));
    LocalMux I__11570 (
            .O(N__50785),
            .I(N__50782));
    Odrv4 I__11569 (
            .O(N__50782),
            .I(n3194));
    InMux I__11568 (
            .O(N__50779),
            .I(n12498));
    InMux I__11567 (
            .O(N__50776),
            .I(N__50772));
    InMux I__11566 (
            .O(N__50775),
            .I(N__50769));
    LocalMux I__11565 (
            .O(N__50772),
            .I(sweep_counter_10));
    LocalMux I__11564 (
            .O(N__50769),
            .I(sweep_counter_10));
    InMux I__11563 (
            .O(N__50764),
            .I(n12615));
    InMux I__11562 (
            .O(N__50761),
            .I(N__50757));
    InMux I__11561 (
            .O(N__50760),
            .I(N__50754));
    LocalMux I__11560 (
            .O(N__50757),
            .I(sweep_counter_11));
    LocalMux I__11559 (
            .O(N__50754),
            .I(sweep_counter_11));
    InMux I__11558 (
            .O(N__50749),
            .I(n12616));
    InMux I__11557 (
            .O(N__50746),
            .I(N__50742));
    InMux I__11556 (
            .O(N__50745),
            .I(N__50739));
    LocalMux I__11555 (
            .O(N__50742),
            .I(sweep_counter_12));
    LocalMux I__11554 (
            .O(N__50739),
            .I(sweep_counter_12));
    InMux I__11553 (
            .O(N__50734),
            .I(n12617));
    InMux I__11552 (
            .O(N__50731),
            .I(N__50727));
    InMux I__11551 (
            .O(N__50730),
            .I(N__50724));
    LocalMux I__11550 (
            .O(N__50727),
            .I(sweep_counter_13));
    LocalMux I__11549 (
            .O(N__50724),
            .I(sweep_counter_13));
    InMux I__11548 (
            .O(N__50719),
            .I(n12618));
    CascadeMux I__11547 (
            .O(N__50716),
            .I(N__50712));
    InMux I__11546 (
            .O(N__50715),
            .I(N__50709));
    InMux I__11545 (
            .O(N__50712),
            .I(N__50706));
    LocalMux I__11544 (
            .O(N__50709),
            .I(sweep_counter_14));
    LocalMux I__11543 (
            .O(N__50706),
            .I(sweep_counter_14));
    InMux I__11542 (
            .O(N__50701),
            .I(n12619));
    CascadeMux I__11541 (
            .O(N__50698),
            .I(N__50694));
    InMux I__11540 (
            .O(N__50697),
            .I(N__50691));
    InMux I__11539 (
            .O(N__50694),
            .I(N__50688));
    LocalMux I__11538 (
            .O(N__50691),
            .I(sweep_counter_15));
    LocalMux I__11537 (
            .O(N__50688),
            .I(sweep_counter_15));
    InMux I__11536 (
            .O(N__50683),
            .I(n12620));
    InMux I__11535 (
            .O(N__50680),
            .I(N__50676));
    InMux I__11534 (
            .O(N__50679),
            .I(N__50673));
    LocalMux I__11533 (
            .O(N__50676),
            .I(sweep_counter_16));
    LocalMux I__11532 (
            .O(N__50673),
            .I(sweep_counter_16));
    InMux I__11531 (
            .O(N__50668),
            .I(bfn_16_19_0_));
    InMux I__11530 (
            .O(N__50665),
            .I(n12622));
    InMux I__11529 (
            .O(N__50662),
            .I(N__50658));
    InMux I__11528 (
            .O(N__50661),
            .I(N__50655));
    LocalMux I__11527 (
            .O(N__50658),
            .I(sweep_counter_17));
    LocalMux I__11526 (
            .O(N__50655),
            .I(sweep_counter_17));
    InMux I__11525 (
            .O(N__50650),
            .I(N__50646));
    InMux I__11524 (
            .O(N__50649),
            .I(N__50643));
    LocalMux I__11523 (
            .O(N__50646),
            .I(sweep_counter_1));
    LocalMux I__11522 (
            .O(N__50643),
            .I(sweep_counter_1));
    InMux I__11521 (
            .O(N__50638),
            .I(n12606));
    CascadeMux I__11520 (
            .O(N__50635),
            .I(N__50631));
    InMux I__11519 (
            .O(N__50634),
            .I(N__50628));
    InMux I__11518 (
            .O(N__50631),
            .I(N__50625));
    LocalMux I__11517 (
            .O(N__50628),
            .I(sweep_counter_2));
    LocalMux I__11516 (
            .O(N__50625),
            .I(sweep_counter_2));
    InMux I__11515 (
            .O(N__50620),
            .I(n12607));
    InMux I__11514 (
            .O(N__50617),
            .I(N__50613));
    InMux I__11513 (
            .O(N__50616),
            .I(N__50610));
    LocalMux I__11512 (
            .O(N__50613),
            .I(sweep_counter_3));
    LocalMux I__11511 (
            .O(N__50610),
            .I(sweep_counter_3));
    InMux I__11510 (
            .O(N__50605),
            .I(n12608));
    InMux I__11509 (
            .O(N__50602),
            .I(N__50598));
    InMux I__11508 (
            .O(N__50601),
            .I(N__50595));
    LocalMux I__11507 (
            .O(N__50598),
            .I(sweep_counter_4));
    LocalMux I__11506 (
            .O(N__50595),
            .I(sweep_counter_4));
    InMux I__11505 (
            .O(N__50590),
            .I(n12609));
    InMux I__11504 (
            .O(N__50587),
            .I(N__50583));
    InMux I__11503 (
            .O(N__50586),
            .I(N__50580));
    LocalMux I__11502 (
            .O(N__50583),
            .I(sweep_counter_5));
    LocalMux I__11501 (
            .O(N__50580),
            .I(sweep_counter_5));
    InMux I__11500 (
            .O(N__50575),
            .I(n12610));
    CascadeMux I__11499 (
            .O(N__50572),
            .I(N__50568));
    InMux I__11498 (
            .O(N__50571),
            .I(N__50565));
    InMux I__11497 (
            .O(N__50568),
            .I(N__50562));
    LocalMux I__11496 (
            .O(N__50565),
            .I(N__50557));
    LocalMux I__11495 (
            .O(N__50562),
            .I(N__50557));
    Odrv4 I__11494 (
            .O(N__50557),
            .I(sweep_counter_6));
    InMux I__11493 (
            .O(N__50554),
            .I(n12611));
    InMux I__11492 (
            .O(N__50551),
            .I(N__50547));
    InMux I__11491 (
            .O(N__50550),
            .I(N__50544));
    LocalMux I__11490 (
            .O(N__50547),
            .I(sweep_counter_7));
    LocalMux I__11489 (
            .O(N__50544),
            .I(sweep_counter_7));
    InMux I__11488 (
            .O(N__50539),
            .I(n12612));
    InMux I__11487 (
            .O(N__50536),
            .I(N__50532));
    InMux I__11486 (
            .O(N__50535),
            .I(N__50529));
    LocalMux I__11485 (
            .O(N__50532),
            .I(sweep_counter_8));
    LocalMux I__11484 (
            .O(N__50529),
            .I(sweep_counter_8));
    InMux I__11483 (
            .O(N__50524),
            .I(bfn_16_18_0_));
    InMux I__11482 (
            .O(N__50521),
            .I(N__50517));
    InMux I__11481 (
            .O(N__50520),
            .I(N__50514));
    LocalMux I__11480 (
            .O(N__50517),
            .I(sweep_counter_9));
    LocalMux I__11479 (
            .O(N__50514),
            .I(sweep_counter_9));
    InMux I__11478 (
            .O(N__50509),
            .I(n12614));
    CascadeMux I__11477 (
            .O(N__50506),
            .I(\quad_counter0.direction_N_534_cascade_ ));
    InMux I__11476 (
            .O(N__50503),
            .I(N__50500));
    LocalMux I__11475 (
            .O(N__50500),
            .I(\quad_counter0.a_prev_N_537 ));
    CascadeMux I__11474 (
            .O(N__50497),
            .I(N__50494));
    InMux I__11473 (
            .O(N__50494),
            .I(N__50488));
    InMux I__11472 (
            .O(N__50493),
            .I(N__50488));
    LocalMux I__11471 (
            .O(N__50488),
            .I(\quad_counter0.a_prev ));
    InMux I__11470 (
            .O(N__50485),
            .I(N__50473));
    InMux I__11469 (
            .O(N__50484),
            .I(N__50473));
    InMux I__11468 (
            .O(N__50483),
            .I(N__50473));
    InMux I__11467 (
            .O(N__50482),
            .I(N__50473));
    LocalMux I__11466 (
            .O(N__50473),
            .I(\quad_counter0.b_new_1 ));
    CascadeMux I__11465 (
            .O(N__50470),
            .I(N__50466));
    InMux I__11464 (
            .O(N__50469),
            .I(N__50462));
    InMux I__11463 (
            .O(N__50466),
            .I(N__50457));
    InMux I__11462 (
            .O(N__50465),
            .I(N__50457));
    LocalMux I__11461 (
            .O(N__50462),
            .I(N__50452));
    LocalMux I__11460 (
            .O(N__50457),
            .I(N__50452));
    Odrv12 I__11459 (
            .O(N__50452),
            .I(\quad_counter0.b_new_0 ));
    InMux I__11458 (
            .O(N__50449),
            .I(N__50440));
    InMux I__11457 (
            .O(N__50448),
            .I(N__50440));
    InMux I__11456 (
            .O(N__50447),
            .I(N__50440));
    LocalMux I__11455 (
            .O(N__50440),
            .I(\quad_counter0.debounce_cnt ));
    CEMux I__11454 (
            .O(N__50437),
            .I(N__50433));
    CEMux I__11453 (
            .O(N__50436),
            .I(N__50428));
    LocalMux I__11452 (
            .O(N__50433),
            .I(N__50425));
    CEMux I__11451 (
            .O(N__50432),
            .I(N__50422));
    CEMux I__11450 (
            .O(N__50431),
            .I(N__50419));
    LocalMux I__11449 (
            .O(N__50428),
            .I(N__50416));
    Span4Mux_v I__11448 (
            .O(N__50425),
            .I(N__50411));
    LocalMux I__11447 (
            .O(N__50422),
            .I(N__50411));
    LocalMux I__11446 (
            .O(N__50419),
            .I(N__50408));
    Span4Mux_v I__11445 (
            .O(N__50416),
            .I(N__50403));
    Span4Mux_h I__11444 (
            .O(N__50411),
            .I(N__50403));
    Span4Mux_h I__11443 (
            .O(N__50408),
            .I(N__50400));
    Span4Mux_h I__11442 (
            .O(N__50403),
            .I(N__50397));
    Span4Mux_h I__11441 (
            .O(N__50400),
            .I(N__50394));
    Span4Mux_h I__11440 (
            .O(N__50397),
            .I(N__50390));
    Span4Mux_h I__11439 (
            .O(N__50394),
            .I(N__50387));
    InMux I__11438 (
            .O(N__50393),
            .I(N__50384));
    Odrv4 I__11437 (
            .O(N__50390),
            .I(direction_N_531));
    Odrv4 I__11436 (
            .O(N__50387),
            .I(direction_N_531));
    LocalMux I__11435 (
            .O(N__50384),
            .I(direction_N_531));
    CascadeMux I__11434 (
            .O(N__50377),
            .I(N__50373));
    InMux I__11433 (
            .O(N__50376),
            .I(N__50368));
    InMux I__11432 (
            .O(N__50373),
            .I(N__50365));
    InMux I__11431 (
            .O(N__50372),
            .I(N__50362));
    InMux I__11430 (
            .O(N__50371),
            .I(N__50359));
    LocalMux I__11429 (
            .O(N__50368),
            .I(N__50356));
    LocalMux I__11428 (
            .O(N__50365),
            .I(b_prev));
    LocalMux I__11427 (
            .O(N__50362),
            .I(b_prev));
    LocalMux I__11426 (
            .O(N__50359),
            .I(b_prev));
    Odrv4 I__11425 (
            .O(N__50356),
            .I(b_prev));
    InMux I__11424 (
            .O(N__50347),
            .I(N__50344));
    LocalMux I__11423 (
            .O(N__50344),
            .I(n1185));
    InMux I__11422 (
            .O(N__50341),
            .I(N__50338));
    LocalMux I__11421 (
            .O(N__50338),
            .I(N__50335));
    Span4Mux_s3_v I__11420 (
            .O(N__50335),
            .I(N__50330));
    InMux I__11419 (
            .O(N__50334),
            .I(N__50325));
    InMux I__11418 (
            .O(N__50333),
            .I(N__50325));
    Sp12to4 I__11417 (
            .O(N__50330),
            .I(N__50320));
    LocalMux I__11416 (
            .O(N__50325),
            .I(N__50320));
    Odrv12 I__11415 (
            .O(N__50320),
            .I(\quad_counter0.a_new_0 ));
    CascadeMux I__11414 (
            .O(N__50317),
            .I(N__50311));
    InMux I__11413 (
            .O(N__50316),
            .I(N__50306));
    InMux I__11412 (
            .O(N__50315),
            .I(N__50303));
    InMux I__11411 (
            .O(N__50314),
            .I(N__50298));
    InMux I__11410 (
            .O(N__50311),
            .I(N__50298));
    InMux I__11409 (
            .O(N__50310),
            .I(N__50293));
    InMux I__11408 (
            .O(N__50309),
            .I(N__50293));
    LocalMux I__11407 (
            .O(N__50306),
            .I(N__50290));
    LocalMux I__11406 (
            .O(N__50303),
            .I(a_new_1));
    LocalMux I__11405 (
            .O(N__50298),
            .I(a_new_1));
    LocalMux I__11404 (
            .O(N__50293),
            .I(a_new_1));
    Odrv4 I__11403 (
            .O(N__50290),
            .I(a_new_1));
    InMux I__11402 (
            .O(N__50281),
            .I(N__50278));
    LocalMux I__11401 (
            .O(N__50278),
            .I(N__50274));
    InMux I__11400 (
            .O(N__50277),
            .I(N__50271));
    Span4Mux_v I__11399 (
            .O(N__50274),
            .I(N__50268));
    LocalMux I__11398 (
            .O(N__50271),
            .I(N__50265));
    Odrv4 I__11397 (
            .O(N__50268),
            .I(duty_19));
    Odrv4 I__11396 (
            .O(N__50265),
            .I(duty_19));
    InMux I__11395 (
            .O(N__50260),
            .I(N__50257));
    LocalMux I__11394 (
            .O(N__50257),
            .I(N__50254));
    Odrv4 I__11393 (
            .O(N__50254),
            .I(n6_adj_572));
    InMux I__11392 (
            .O(N__50251),
            .I(N__50247));
    InMux I__11391 (
            .O(N__50250),
            .I(N__50244));
    LocalMux I__11390 (
            .O(N__50247),
            .I(N__50241));
    LocalMux I__11389 (
            .O(N__50244),
            .I(N__50238));
    Odrv4 I__11388 (
            .O(N__50241),
            .I(duty_18));
    Odrv4 I__11387 (
            .O(N__50238),
            .I(duty_18));
    InMux I__11386 (
            .O(N__50233),
            .I(N__50230));
    LocalMux I__11385 (
            .O(N__50230),
            .I(N__50227));
    Span4Mux_h I__11384 (
            .O(N__50227),
            .I(N__50224));
    Odrv4 I__11383 (
            .O(N__50224),
            .I(n7_adj_573));
    InMux I__11382 (
            .O(N__50221),
            .I(N__50217));
    InMux I__11381 (
            .O(N__50220),
            .I(N__50214));
    LocalMux I__11380 (
            .O(N__50217),
            .I(sweep_counter_0));
    LocalMux I__11379 (
            .O(N__50214),
            .I(sweep_counter_0));
    InMux I__11378 (
            .O(N__50209),
            .I(bfn_16_17_0_));
    InMux I__11377 (
            .O(N__50206),
            .I(N__50203));
    LocalMux I__11376 (
            .O(N__50203),
            .I(N__50200));
    Odrv4 I__11375 (
            .O(N__50200),
            .I(n24_adj_590));
    InMux I__11374 (
            .O(N__50197),
            .I(N__50194));
    LocalMux I__11373 (
            .O(N__50194),
            .I(N__50191));
    Span4Mux_v I__11372 (
            .O(N__50191),
            .I(N__50187));
    InMux I__11371 (
            .O(N__50190),
            .I(N__50184));
    Span4Mux_h I__11370 (
            .O(N__50187),
            .I(N__50181));
    LocalMux I__11369 (
            .O(N__50184),
            .I(N__50178));
    Odrv4 I__11368 (
            .O(N__50181),
            .I(duty_3));
    Odrv4 I__11367 (
            .O(N__50178),
            .I(duty_3));
    InMux I__11366 (
            .O(N__50173),
            .I(N__50170));
    LocalMux I__11365 (
            .O(N__50170),
            .I(N__50167));
    Odrv4 I__11364 (
            .O(N__50167),
            .I(n22_adj_588));
    CascadeMux I__11363 (
            .O(N__50164),
            .I(n21_adj_700_cascade_));
    InMux I__11362 (
            .O(N__50161),
            .I(N__50158));
    LocalMux I__11361 (
            .O(N__50158),
            .I(n22_adj_699));
    InMux I__11360 (
            .O(N__50155),
            .I(N__50151));
    InMux I__11359 (
            .O(N__50154),
            .I(N__50148));
    LocalMux I__11358 (
            .O(N__50151),
            .I(N__50143));
    LocalMux I__11357 (
            .O(N__50148),
            .I(N__50143));
    Span4Mux_h I__11356 (
            .O(N__50143),
            .I(N__50140));
    Odrv4 I__11355 (
            .O(N__50140),
            .I(duty_1));
    InMux I__11354 (
            .O(N__50137),
            .I(N__50134));
    LocalMux I__11353 (
            .O(N__50134),
            .I(N__50131));
    Odrv4 I__11352 (
            .O(N__50131),
            .I(pwm_setpoint_23_N_171_1));
    InMux I__11351 (
            .O(N__50128),
            .I(N__50125));
    LocalMux I__11350 (
            .O(N__50125),
            .I(pwm_setpoint_1));
    CascadeMux I__11349 (
            .O(N__50122),
            .I(\quad_counter0.a_prev_N_537_cascade_ ));
    CascadeMux I__11348 (
            .O(N__50119),
            .I(N__50114));
    CascadeMux I__11347 (
            .O(N__50118),
            .I(N__50110));
    InMux I__11346 (
            .O(N__50117),
            .I(N__50098));
    InMux I__11345 (
            .O(N__50114),
            .I(N__50098));
    InMux I__11344 (
            .O(N__50113),
            .I(N__50098));
    InMux I__11343 (
            .O(N__50110),
            .I(N__50090));
    InMux I__11342 (
            .O(N__50109),
            .I(N__50090));
    InMux I__11341 (
            .O(N__50108),
            .I(N__50087));
    InMux I__11340 (
            .O(N__50107),
            .I(N__50082));
    InMux I__11339 (
            .O(N__50106),
            .I(N__50079));
    CascadeMux I__11338 (
            .O(N__50105),
            .I(N__50074));
    LocalMux I__11337 (
            .O(N__50098),
            .I(N__50065));
    InMux I__11336 (
            .O(N__50097),
            .I(N__50058));
    InMux I__11335 (
            .O(N__50096),
            .I(N__50058));
    InMux I__11334 (
            .O(N__50095),
            .I(N__50058));
    LocalMux I__11333 (
            .O(N__50090),
            .I(N__50053));
    LocalMux I__11332 (
            .O(N__50087),
            .I(N__50053));
    InMux I__11331 (
            .O(N__50086),
            .I(N__50048));
    InMux I__11330 (
            .O(N__50085),
            .I(N__50048));
    LocalMux I__11329 (
            .O(N__50082),
            .I(N__50045));
    LocalMux I__11328 (
            .O(N__50079),
            .I(N__50042));
    InMux I__11327 (
            .O(N__50078),
            .I(N__50033));
    InMux I__11326 (
            .O(N__50077),
            .I(N__50033));
    InMux I__11325 (
            .O(N__50074),
            .I(N__50033));
    InMux I__11324 (
            .O(N__50073),
            .I(N__50033));
    CascadeMux I__11323 (
            .O(N__50072),
            .I(N__50029));
    CascadeMux I__11322 (
            .O(N__50071),
            .I(N__50026));
    CascadeMux I__11321 (
            .O(N__50070),
            .I(N__50020));
    CascadeMux I__11320 (
            .O(N__50069),
            .I(N__50016));
    InMux I__11319 (
            .O(N__50068),
            .I(N__50010));
    Sp12to4 I__11318 (
            .O(N__50065),
            .I(N__50005));
    LocalMux I__11317 (
            .O(N__50058),
            .I(N__50005));
    Span4Mux_h I__11316 (
            .O(N__50053),
            .I(N__50002));
    LocalMux I__11315 (
            .O(N__50048),
            .I(N__49999));
    Span4Mux_v I__11314 (
            .O(N__50045),
            .I(N__49992));
    Span4Mux_v I__11313 (
            .O(N__50042),
            .I(N__49992));
    LocalMux I__11312 (
            .O(N__50033),
            .I(N__49992));
    InMux I__11311 (
            .O(N__50032),
            .I(N__49989));
    InMux I__11310 (
            .O(N__50029),
            .I(N__49980));
    InMux I__11309 (
            .O(N__50026),
            .I(N__49980));
    InMux I__11308 (
            .O(N__50025),
            .I(N__49980));
    InMux I__11307 (
            .O(N__50024),
            .I(N__49980));
    InMux I__11306 (
            .O(N__50023),
            .I(N__49977));
    InMux I__11305 (
            .O(N__50020),
            .I(N__49972));
    InMux I__11304 (
            .O(N__50019),
            .I(N__49972));
    InMux I__11303 (
            .O(N__50016),
            .I(N__49963));
    InMux I__11302 (
            .O(N__50015),
            .I(N__49963));
    InMux I__11301 (
            .O(N__50014),
            .I(N__49963));
    InMux I__11300 (
            .O(N__50013),
            .I(N__49963));
    LocalMux I__11299 (
            .O(N__50010),
            .I(N__49958));
    Span12Mux_s8_v I__11298 (
            .O(N__50005),
            .I(N__49958));
    Span4Mux_h I__11297 (
            .O(N__50002),
            .I(N__49955));
    Span4Mux_h I__11296 (
            .O(N__49999),
            .I(N__49950));
    Span4Mux_h I__11295 (
            .O(N__49992),
            .I(N__49950));
    LocalMux I__11294 (
            .O(N__49989),
            .I(n3138));
    LocalMux I__11293 (
            .O(N__49980),
            .I(n3138));
    LocalMux I__11292 (
            .O(N__49977),
            .I(n3138));
    LocalMux I__11291 (
            .O(N__49972),
            .I(n3138));
    LocalMux I__11290 (
            .O(N__49963),
            .I(n3138));
    Odrv12 I__11289 (
            .O(N__49958),
            .I(n3138));
    Odrv4 I__11288 (
            .O(N__49955),
            .I(n3138));
    Odrv4 I__11287 (
            .O(N__49950),
            .I(n3138));
    CascadeMux I__11286 (
            .O(N__49933),
            .I(n3114_cascade_));
    InMux I__11285 (
            .O(N__49930),
            .I(N__49925));
    InMux I__11284 (
            .O(N__49929),
            .I(N__49922));
    InMux I__11283 (
            .O(N__49928),
            .I(N__49919));
    LocalMux I__11282 (
            .O(N__49925),
            .I(N__49916));
    LocalMux I__11281 (
            .O(N__49922),
            .I(N__49913));
    LocalMux I__11280 (
            .O(N__49919),
            .I(N__49910));
    Span4Mux_h I__11279 (
            .O(N__49916),
            .I(N__49907));
    Odrv4 I__11278 (
            .O(N__49913),
            .I(n3213));
    Odrv4 I__11277 (
            .O(N__49910),
            .I(n3213));
    Odrv4 I__11276 (
            .O(N__49907),
            .I(n3213));
    CascadeMux I__11275 (
            .O(N__49900),
            .I(n7_adj_712_cascade_));
    InMux I__11274 (
            .O(N__49897),
            .I(N__49894));
    LocalMux I__11273 (
            .O(N__49894),
            .I(n8_adj_711));
    CascadeMux I__11272 (
            .O(N__49891),
            .I(N__49876));
    CascadeMux I__11271 (
            .O(N__49890),
            .I(N__49872));
    CascadeMux I__11270 (
            .O(N__49889),
            .I(N__49868));
    CascadeMux I__11269 (
            .O(N__49888),
            .I(N__49864));
    CascadeMux I__11268 (
            .O(N__49887),
            .I(N__49861));
    CascadeMux I__11267 (
            .O(N__49886),
            .I(N__49857));
    CascadeMux I__11266 (
            .O(N__49885),
            .I(N__49853));
    CascadeMux I__11265 (
            .O(N__49884),
            .I(N__49849));
    CascadeMux I__11264 (
            .O(N__49883),
            .I(N__49845));
    CascadeMux I__11263 (
            .O(N__49882),
            .I(N__49841));
    CascadeMux I__11262 (
            .O(N__49881),
            .I(N__49837));
    CascadeMux I__11261 (
            .O(N__49880),
            .I(N__49833));
    InMux I__11260 (
            .O(N__49879),
            .I(N__49812));
    InMux I__11259 (
            .O(N__49876),
            .I(N__49812));
    InMux I__11258 (
            .O(N__49875),
            .I(N__49812));
    InMux I__11257 (
            .O(N__49872),
            .I(N__49812));
    InMux I__11256 (
            .O(N__49871),
            .I(N__49812));
    InMux I__11255 (
            .O(N__49868),
            .I(N__49812));
    InMux I__11254 (
            .O(N__49867),
            .I(N__49812));
    InMux I__11253 (
            .O(N__49864),
            .I(N__49812));
    InMux I__11252 (
            .O(N__49861),
            .I(N__49795));
    InMux I__11251 (
            .O(N__49860),
            .I(N__49795));
    InMux I__11250 (
            .O(N__49857),
            .I(N__49795));
    InMux I__11249 (
            .O(N__49856),
            .I(N__49795));
    InMux I__11248 (
            .O(N__49853),
            .I(N__49795));
    InMux I__11247 (
            .O(N__49852),
            .I(N__49795));
    InMux I__11246 (
            .O(N__49849),
            .I(N__49795));
    InMux I__11245 (
            .O(N__49848),
            .I(N__49795));
    InMux I__11244 (
            .O(N__49845),
            .I(N__49778));
    InMux I__11243 (
            .O(N__49844),
            .I(N__49778));
    InMux I__11242 (
            .O(N__49841),
            .I(N__49778));
    InMux I__11241 (
            .O(N__49840),
            .I(N__49778));
    InMux I__11240 (
            .O(N__49837),
            .I(N__49778));
    InMux I__11239 (
            .O(N__49836),
            .I(N__49778));
    InMux I__11238 (
            .O(N__49833),
            .I(N__49778));
    InMux I__11237 (
            .O(N__49832),
            .I(N__49778));
    CascadeMux I__11236 (
            .O(N__49831),
            .I(N__49774));
    CascadeMux I__11235 (
            .O(N__49830),
            .I(N__49770));
    CascadeMux I__11234 (
            .O(N__49829),
            .I(N__49766));
    LocalMux I__11233 (
            .O(N__49812),
            .I(N__49758));
    LocalMux I__11232 (
            .O(N__49795),
            .I(N__49758));
    LocalMux I__11231 (
            .O(N__49778),
            .I(N__49758));
    InMux I__11230 (
            .O(N__49777),
            .I(N__49743));
    InMux I__11229 (
            .O(N__49774),
            .I(N__49743));
    InMux I__11228 (
            .O(N__49773),
            .I(N__49743));
    InMux I__11227 (
            .O(N__49770),
            .I(N__49743));
    InMux I__11226 (
            .O(N__49769),
            .I(N__49743));
    InMux I__11225 (
            .O(N__49766),
            .I(N__49743));
    InMux I__11224 (
            .O(N__49765),
            .I(N__49743));
    Span4Mux_v I__11223 (
            .O(N__49758),
            .I(N__49740));
    LocalMux I__11222 (
            .O(N__49743),
            .I(N__49737));
    Span4Mux_h I__11221 (
            .O(N__49740),
            .I(N__49732));
    Span4Mux_h I__11220 (
            .O(N__49737),
            .I(N__49732));
    Span4Mux_v I__11219 (
            .O(N__49732),
            .I(N__49729));
    Span4Mux_h I__11218 (
            .O(N__49729),
            .I(N__49726));
    Odrv4 I__11217 (
            .O(N__49726),
            .I(\quad_counter0.direction_N_530 ));
    InMux I__11216 (
            .O(N__49723),
            .I(N__49720));
    LocalMux I__11215 (
            .O(N__49720),
            .I(n13676));
    CascadeMux I__11214 (
            .O(N__49717),
            .I(n10_adj_714_cascade_));
    CascadeMux I__11213 (
            .O(N__49714),
            .I(n16_adj_702_cascade_));
    InMux I__11212 (
            .O(N__49711),
            .I(N__49708));
    LocalMux I__11211 (
            .O(N__49708),
            .I(n19_adj_701));
    InMux I__11210 (
            .O(N__49705),
            .I(N__49702));
    LocalMux I__11209 (
            .O(N__49702),
            .I(N__49699));
    Span4Mux_v I__11208 (
            .O(N__49699),
            .I(N__49696));
    Odrv4 I__11207 (
            .O(N__49696),
            .I(n3286));
    CascadeMux I__11206 (
            .O(N__49693),
            .I(n27_adj_709_cascade_));
    InMux I__11205 (
            .O(N__49690),
            .I(N__49685));
    InMux I__11204 (
            .O(N__49689),
            .I(N__49682));
    InMux I__11203 (
            .O(N__49688),
            .I(N__49679));
    LocalMux I__11202 (
            .O(N__49685),
            .I(n3219));
    LocalMux I__11201 (
            .O(N__49682),
            .I(n3219));
    LocalMux I__11200 (
            .O(N__49679),
            .I(n3219));
    InMux I__11199 (
            .O(N__49672),
            .I(N__49669));
    LocalMux I__11198 (
            .O(N__49669),
            .I(n13830));
    InMux I__11197 (
            .O(N__49666),
            .I(N__49663));
    LocalMux I__11196 (
            .O(N__49663),
            .I(N__49660));
    Odrv4 I__11195 (
            .O(N__49660),
            .I(n3292));
    CascadeMux I__11194 (
            .O(N__49657),
            .I(N__49652));
    InMux I__11193 (
            .O(N__49656),
            .I(N__49649));
    InMux I__11192 (
            .O(N__49655),
            .I(N__49646));
    InMux I__11191 (
            .O(N__49652),
            .I(N__49643));
    LocalMux I__11190 (
            .O(N__49649),
            .I(N__49640));
    LocalMux I__11189 (
            .O(N__49646),
            .I(N__49637));
    LocalMux I__11188 (
            .O(N__49643),
            .I(N__49634));
    Span4Mux_v I__11187 (
            .O(N__49640),
            .I(N__49629));
    Span4Mux_h I__11186 (
            .O(N__49637),
            .I(N__49629));
    Span4Mux_h I__11185 (
            .O(N__49634),
            .I(N__49626));
    Span4Mux_h I__11184 (
            .O(N__49629),
            .I(N__49623));
    Odrv4 I__11183 (
            .O(N__49626),
            .I(n3225));
    Odrv4 I__11182 (
            .O(N__49623),
            .I(n3225));
    InMux I__11181 (
            .O(N__49618),
            .I(N__49609));
    InMux I__11180 (
            .O(N__49617),
            .I(N__49593));
    InMux I__11179 (
            .O(N__49616),
            .I(N__49593));
    InMux I__11178 (
            .O(N__49615),
            .I(N__49593));
    InMux I__11177 (
            .O(N__49614),
            .I(N__49593));
    InMux I__11176 (
            .O(N__49613),
            .I(N__49593));
    CascadeMux I__11175 (
            .O(N__49612),
            .I(N__49590));
    LocalMux I__11174 (
            .O(N__49609),
            .I(N__49586));
    CascadeMux I__11173 (
            .O(N__49608),
            .I(N__49578));
    CascadeMux I__11172 (
            .O(N__49607),
            .I(N__49574));
    CascadeMux I__11171 (
            .O(N__49606),
            .I(N__49570));
    CascadeMux I__11170 (
            .O(N__49605),
            .I(N__49558));
    CascadeMux I__11169 (
            .O(N__49604),
            .I(N__49555));
    LocalMux I__11168 (
            .O(N__49593),
            .I(N__49551));
    InMux I__11167 (
            .O(N__49590),
            .I(N__49546));
    InMux I__11166 (
            .O(N__49589),
            .I(N__49546));
    Span4Mux_v I__11165 (
            .O(N__49586),
            .I(N__49543));
    InMux I__11164 (
            .O(N__49585),
            .I(N__49530));
    InMux I__11163 (
            .O(N__49584),
            .I(N__49530));
    InMux I__11162 (
            .O(N__49583),
            .I(N__49530));
    InMux I__11161 (
            .O(N__49582),
            .I(N__49530));
    InMux I__11160 (
            .O(N__49581),
            .I(N__49530));
    InMux I__11159 (
            .O(N__49578),
            .I(N__49530));
    InMux I__11158 (
            .O(N__49577),
            .I(N__49519));
    InMux I__11157 (
            .O(N__49574),
            .I(N__49519));
    InMux I__11156 (
            .O(N__49573),
            .I(N__49519));
    InMux I__11155 (
            .O(N__49570),
            .I(N__49519));
    InMux I__11154 (
            .O(N__49569),
            .I(N__49519));
    InMux I__11153 (
            .O(N__49568),
            .I(N__49506));
    InMux I__11152 (
            .O(N__49567),
            .I(N__49506));
    InMux I__11151 (
            .O(N__49566),
            .I(N__49506));
    InMux I__11150 (
            .O(N__49565),
            .I(N__49506));
    InMux I__11149 (
            .O(N__49564),
            .I(N__49506));
    InMux I__11148 (
            .O(N__49563),
            .I(N__49506));
    InMux I__11147 (
            .O(N__49562),
            .I(N__49495));
    InMux I__11146 (
            .O(N__49561),
            .I(N__49495));
    InMux I__11145 (
            .O(N__49558),
            .I(N__49495));
    InMux I__11144 (
            .O(N__49555),
            .I(N__49495));
    InMux I__11143 (
            .O(N__49554),
            .I(N__49495));
    Span4Mux_h I__11142 (
            .O(N__49551),
            .I(N__49490));
    LocalMux I__11141 (
            .O(N__49546),
            .I(N__49490));
    Odrv4 I__11140 (
            .O(N__49543),
            .I(n3237));
    LocalMux I__11139 (
            .O(N__49530),
            .I(n3237));
    LocalMux I__11138 (
            .O(N__49519),
            .I(n3237));
    LocalMux I__11137 (
            .O(N__49506),
            .I(n3237));
    LocalMux I__11136 (
            .O(N__49495),
            .I(n3237));
    Odrv4 I__11135 (
            .O(N__49490),
            .I(n3237));
    InMux I__11134 (
            .O(N__49477),
            .I(N__49474));
    LocalMux I__11133 (
            .O(N__49474),
            .I(n21_adj_706));
    InMux I__11132 (
            .O(N__49471),
            .I(N__49467));
    InMux I__11131 (
            .O(N__49470),
            .I(N__49464));
    LocalMux I__11130 (
            .O(N__49467),
            .I(N__49458));
    LocalMux I__11129 (
            .O(N__49464),
            .I(N__49458));
    InMux I__11128 (
            .O(N__49463),
            .I(N__49455));
    Span4Mux_v I__11127 (
            .O(N__49458),
            .I(N__49450));
    LocalMux I__11126 (
            .O(N__49455),
            .I(N__49450));
    Odrv4 I__11125 (
            .O(N__49450),
            .I(n3011));
    CascadeMux I__11124 (
            .O(N__49447),
            .I(N__49444));
    InMux I__11123 (
            .O(N__49444),
            .I(N__49441));
    LocalMux I__11122 (
            .O(N__49441),
            .I(N__49438));
    Span4Mux_h I__11121 (
            .O(N__49438),
            .I(N__49435));
    Odrv4 I__11120 (
            .O(N__49435),
            .I(n3078));
    CascadeMux I__11119 (
            .O(N__49432),
            .I(n3110_cascade_));
    InMux I__11118 (
            .O(N__49429),
            .I(N__49424));
    InMux I__11117 (
            .O(N__49428),
            .I(N__49421));
    InMux I__11116 (
            .O(N__49427),
            .I(N__49418));
    LocalMux I__11115 (
            .O(N__49424),
            .I(N__49413));
    LocalMux I__11114 (
            .O(N__49421),
            .I(N__49413));
    LocalMux I__11113 (
            .O(N__49418),
            .I(N__49408));
    Span4Mux_v I__11112 (
            .O(N__49413),
            .I(N__49408));
    Span4Mux_h I__11111 (
            .O(N__49408),
            .I(N__49405));
    Odrv4 I__11110 (
            .O(N__49405),
            .I(n3209));
    CascadeMux I__11109 (
            .O(N__49402),
            .I(N__49399));
    InMux I__11108 (
            .O(N__49399),
            .I(N__49395));
    InMux I__11107 (
            .O(N__49398),
            .I(N__49392));
    LocalMux I__11106 (
            .O(N__49395),
            .I(N__49387));
    LocalMux I__11105 (
            .O(N__49392),
            .I(N__49387));
    Span4Mux_h I__11104 (
            .O(N__49387),
            .I(N__49383));
    InMux I__11103 (
            .O(N__49386),
            .I(N__49380));
    Odrv4 I__11102 (
            .O(N__49383),
            .I(n3226));
    LocalMux I__11101 (
            .O(N__49380),
            .I(n3226));
    CascadeMux I__11100 (
            .O(N__49375),
            .I(N__49368));
    InMux I__11099 (
            .O(N__49374),
            .I(N__49363));
    InMux I__11098 (
            .O(N__49373),
            .I(N__49360));
    InMux I__11097 (
            .O(N__49372),
            .I(N__49355));
    InMux I__11096 (
            .O(N__49371),
            .I(N__49350));
    InMux I__11095 (
            .O(N__49368),
            .I(N__49347));
    InMux I__11094 (
            .O(N__49367),
            .I(N__49344));
    InMux I__11093 (
            .O(N__49366),
            .I(N__49341));
    LocalMux I__11092 (
            .O(N__49363),
            .I(N__49337));
    LocalMux I__11091 (
            .O(N__49360),
            .I(N__49333));
    InMux I__11090 (
            .O(N__49359),
            .I(N__49330));
    CascadeMux I__11089 (
            .O(N__49358),
            .I(N__49327));
    LocalMux I__11088 (
            .O(N__49355),
            .I(N__49321));
    CascadeMux I__11087 (
            .O(N__49354),
            .I(N__49317));
    CascadeMux I__11086 (
            .O(N__49353),
            .I(N__49313));
    LocalMux I__11085 (
            .O(N__49350),
            .I(N__49303));
    LocalMux I__11084 (
            .O(N__49347),
            .I(N__49303));
    LocalMux I__11083 (
            .O(N__49344),
            .I(N__49303));
    LocalMux I__11082 (
            .O(N__49341),
            .I(N__49303));
    CascadeMux I__11081 (
            .O(N__49340),
            .I(N__49299));
    Span4Mux_v I__11080 (
            .O(N__49337),
            .I(N__49289));
    InMux I__11079 (
            .O(N__49336),
            .I(N__49286));
    Span4Mux_h I__11078 (
            .O(N__49333),
            .I(N__49281));
    LocalMux I__11077 (
            .O(N__49330),
            .I(N__49281));
    InMux I__11076 (
            .O(N__49327),
            .I(N__49274));
    InMux I__11075 (
            .O(N__49326),
            .I(N__49274));
    InMux I__11074 (
            .O(N__49325),
            .I(N__49274));
    InMux I__11073 (
            .O(N__49324),
            .I(N__49270));
    Span4Mux_v I__11072 (
            .O(N__49321),
            .I(N__49267));
    InMux I__11071 (
            .O(N__49320),
            .I(N__49264));
    InMux I__11070 (
            .O(N__49317),
            .I(N__49255));
    InMux I__11069 (
            .O(N__49316),
            .I(N__49255));
    InMux I__11068 (
            .O(N__49313),
            .I(N__49255));
    InMux I__11067 (
            .O(N__49312),
            .I(N__49255));
    Span4Mux_v I__11066 (
            .O(N__49303),
            .I(N__49252));
    InMux I__11065 (
            .O(N__49302),
            .I(N__49245));
    InMux I__11064 (
            .O(N__49299),
            .I(N__49245));
    InMux I__11063 (
            .O(N__49298),
            .I(N__49245));
    InMux I__11062 (
            .O(N__49297),
            .I(N__49232));
    InMux I__11061 (
            .O(N__49296),
            .I(N__49232));
    InMux I__11060 (
            .O(N__49295),
            .I(N__49232));
    InMux I__11059 (
            .O(N__49294),
            .I(N__49232));
    InMux I__11058 (
            .O(N__49293),
            .I(N__49232));
    InMux I__11057 (
            .O(N__49292),
            .I(N__49232));
    Span4Mux_h I__11056 (
            .O(N__49289),
            .I(N__49223));
    LocalMux I__11055 (
            .O(N__49286),
            .I(N__49223));
    Span4Mux_v I__11054 (
            .O(N__49281),
            .I(N__49223));
    LocalMux I__11053 (
            .O(N__49274),
            .I(N__49223));
    InMux I__11052 (
            .O(N__49273),
            .I(N__49220));
    LocalMux I__11051 (
            .O(N__49270),
            .I(n2841));
    Odrv4 I__11050 (
            .O(N__49267),
            .I(n2841));
    LocalMux I__11049 (
            .O(N__49264),
            .I(n2841));
    LocalMux I__11048 (
            .O(N__49255),
            .I(n2841));
    Odrv4 I__11047 (
            .O(N__49252),
            .I(n2841));
    LocalMux I__11046 (
            .O(N__49245),
            .I(n2841));
    LocalMux I__11045 (
            .O(N__49232),
            .I(n2841));
    Odrv4 I__11044 (
            .O(N__49223),
            .I(n2841));
    LocalMux I__11043 (
            .O(N__49220),
            .I(n2841));
    InMux I__11042 (
            .O(N__49201),
            .I(N__49198));
    LocalMux I__11041 (
            .O(N__49198),
            .I(N__49195));
    Span4Mux_h I__11040 (
            .O(N__49195),
            .I(N__49192));
    Odrv4 I__11039 (
            .O(N__49192),
            .I(n14921));
    InMux I__11038 (
            .O(N__49189),
            .I(N__49186));
    LocalMux I__11037 (
            .O(N__49186),
            .I(N__49182));
    InMux I__11036 (
            .O(N__49185),
            .I(N__49179));
    Span4Mux_h I__11035 (
            .O(N__49182),
            .I(N__49174));
    LocalMux I__11034 (
            .O(N__49179),
            .I(N__49174));
    Span4Mux_v I__11033 (
            .O(N__49174),
            .I(N__49170));
    InMux I__11032 (
            .O(N__49173),
            .I(N__49167));
    Odrv4 I__11031 (
            .O(N__49170),
            .I(n3009));
    LocalMux I__11030 (
            .O(N__49167),
            .I(n3009));
    CascadeMux I__11029 (
            .O(N__49162),
            .I(N__49159));
    InMux I__11028 (
            .O(N__49159),
            .I(N__49156));
    LocalMux I__11027 (
            .O(N__49156),
            .I(n3076));
    InMux I__11026 (
            .O(N__49153),
            .I(N__49150));
    LocalMux I__11025 (
            .O(N__49150),
            .I(N__49147));
    Span4Mux_v I__11024 (
            .O(N__49147),
            .I(N__49144));
    Span4Mux_h I__11023 (
            .O(N__49144),
            .I(N__49141));
    Span4Mux_h I__11022 (
            .O(N__49141),
            .I(N__49138));
    Span4Mux_v I__11021 (
            .O(N__49138),
            .I(N__49135));
    Sp12to4 I__11020 (
            .O(N__49135),
            .I(N__49132));
    Odrv12 I__11019 (
            .O(N__49132),
            .I(ENCODER0_B_N));
    InMux I__11018 (
            .O(N__49129),
            .I(N__49126));
    LocalMux I__11017 (
            .O(N__49126),
            .I(N__49122));
    InMux I__11016 (
            .O(N__49125),
            .I(N__49119));
    Span4Mux_v I__11015 (
            .O(N__49122),
            .I(N__49115));
    LocalMux I__11014 (
            .O(N__49119),
            .I(N__49112));
    InMux I__11013 (
            .O(N__49118),
            .I(N__49109));
    Span4Mux_h I__11012 (
            .O(N__49115),
            .I(N__49106));
    Span4Mux_v I__11011 (
            .O(N__49112),
            .I(N__49101));
    LocalMux I__11010 (
            .O(N__49109),
            .I(N__49101));
    Odrv4 I__11009 (
            .O(N__49106),
            .I(n3015));
    Odrv4 I__11008 (
            .O(N__49101),
            .I(n3015));
    CascadeMux I__11007 (
            .O(N__49096),
            .I(N__49093));
    InMux I__11006 (
            .O(N__49093),
            .I(N__49090));
    LocalMux I__11005 (
            .O(N__49090),
            .I(N__49087));
    Odrv4 I__11004 (
            .O(N__49087),
            .I(n3082));
    CascadeMux I__11003 (
            .O(N__49084),
            .I(N__49070));
    CascadeMux I__11002 (
            .O(N__49083),
            .I(N__49066));
    CascadeMux I__11001 (
            .O(N__49082),
            .I(N__49060));
    CascadeMux I__11000 (
            .O(N__49081),
            .I(N__49057));
    InMux I__10999 (
            .O(N__49080),
            .I(N__49054));
    CascadeMux I__10998 (
            .O(N__49079),
            .I(N__49051));
    InMux I__10997 (
            .O(N__49078),
            .I(N__49044));
    InMux I__10996 (
            .O(N__49077),
            .I(N__49044));
    InMux I__10995 (
            .O(N__49076),
            .I(N__49044));
    InMux I__10994 (
            .O(N__49075),
            .I(N__49036));
    InMux I__10993 (
            .O(N__49074),
            .I(N__49031));
    InMux I__10992 (
            .O(N__49073),
            .I(N__49031));
    InMux I__10991 (
            .O(N__49070),
            .I(N__49026));
    InMux I__10990 (
            .O(N__49069),
            .I(N__49026));
    InMux I__10989 (
            .O(N__49066),
            .I(N__49021));
    InMux I__10988 (
            .O(N__49065),
            .I(N__49021));
    InMux I__10987 (
            .O(N__49064),
            .I(N__49010));
    InMux I__10986 (
            .O(N__49063),
            .I(N__49010));
    InMux I__10985 (
            .O(N__49060),
            .I(N__49010));
    InMux I__10984 (
            .O(N__49057),
            .I(N__49010));
    LocalMux I__10983 (
            .O(N__49054),
            .I(N__49007));
    InMux I__10982 (
            .O(N__49051),
            .I(N__49004));
    LocalMux I__10981 (
            .O(N__49044),
            .I(N__49001));
    CascadeMux I__10980 (
            .O(N__49043),
            .I(N__48996));
    CascadeMux I__10979 (
            .O(N__49042),
            .I(N__48992));
    CascadeMux I__10978 (
            .O(N__49041),
            .I(N__48989));
    CascadeMux I__10977 (
            .O(N__49040),
            .I(N__48985));
    CascadeMux I__10976 (
            .O(N__49039),
            .I(N__48982));
    LocalMux I__10975 (
            .O(N__49036),
            .I(N__48973));
    LocalMux I__10974 (
            .O(N__49031),
            .I(N__48973));
    LocalMux I__10973 (
            .O(N__49026),
            .I(N__48973));
    LocalMux I__10972 (
            .O(N__49021),
            .I(N__48970));
    InMux I__10971 (
            .O(N__49020),
            .I(N__48967));
    InMux I__10970 (
            .O(N__49019),
            .I(N__48964));
    LocalMux I__10969 (
            .O(N__49010),
            .I(N__48961));
    Span4Mux_h I__10968 (
            .O(N__49007),
            .I(N__48954));
    LocalMux I__10967 (
            .O(N__49004),
            .I(N__48954));
    Span4Mux_h I__10966 (
            .O(N__49001),
            .I(N__48954));
    InMux I__10965 (
            .O(N__49000),
            .I(N__48945));
    InMux I__10964 (
            .O(N__48999),
            .I(N__48945));
    InMux I__10963 (
            .O(N__48996),
            .I(N__48945));
    InMux I__10962 (
            .O(N__48995),
            .I(N__48945));
    InMux I__10961 (
            .O(N__48992),
            .I(N__48938));
    InMux I__10960 (
            .O(N__48989),
            .I(N__48938));
    InMux I__10959 (
            .O(N__48988),
            .I(N__48938));
    InMux I__10958 (
            .O(N__48985),
            .I(N__48929));
    InMux I__10957 (
            .O(N__48982),
            .I(N__48929));
    InMux I__10956 (
            .O(N__48981),
            .I(N__48929));
    InMux I__10955 (
            .O(N__48980),
            .I(N__48929));
    Span4Mux_h I__10954 (
            .O(N__48973),
            .I(N__48924));
    Span4Mux_h I__10953 (
            .O(N__48970),
            .I(N__48924));
    LocalMux I__10952 (
            .O(N__48967),
            .I(n3039));
    LocalMux I__10951 (
            .O(N__48964),
            .I(n3039));
    Odrv4 I__10950 (
            .O(N__48961),
            .I(n3039));
    Odrv4 I__10949 (
            .O(N__48954),
            .I(n3039));
    LocalMux I__10948 (
            .O(N__48945),
            .I(n3039));
    LocalMux I__10947 (
            .O(N__48938),
            .I(n3039));
    LocalMux I__10946 (
            .O(N__48929),
            .I(n3039));
    Odrv4 I__10945 (
            .O(N__48924),
            .I(n3039));
    InMux I__10944 (
            .O(N__48907),
            .I(N__48903));
    CascadeMux I__10943 (
            .O(N__48906),
            .I(N__48900));
    LocalMux I__10942 (
            .O(N__48903),
            .I(N__48897));
    InMux I__10941 (
            .O(N__48900),
            .I(N__48893));
    Span4Mux_v I__10940 (
            .O(N__48897),
            .I(N__48890));
    InMux I__10939 (
            .O(N__48896),
            .I(N__48887));
    LocalMux I__10938 (
            .O(N__48893),
            .I(n2810));
    Odrv4 I__10937 (
            .O(N__48890),
            .I(n2810));
    LocalMux I__10936 (
            .O(N__48887),
            .I(n2810));
    InMux I__10935 (
            .O(N__48880),
            .I(N__48877));
    LocalMux I__10934 (
            .O(N__48877),
            .I(N__48874));
    Span4Mux_h I__10933 (
            .O(N__48874),
            .I(N__48871));
    Odrv4 I__10932 (
            .O(N__48871),
            .I(n2877));
    InMux I__10931 (
            .O(N__48868),
            .I(bfn_15_23_0_));
    InMux I__10930 (
            .O(N__48865),
            .I(N__48860));
    InMux I__10929 (
            .O(N__48864),
            .I(N__48857));
    CascadeMux I__10928 (
            .O(N__48863),
            .I(N__48854));
    LocalMux I__10927 (
            .O(N__48860),
            .I(N__48851));
    LocalMux I__10926 (
            .O(N__48857),
            .I(N__48848));
    InMux I__10925 (
            .O(N__48854),
            .I(N__48845));
    Span4Mux_h I__10924 (
            .O(N__48851),
            .I(N__48842));
    Span4Mux_h I__10923 (
            .O(N__48848),
            .I(N__48839));
    LocalMux I__10922 (
            .O(N__48845),
            .I(N__48836));
    Span4Mux_h I__10921 (
            .O(N__48842),
            .I(N__48833));
    Span4Mux_h I__10920 (
            .O(N__48839),
            .I(N__48830));
    Odrv4 I__10919 (
            .O(N__48836),
            .I(n2809));
    Odrv4 I__10918 (
            .O(N__48833),
            .I(n2809));
    Odrv4 I__10917 (
            .O(N__48830),
            .I(n2809));
    InMux I__10916 (
            .O(N__48823),
            .I(N__48820));
    LocalMux I__10915 (
            .O(N__48820),
            .I(N__48817));
    Span4Mux_v I__10914 (
            .O(N__48817),
            .I(N__48814));
    Odrv4 I__10913 (
            .O(N__48814),
            .I(n2876));
    InMux I__10912 (
            .O(N__48811),
            .I(n12435));
    InMux I__10911 (
            .O(N__48808),
            .I(n12436));
    CascadeMux I__10910 (
            .O(N__48805),
            .I(N__48801));
    InMux I__10909 (
            .O(N__48804),
            .I(N__48795));
    InMux I__10908 (
            .O(N__48801),
            .I(N__48795));
    InMux I__10907 (
            .O(N__48800),
            .I(N__48792));
    LocalMux I__10906 (
            .O(N__48795),
            .I(N__48789));
    LocalMux I__10905 (
            .O(N__48792),
            .I(N__48786));
    Span4Mux_v I__10904 (
            .O(N__48789),
            .I(N__48783));
    Span4Mux_h I__10903 (
            .O(N__48786),
            .I(N__48780));
    Odrv4 I__10902 (
            .O(N__48783),
            .I(n2808));
    Odrv4 I__10901 (
            .O(N__48780),
            .I(n2808));
    CascadeMux I__10900 (
            .O(N__48775),
            .I(N__48772));
    InMux I__10899 (
            .O(N__48772),
            .I(N__48769));
    LocalMux I__10898 (
            .O(N__48769),
            .I(n2875));
    CascadeMux I__10897 (
            .O(N__48766),
            .I(N__48763));
    InMux I__10896 (
            .O(N__48763),
            .I(N__48760));
    LocalMux I__10895 (
            .O(N__48760),
            .I(N__48756));
    InMux I__10894 (
            .O(N__48759),
            .I(N__48753));
    Span4Mux_v I__10893 (
            .O(N__48756),
            .I(N__48748));
    LocalMux I__10892 (
            .O(N__48753),
            .I(N__48748));
    Span4Mux_h I__10891 (
            .O(N__48748),
            .I(N__48745));
    Odrv4 I__10890 (
            .O(N__48745),
            .I(n2907));
    InMux I__10889 (
            .O(N__48742),
            .I(N__48738));
    InMux I__10888 (
            .O(N__48741),
            .I(N__48735));
    LocalMux I__10887 (
            .O(N__48738),
            .I(N__48729));
    LocalMux I__10886 (
            .O(N__48735),
            .I(N__48729));
    InMux I__10885 (
            .O(N__48734),
            .I(N__48726));
    Span4Mux_v I__10884 (
            .O(N__48729),
            .I(N__48723));
    LocalMux I__10883 (
            .O(N__48726),
            .I(n3220));
    Odrv4 I__10882 (
            .O(N__48723),
            .I(n3220));
    CascadeMux I__10881 (
            .O(N__48718),
            .I(N__48715));
    InMux I__10880 (
            .O(N__48715),
            .I(N__48712));
    LocalMux I__10879 (
            .O(N__48712),
            .I(N__48709));
    Odrv12 I__10878 (
            .O(N__48709),
            .I(n3287));
    InMux I__10877 (
            .O(N__48706),
            .I(N__48703));
    LocalMux I__10876 (
            .O(N__48703),
            .I(n17_adj_705));
    InMux I__10875 (
            .O(N__48700),
            .I(N__48697));
    LocalMux I__10874 (
            .O(N__48697),
            .I(N__48694));
    Span4Mux_h I__10873 (
            .O(N__48694),
            .I(N__48691));
    Span4Mux_h I__10872 (
            .O(N__48691),
            .I(N__48688));
    Odrv4 I__10871 (
            .O(N__48688),
            .I(n3296));
    CascadeMux I__10870 (
            .O(N__48685),
            .I(n13822_cascade_));
    InMux I__10869 (
            .O(N__48682),
            .I(N__48678));
    InMux I__10868 (
            .O(N__48681),
            .I(N__48675));
    LocalMux I__10867 (
            .O(N__48678),
            .I(N__48672));
    LocalMux I__10866 (
            .O(N__48675),
            .I(N__48669));
    Span4Mux_h I__10865 (
            .O(N__48672),
            .I(N__48666));
    Odrv12 I__10864 (
            .O(N__48669),
            .I(n3229));
    Odrv4 I__10863 (
            .O(N__48666),
            .I(n3229));
    InMux I__10862 (
            .O(N__48661),
            .I(N__48658));
    LocalMux I__10861 (
            .O(N__48658),
            .I(n15_adj_704));
    CascadeMux I__10860 (
            .O(N__48655),
            .I(n13834_cascade_));
    InMux I__10859 (
            .O(N__48652),
            .I(N__48649));
    LocalMux I__10858 (
            .O(N__48649),
            .I(N__48646));
    Odrv4 I__10857 (
            .O(N__48646),
            .I(n13842));
    InMux I__10856 (
            .O(N__48643),
            .I(N__48640));
    LocalMux I__10855 (
            .O(N__48640),
            .I(N__48636));
    InMux I__10854 (
            .O(N__48639),
            .I(N__48632));
    Span4Mux_h I__10853 (
            .O(N__48636),
            .I(N__48629));
    InMux I__10852 (
            .O(N__48635),
            .I(N__48626));
    LocalMux I__10851 (
            .O(N__48632),
            .I(N__48623));
    Odrv4 I__10850 (
            .O(N__48629),
            .I(n3222));
    LocalMux I__10849 (
            .O(N__48626),
            .I(n3222));
    Odrv12 I__10848 (
            .O(N__48623),
            .I(n3222));
    CascadeMux I__10847 (
            .O(N__48616),
            .I(N__48613));
    InMux I__10846 (
            .O(N__48613),
            .I(N__48610));
    LocalMux I__10845 (
            .O(N__48610),
            .I(N__48607));
    Odrv4 I__10844 (
            .O(N__48607),
            .I(n3289));
    InMux I__10843 (
            .O(N__48604),
            .I(N__48601));
    LocalMux I__10842 (
            .O(N__48601),
            .I(N__48598));
    Span4Mux_h I__10841 (
            .O(N__48598),
            .I(N__48595));
    Odrv4 I__10840 (
            .O(N__48595),
            .I(n2885));
    InMux I__10839 (
            .O(N__48592),
            .I(bfn_15_22_0_));
    InMux I__10838 (
            .O(N__48589),
            .I(N__48586));
    LocalMux I__10837 (
            .O(N__48586),
            .I(N__48582));
    InMux I__10836 (
            .O(N__48585),
            .I(N__48579));
    Span4Mux_v I__10835 (
            .O(N__48582),
            .I(N__48574));
    LocalMux I__10834 (
            .O(N__48579),
            .I(N__48574));
    Span4Mux_h I__10833 (
            .O(N__48574),
            .I(N__48571));
    Odrv4 I__10832 (
            .O(N__48571),
            .I(n2817));
    InMux I__10831 (
            .O(N__48568),
            .I(N__48565));
    LocalMux I__10830 (
            .O(N__48565),
            .I(N__48562));
    Span4Mux_h I__10829 (
            .O(N__48562),
            .I(N__48559));
    Odrv4 I__10828 (
            .O(N__48559),
            .I(n2884));
    InMux I__10827 (
            .O(N__48556),
            .I(n12427));
    InMux I__10826 (
            .O(N__48553),
            .I(N__48549));
    InMux I__10825 (
            .O(N__48552),
            .I(N__48546));
    LocalMux I__10824 (
            .O(N__48549),
            .I(N__48542));
    LocalMux I__10823 (
            .O(N__48546),
            .I(N__48539));
    InMux I__10822 (
            .O(N__48545),
            .I(N__48536));
    Span4Mux_h I__10821 (
            .O(N__48542),
            .I(N__48533));
    Span4Mux_v I__10820 (
            .O(N__48539),
            .I(N__48528));
    LocalMux I__10819 (
            .O(N__48536),
            .I(N__48528));
    Odrv4 I__10818 (
            .O(N__48533),
            .I(n2816));
    Odrv4 I__10817 (
            .O(N__48528),
            .I(n2816));
    CascadeMux I__10816 (
            .O(N__48523),
            .I(N__48520));
    InMux I__10815 (
            .O(N__48520),
            .I(N__48517));
    LocalMux I__10814 (
            .O(N__48517),
            .I(N__48514));
    Span4Mux_h I__10813 (
            .O(N__48514),
            .I(N__48511));
    Odrv4 I__10812 (
            .O(N__48511),
            .I(n2883));
    InMux I__10811 (
            .O(N__48508),
            .I(n12428));
    InMux I__10810 (
            .O(N__48505),
            .I(N__48501));
    InMux I__10809 (
            .O(N__48504),
            .I(N__48498));
    LocalMux I__10808 (
            .O(N__48501),
            .I(N__48495));
    LocalMux I__10807 (
            .O(N__48498),
            .I(N__48489));
    Span4Mux_v I__10806 (
            .O(N__48495),
            .I(N__48489));
    InMux I__10805 (
            .O(N__48494),
            .I(N__48486));
    Odrv4 I__10804 (
            .O(N__48489),
            .I(n2815));
    LocalMux I__10803 (
            .O(N__48486),
            .I(n2815));
    InMux I__10802 (
            .O(N__48481),
            .I(N__48478));
    LocalMux I__10801 (
            .O(N__48478),
            .I(N__48475));
    Odrv4 I__10800 (
            .O(N__48475),
            .I(n2882));
    InMux I__10799 (
            .O(N__48472),
            .I(n12429));
    CascadeMux I__10798 (
            .O(N__48469),
            .I(N__48466));
    InMux I__10797 (
            .O(N__48466),
            .I(N__48462));
    InMux I__10796 (
            .O(N__48465),
            .I(N__48459));
    LocalMux I__10795 (
            .O(N__48462),
            .I(N__48456));
    LocalMux I__10794 (
            .O(N__48459),
            .I(N__48453));
    Span4Mux_v I__10793 (
            .O(N__48456),
            .I(N__48450));
    Span4Mux_v I__10792 (
            .O(N__48453),
            .I(N__48447));
    Odrv4 I__10791 (
            .O(N__48450),
            .I(n2814));
    Odrv4 I__10790 (
            .O(N__48447),
            .I(n2814));
    InMux I__10789 (
            .O(N__48442),
            .I(N__48439));
    LocalMux I__10788 (
            .O(N__48439),
            .I(N__48436));
    Odrv4 I__10787 (
            .O(N__48436),
            .I(n2881));
    InMux I__10786 (
            .O(N__48433),
            .I(n12430));
    InMux I__10785 (
            .O(N__48430),
            .I(N__48426));
    InMux I__10784 (
            .O(N__48429),
            .I(N__48422));
    LocalMux I__10783 (
            .O(N__48426),
            .I(N__48419));
    InMux I__10782 (
            .O(N__48425),
            .I(N__48416));
    LocalMux I__10781 (
            .O(N__48422),
            .I(N__48413));
    Span4Mux_v I__10780 (
            .O(N__48419),
            .I(N__48410));
    LocalMux I__10779 (
            .O(N__48416),
            .I(N__48407));
    Span4Mux_v I__10778 (
            .O(N__48413),
            .I(N__48400));
    Span4Mux_h I__10777 (
            .O(N__48410),
            .I(N__48400));
    Span4Mux_h I__10776 (
            .O(N__48407),
            .I(N__48400));
    Odrv4 I__10775 (
            .O(N__48400),
            .I(n2813));
    InMux I__10774 (
            .O(N__48397),
            .I(N__48394));
    LocalMux I__10773 (
            .O(N__48394),
            .I(N__48391));
    Odrv12 I__10772 (
            .O(N__48391),
            .I(n2880));
    InMux I__10771 (
            .O(N__48388),
            .I(n12431));
    InMux I__10770 (
            .O(N__48385),
            .I(N__48381));
    InMux I__10769 (
            .O(N__48384),
            .I(N__48378));
    LocalMux I__10768 (
            .O(N__48381),
            .I(N__48374));
    LocalMux I__10767 (
            .O(N__48378),
            .I(N__48371));
    InMux I__10766 (
            .O(N__48377),
            .I(N__48368));
    Span4Mux_h I__10765 (
            .O(N__48374),
            .I(N__48365));
    Span4Mux_h I__10764 (
            .O(N__48371),
            .I(N__48362));
    LocalMux I__10763 (
            .O(N__48368),
            .I(n2812));
    Odrv4 I__10762 (
            .O(N__48365),
            .I(n2812));
    Odrv4 I__10761 (
            .O(N__48362),
            .I(n2812));
    CascadeMux I__10760 (
            .O(N__48355),
            .I(N__48352));
    InMux I__10759 (
            .O(N__48352),
            .I(N__48349));
    LocalMux I__10758 (
            .O(N__48349),
            .I(N__48346));
    Span4Mux_h I__10757 (
            .O(N__48346),
            .I(N__48343));
    Odrv4 I__10756 (
            .O(N__48343),
            .I(n2879));
    InMux I__10755 (
            .O(N__48340),
            .I(n12432));
    InMux I__10754 (
            .O(N__48337),
            .I(N__48333));
    CascadeMux I__10753 (
            .O(N__48336),
            .I(N__48330));
    LocalMux I__10752 (
            .O(N__48333),
            .I(N__48327));
    InMux I__10751 (
            .O(N__48330),
            .I(N__48324));
    Span4Mux_v I__10750 (
            .O(N__48327),
            .I(N__48321));
    LocalMux I__10749 (
            .O(N__48324),
            .I(n2811));
    Odrv4 I__10748 (
            .O(N__48321),
            .I(n2811));
    InMux I__10747 (
            .O(N__48316),
            .I(N__48313));
    LocalMux I__10746 (
            .O(N__48313),
            .I(N__48310));
    Odrv12 I__10745 (
            .O(N__48310),
            .I(n2878));
    InMux I__10744 (
            .O(N__48307),
            .I(n12433));
    CascadeMux I__10743 (
            .O(N__48304),
            .I(N__48300));
    InMux I__10742 (
            .O(N__48303),
            .I(N__48297));
    InMux I__10741 (
            .O(N__48300),
            .I(N__48294));
    LocalMux I__10740 (
            .O(N__48297),
            .I(N__48291));
    LocalMux I__10739 (
            .O(N__48294),
            .I(n2825));
    Odrv4 I__10738 (
            .O(N__48291),
            .I(n2825));
    InMux I__10737 (
            .O(N__48286),
            .I(N__48283));
    LocalMux I__10736 (
            .O(N__48283),
            .I(n2892));
    InMux I__10735 (
            .O(N__48280),
            .I(n12419));
    CascadeMux I__10734 (
            .O(N__48277),
            .I(N__48274));
    InMux I__10733 (
            .O(N__48274),
            .I(N__48270));
    InMux I__10732 (
            .O(N__48273),
            .I(N__48267));
    LocalMux I__10731 (
            .O(N__48270),
            .I(N__48264));
    LocalMux I__10730 (
            .O(N__48267),
            .I(N__48260));
    Span4Mux_v I__10729 (
            .O(N__48264),
            .I(N__48257));
    InMux I__10728 (
            .O(N__48263),
            .I(N__48254));
    Odrv4 I__10727 (
            .O(N__48260),
            .I(n2824));
    Odrv4 I__10726 (
            .O(N__48257),
            .I(n2824));
    LocalMux I__10725 (
            .O(N__48254),
            .I(n2824));
    InMux I__10724 (
            .O(N__48247),
            .I(N__48244));
    LocalMux I__10723 (
            .O(N__48244),
            .I(N__48241));
    Odrv4 I__10722 (
            .O(N__48241),
            .I(n2891));
    InMux I__10721 (
            .O(N__48238),
            .I(n12420));
    CascadeMux I__10720 (
            .O(N__48235),
            .I(N__48231));
    CascadeMux I__10719 (
            .O(N__48234),
            .I(N__48228));
    InMux I__10718 (
            .O(N__48231),
            .I(N__48225));
    InMux I__10717 (
            .O(N__48228),
            .I(N__48221));
    LocalMux I__10716 (
            .O(N__48225),
            .I(N__48218));
    CascadeMux I__10715 (
            .O(N__48224),
            .I(N__48215));
    LocalMux I__10714 (
            .O(N__48221),
            .I(N__48210));
    Span4Mux_h I__10713 (
            .O(N__48218),
            .I(N__48210));
    InMux I__10712 (
            .O(N__48215),
            .I(N__48207));
    Odrv4 I__10711 (
            .O(N__48210),
            .I(n2823));
    LocalMux I__10710 (
            .O(N__48207),
            .I(n2823));
    InMux I__10709 (
            .O(N__48202),
            .I(N__48199));
    LocalMux I__10708 (
            .O(N__48199),
            .I(N__48196));
    Odrv4 I__10707 (
            .O(N__48196),
            .I(n2890));
    InMux I__10706 (
            .O(N__48193),
            .I(n12421));
    CascadeMux I__10705 (
            .O(N__48190),
            .I(N__48187));
    InMux I__10704 (
            .O(N__48187),
            .I(N__48183));
    InMux I__10703 (
            .O(N__48186),
            .I(N__48180));
    LocalMux I__10702 (
            .O(N__48183),
            .I(N__48177));
    LocalMux I__10701 (
            .O(N__48180),
            .I(N__48173));
    Span4Mux_v I__10700 (
            .O(N__48177),
            .I(N__48170));
    InMux I__10699 (
            .O(N__48176),
            .I(N__48167));
    Odrv4 I__10698 (
            .O(N__48173),
            .I(n2822));
    Odrv4 I__10697 (
            .O(N__48170),
            .I(n2822));
    LocalMux I__10696 (
            .O(N__48167),
            .I(n2822));
    CascadeMux I__10695 (
            .O(N__48160),
            .I(N__48157));
    InMux I__10694 (
            .O(N__48157),
            .I(N__48154));
    LocalMux I__10693 (
            .O(N__48154),
            .I(N__48151));
    Span4Mux_h I__10692 (
            .O(N__48151),
            .I(N__48148));
    Odrv4 I__10691 (
            .O(N__48148),
            .I(n2889));
    InMux I__10690 (
            .O(N__48145),
            .I(n12422));
    CascadeMux I__10689 (
            .O(N__48142),
            .I(N__48139));
    InMux I__10688 (
            .O(N__48139),
            .I(N__48135));
    CascadeMux I__10687 (
            .O(N__48138),
            .I(N__48132));
    LocalMux I__10686 (
            .O(N__48135),
            .I(N__48129));
    InMux I__10685 (
            .O(N__48132),
            .I(N__48125));
    Span4Mux_h I__10684 (
            .O(N__48129),
            .I(N__48122));
    InMux I__10683 (
            .O(N__48128),
            .I(N__48119));
    LocalMux I__10682 (
            .O(N__48125),
            .I(n2821));
    Odrv4 I__10681 (
            .O(N__48122),
            .I(n2821));
    LocalMux I__10680 (
            .O(N__48119),
            .I(n2821));
    InMux I__10679 (
            .O(N__48112),
            .I(N__48109));
    LocalMux I__10678 (
            .O(N__48109),
            .I(N__48106));
    Odrv4 I__10677 (
            .O(N__48106),
            .I(n2888));
    InMux I__10676 (
            .O(N__48103),
            .I(n12423));
    CascadeMux I__10675 (
            .O(N__48100),
            .I(N__48096));
    CascadeMux I__10674 (
            .O(N__48099),
            .I(N__48093));
    InMux I__10673 (
            .O(N__48096),
            .I(N__48090));
    InMux I__10672 (
            .O(N__48093),
            .I(N__48087));
    LocalMux I__10671 (
            .O(N__48090),
            .I(N__48084));
    LocalMux I__10670 (
            .O(N__48087),
            .I(N__48081));
    Span4Mux_v I__10669 (
            .O(N__48084),
            .I(N__48077));
    Span4Mux_v I__10668 (
            .O(N__48081),
            .I(N__48074));
    InMux I__10667 (
            .O(N__48080),
            .I(N__48071));
    Sp12to4 I__10666 (
            .O(N__48077),
            .I(N__48064));
    Sp12to4 I__10665 (
            .O(N__48074),
            .I(N__48064));
    LocalMux I__10664 (
            .O(N__48071),
            .I(N__48064));
    Odrv12 I__10663 (
            .O(N__48064),
            .I(n2820));
    InMux I__10662 (
            .O(N__48061),
            .I(N__48058));
    LocalMux I__10661 (
            .O(N__48058),
            .I(N__48055));
    Odrv4 I__10660 (
            .O(N__48055),
            .I(n2887));
    InMux I__10659 (
            .O(N__48052),
            .I(n12424));
    CascadeMux I__10658 (
            .O(N__48049),
            .I(N__48046));
    InMux I__10657 (
            .O(N__48046),
            .I(N__48043));
    LocalMux I__10656 (
            .O(N__48043),
            .I(N__48039));
    InMux I__10655 (
            .O(N__48042),
            .I(N__48035));
    Span4Mux_h I__10654 (
            .O(N__48039),
            .I(N__48032));
    InMux I__10653 (
            .O(N__48038),
            .I(N__48029));
    LocalMux I__10652 (
            .O(N__48035),
            .I(n2819));
    Odrv4 I__10651 (
            .O(N__48032),
            .I(n2819));
    LocalMux I__10650 (
            .O(N__48029),
            .I(n2819));
    InMux I__10649 (
            .O(N__48022),
            .I(N__48019));
    LocalMux I__10648 (
            .O(N__48019),
            .I(N__48016));
    Span4Mux_h I__10647 (
            .O(N__48016),
            .I(N__48013));
    Odrv4 I__10646 (
            .O(N__48013),
            .I(n2886));
    InMux I__10645 (
            .O(N__48010),
            .I(n12425));
    InMux I__10644 (
            .O(N__48007),
            .I(N__48004));
    LocalMux I__10643 (
            .O(N__48004),
            .I(N__48000));
    InMux I__10642 (
            .O(N__48003),
            .I(N__47996));
    Span4Mux_v I__10641 (
            .O(N__48000),
            .I(N__47993));
    InMux I__10640 (
            .O(N__47999),
            .I(N__47990));
    LocalMux I__10639 (
            .O(N__47996),
            .I(n2818));
    Odrv4 I__10638 (
            .O(N__47993),
            .I(n2818));
    LocalMux I__10637 (
            .O(N__47990),
            .I(n2818));
    CascadeMux I__10636 (
            .O(N__47983),
            .I(N__47979));
    InMux I__10635 (
            .O(N__47982),
            .I(N__47976));
    InMux I__10634 (
            .O(N__47979),
            .I(N__47973));
    LocalMux I__10633 (
            .O(N__47976),
            .I(n2833));
    LocalMux I__10632 (
            .O(N__47973),
            .I(n2833));
    CascadeMux I__10631 (
            .O(N__47968),
            .I(N__47965));
    InMux I__10630 (
            .O(N__47965),
            .I(N__47962));
    LocalMux I__10629 (
            .O(N__47962),
            .I(n2900));
    InMux I__10628 (
            .O(N__47959),
            .I(n12411));
    CascadeMux I__10627 (
            .O(N__47956),
            .I(N__47953));
    InMux I__10626 (
            .O(N__47953),
            .I(N__47948));
    InMux I__10625 (
            .O(N__47952),
            .I(N__47943));
    InMux I__10624 (
            .O(N__47951),
            .I(N__47943));
    LocalMux I__10623 (
            .O(N__47948),
            .I(N__47940));
    LocalMux I__10622 (
            .O(N__47943),
            .I(n2832));
    Odrv4 I__10621 (
            .O(N__47940),
            .I(n2832));
    InMux I__10620 (
            .O(N__47935),
            .I(N__47932));
    LocalMux I__10619 (
            .O(N__47932),
            .I(n2899));
    InMux I__10618 (
            .O(N__47929),
            .I(n12412));
    CascadeMux I__10617 (
            .O(N__47926),
            .I(N__47923));
    InMux I__10616 (
            .O(N__47923),
            .I(N__47918));
    InMux I__10615 (
            .O(N__47922),
            .I(N__47913));
    InMux I__10614 (
            .O(N__47921),
            .I(N__47913));
    LocalMux I__10613 (
            .O(N__47918),
            .I(N__47910));
    LocalMux I__10612 (
            .O(N__47913),
            .I(n2831));
    Odrv4 I__10611 (
            .O(N__47910),
            .I(n2831));
    CascadeMux I__10610 (
            .O(N__47905),
            .I(N__47902));
    InMux I__10609 (
            .O(N__47902),
            .I(N__47899));
    LocalMux I__10608 (
            .O(N__47899),
            .I(n2898));
    InMux I__10607 (
            .O(N__47896),
            .I(n12413));
    CascadeMux I__10606 (
            .O(N__47893),
            .I(N__47890));
    InMux I__10605 (
            .O(N__47890),
            .I(N__47886));
    CascadeMux I__10604 (
            .O(N__47889),
            .I(N__47883));
    LocalMux I__10603 (
            .O(N__47886),
            .I(N__47879));
    InMux I__10602 (
            .O(N__47883),
            .I(N__47874));
    InMux I__10601 (
            .O(N__47882),
            .I(N__47874));
    Span4Mux_h I__10600 (
            .O(N__47879),
            .I(N__47871));
    LocalMux I__10599 (
            .O(N__47874),
            .I(n2830));
    Odrv4 I__10598 (
            .O(N__47871),
            .I(n2830));
    InMux I__10597 (
            .O(N__47866),
            .I(N__47863));
    LocalMux I__10596 (
            .O(N__47863),
            .I(N__47860));
    Odrv4 I__10595 (
            .O(N__47860),
            .I(n2897));
    InMux I__10594 (
            .O(N__47857),
            .I(n12414));
    CascadeMux I__10593 (
            .O(N__47854),
            .I(N__47851));
    InMux I__10592 (
            .O(N__47851),
            .I(N__47847));
    CascadeMux I__10591 (
            .O(N__47850),
            .I(N__47843));
    LocalMux I__10590 (
            .O(N__47847),
            .I(N__47840));
    InMux I__10589 (
            .O(N__47846),
            .I(N__47837));
    InMux I__10588 (
            .O(N__47843),
            .I(N__47834));
    Span4Mux_h I__10587 (
            .O(N__47840),
            .I(N__47831));
    LocalMux I__10586 (
            .O(N__47837),
            .I(n2829));
    LocalMux I__10585 (
            .O(N__47834),
            .I(n2829));
    Odrv4 I__10584 (
            .O(N__47831),
            .I(n2829));
    InMux I__10583 (
            .O(N__47824),
            .I(N__47821));
    LocalMux I__10582 (
            .O(N__47821),
            .I(n2896));
    InMux I__10581 (
            .O(N__47818),
            .I(n12415));
    CascadeMux I__10580 (
            .O(N__47815),
            .I(N__47811));
    InMux I__10579 (
            .O(N__47814),
            .I(N__47807));
    InMux I__10578 (
            .O(N__47811),
            .I(N__47804));
    InMux I__10577 (
            .O(N__47810),
            .I(N__47801));
    LocalMux I__10576 (
            .O(N__47807),
            .I(N__47796));
    LocalMux I__10575 (
            .O(N__47804),
            .I(N__47796));
    LocalMux I__10574 (
            .O(N__47801),
            .I(n2828));
    Odrv4 I__10573 (
            .O(N__47796),
            .I(n2828));
    InMux I__10572 (
            .O(N__47791),
            .I(N__47788));
    LocalMux I__10571 (
            .O(N__47788),
            .I(n2895));
    InMux I__10570 (
            .O(N__47785),
            .I(n12416));
    CascadeMux I__10569 (
            .O(N__47782),
            .I(N__47778));
    CascadeMux I__10568 (
            .O(N__47781),
            .I(N__47775));
    InMux I__10567 (
            .O(N__47778),
            .I(N__47772));
    InMux I__10566 (
            .O(N__47775),
            .I(N__47769));
    LocalMux I__10565 (
            .O(N__47772),
            .I(N__47766));
    LocalMux I__10564 (
            .O(N__47769),
            .I(N__47763));
    Span4Mux_h I__10563 (
            .O(N__47766),
            .I(N__47759));
    Span4Mux_h I__10562 (
            .O(N__47763),
            .I(N__47756));
    InMux I__10561 (
            .O(N__47762),
            .I(N__47753));
    Odrv4 I__10560 (
            .O(N__47759),
            .I(n2827));
    Odrv4 I__10559 (
            .O(N__47756),
            .I(n2827));
    LocalMux I__10558 (
            .O(N__47753),
            .I(n2827));
    InMux I__10557 (
            .O(N__47746),
            .I(N__47743));
    LocalMux I__10556 (
            .O(N__47743),
            .I(n2894));
    InMux I__10555 (
            .O(N__47740),
            .I(n12417));
    CascadeMux I__10554 (
            .O(N__47737),
            .I(N__47733));
    InMux I__10553 (
            .O(N__47736),
            .I(N__47730));
    InMux I__10552 (
            .O(N__47733),
            .I(N__47727));
    LocalMux I__10551 (
            .O(N__47730),
            .I(N__47721));
    LocalMux I__10550 (
            .O(N__47727),
            .I(N__47721));
    InMux I__10549 (
            .O(N__47726),
            .I(N__47718));
    Span4Mux_v I__10548 (
            .O(N__47721),
            .I(N__47715));
    LocalMux I__10547 (
            .O(N__47718),
            .I(N__47712));
    Odrv4 I__10546 (
            .O(N__47715),
            .I(n2826));
    Odrv4 I__10545 (
            .O(N__47712),
            .I(n2826));
    CascadeMux I__10544 (
            .O(N__47707),
            .I(N__47704));
    InMux I__10543 (
            .O(N__47704),
            .I(N__47701));
    LocalMux I__10542 (
            .O(N__47701),
            .I(n2893));
    InMux I__10541 (
            .O(N__47698),
            .I(bfn_15_21_0_));
    InMux I__10540 (
            .O(N__47695),
            .I(N__47692));
    LocalMux I__10539 (
            .O(N__47692),
            .I(N__47689));
    Span4Mux_h I__10538 (
            .O(N__47689),
            .I(N__47686));
    Odrv4 I__10537 (
            .O(N__47686),
            .I(n2801));
    InMux I__10536 (
            .O(N__47683),
            .I(N__47679));
    InMux I__10535 (
            .O(N__47682),
            .I(N__47675));
    LocalMux I__10534 (
            .O(N__47679),
            .I(N__47672));
    InMux I__10533 (
            .O(N__47678),
            .I(N__47669));
    LocalMux I__10532 (
            .O(N__47675),
            .I(N__47666));
    Span4Mux_v I__10531 (
            .O(N__47672),
            .I(N__47661));
    LocalMux I__10530 (
            .O(N__47669),
            .I(N__47661));
    Span4Mux_h I__10529 (
            .O(N__47666),
            .I(N__47658));
    Span4Mux_h I__10528 (
            .O(N__47661),
            .I(N__47655));
    Span4Mux_h I__10527 (
            .O(N__47658),
            .I(N__47652));
    Span4Mux_v I__10526 (
            .O(N__47655),
            .I(N__47649));
    Odrv4 I__10525 (
            .O(N__47652),
            .I(n313));
    Odrv4 I__10524 (
            .O(N__47649),
            .I(n313));
    CascadeMux I__10523 (
            .O(N__47644),
            .I(N__47641));
    InMux I__10522 (
            .O(N__47641),
            .I(N__47638));
    LocalMux I__10521 (
            .O(N__47638),
            .I(N__47634));
    InMux I__10520 (
            .O(N__47637),
            .I(N__47631));
    Span4Mux_v I__10519 (
            .O(N__47634),
            .I(N__47620));
    LocalMux I__10518 (
            .O(N__47631),
            .I(N__47620));
    InMux I__10517 (
            .O(N__47630),
            .I(N__47617));
    InMux I__10516 (
            .O(N__47629),
            .I(N__47613));
    InMux I__10515 (
            .O(N__47628),
            .I(N__47608));
    InMux I__10514 (
            .O(N__47627),
            .I(N__47608));
    CascadeMux I__10513 (
            .O(N__47626),
            .I(N__47599));
    CascadeMux I__10512 (
            .O(N__47625),
            .I(N__47596));
    Span4Mux_v I__10511 (
            .O(N__47620),
            .I(N__47589));
    LocalMux I__10510 (
            .O(N__47617),
            .I(N__47589));
    InMux I__10509 (
            .O(N__47616),
            .I(N__47586));
    LocalMux I__10508 (
            .O(N__47613),
            .I(N__47581));
    LocalMux I__10507 (
            .O(N__47608),
            .I(N__47581));
    CascadeMux I__10506 (
            .O(N__47607),
            .I(N__47578));
    CascadeMux I__10505 (
            .O(N__47606),
            .I(N__47574));
    CascadeMux I__10504 (
            .O(N__47605),
            .I(N__47569));
    CascadeMux I__10503 (
            .O(N__47604),
            .I(N__47564));
    CascadeMux I__10502 (
            .O(N__47603),
            .I(N__47559));
    CascadeMux I__10501 (
            .O(N__47602),
            .I(N__47555));
    InMux I__10500 (
            .O(N__47599),
            .I(N__47549));
    InMux I__10499 (
            .O(N__47596),
            .I(N__47549));
    InMux I__10498 (
            .O(N__47595),
            .I(N__47546));
    InMux I__10497 (
            .O(N__47594),
            .I(N__47543));
    Span4Mux_v I__10496 (
            .O(N__47589),
            .I(N__47540));
    LocalMux I__10495 (
            .O(N__47586),
            .I(N__47537));
    Span4Mux_v I__10494 (
            .O(N__47581),
            .I(N__47534));
    InMux I__10493 (
            .O(N__47578),
            .I(N__47523));
    InMux I__10492 (
            .O(N__47577),
            .I(N__47523));
    InMux I__10491 (
            .O(N__47574),
            .I(N__47523));
    InMux I__10490 (
            .O(N__47573),
            .I(N__47523));
    InMux I__10489 (
            .O(N__47572),
            .I(N__47523));
    InMux I__10488 (
            .O(N__47569),
            .I(N__47516));
    InMux I__10487 (
            .O(N__47568),
            .I(N__47516));
    InMux I__10486 (
            .O(N__47567),
            .I(N__47516));
    InMux I__10485 (
            .O(N__47564),
            .I(N__47511));
    InMux I__10484 (
            .O(N__47563),
            .I(N__47511));
    InMux I__10483 (
            .O(N__47562),
            .I(N__47500));
    InMux I__10482 (
            .O(N__47559),
            .I(N__47500));
    InMux I__10481 (
            .O(N__47558),
            .I(N__47500));
    InMux I__10480 (
            .O(N__47555),
            .I(N__47500));
    InMux I__10479 (
            .O(N__47554),
            .I(N__47500));
    LocalMux I__10478 (
            .O(N__47549),
            .I(N__47495));
    LocalMux I__10477 (
            .O(N__47546),
            .I(N__47495));
    LocalMux I__10476 (
            .O(N__47543),
            .I(N__47488));
    Span4Mux_h I__10475 (
            .O(N__47540),
            .I(N__47488));
    Span4Mux_h I__10474 (
            .O(N__47537),
            .I(N__47488));
    Odrv4 I__10473 (
            .O(N__47534),
            .I(n2742));
    LocalMux I__10472 (
            .O(N__47523),
            .I(n2742));
    LocalMux I__10471 (
            .O(N__47516),
            .I(n2742));
    LocalMux I__10470 (
            .O(N__47511),
            .I(n2742));
    LocalMux I__10469 (
            .O(N__47500),
            .I(n2742));
    Odrv4 I__10468 (
            .O(N__47495),
            .I(n2742));
    Odrv4 I__10467 (
            .O(N__47488),
            .I(n2742));
    CascadeMux I__10466 (
            .O(N__47473),
            .I(n2833_cascade_));
    InMux I__10465 (
            .O(N__47470),
            .I(N__47467));
    LocalMux I__10464 (
            .O(N__47467),
            .I(n11756));
    CascadeMux I__10463 (
            .O(N__47464),
            .I(N__47461));
    InMux I__10462 (
            .O(N__47461),
            .I(N__47457));
    InMux I__10461 (
            .O(N__47460),
            .I(N__47454));
    LocalMux I__10460 (
            .O(N__47457),
            .I(N__47451));
    LocalMux I__10459 (
            .O(N__47454),
            .I(N__47448));
    Span4Mux_v I__10458 (
            .O(N__47451),
            .I(N__47445));
    Span4Mux_v I__10457 (
            .O(N__47448),
            .I(N__47442));
    Span4Mux_h I__10456 (
            .O(N__47445),
            .I(N__47439));
    Odrv4 I__10455 (
            .O(N__47442),
            .I(n2932));
    Odrv4 I__10454 (
            .O(N__47439),
            .I(n2932));
    InMux I__10453 (
            .O(N__47434),
            .I(N__47431));
    LocalMux I__10452 (
            .O(N__47431),
            .I(N__47427));
    CascadeMux I__10451 (
            .O(N__47430),
            .I(N__47424));
    Span4Mux_v I__10450 (
            .O(N__47427),
            .I(N__47421));
    InMux I__10449 (
            .O(N__47424),
            .I(N__47418));
    Span4Mux_h I__10448 (
            .O(N__47421),
            .I(N__47415));
    LocalMux I__10447 (
            .O(N__47418),
            .I(n315));
    Odrv4 I__10446 (
            .O(N__47415),
            .I(n315));
    CascadeMux I__10445 (
            .O(N__47410),
            .I(n2932_cascade_));
    CascadeMux I__10444 (
            .O(N__47407),
            .I(N__47403));
    InMux I__10443 (
            .O(N__47406),
            .I(N__47400));
    InMux I__10442 (
            .O(N__47403),
            .I(N__47397));
    LocalMux I__10441 (
            .O(N__47400),
            .I(N__47391));
    LocalMux I__10440 (
            .O(N__47397),
            .I(N__47391));
    InMux I__10439 (
            .O(N__47396),
            .I(N__47388));
    Span4Mux_v I__10438 (
            .O(N__47391),
            .I(N__47385));
    LocalMux I__10437 (
            .O(N__47388),
            .I(N__47382));
    Odrv4 I__10436 (
            .O(N__47385),
            .I(n2933));
    Odrv4 I__10435 (
            .O(N__47382),
            .I(n2933));
    CascadeMux I__10434 (
            .O(N__47377),
            .I(N__47373));
    InMux I__10433 (
            .O(N__47376),
            .I(N__47370));
    InMux I__10432 (
            .O(N__47373),
            .I(N__47367));
    LocalMux I__10431 (
            .O(N__47370),
            .I(N__47364));
    LocalMux I__10430 (
            .O(N__47367),
            .I(N__47361));
    Span4Mux_v I__10429 (
            .O(N__47364),
            .I(N__47356));
    Span4Mux_h I__10428 (
            .O(N__47361),
            .I(N__47356));
    Span4Mux_h I__10427 (
            .O(N__47356),
            .I(N__47353));
    Odrv4 I__10426 (
            .O(N__47353),
            .I(n2930));
    CascadeMux I__10425 (
            .O(N__47350),
            .I(N__47347));
    InMux I__10424 (
            .O(N__47347),
            .I(N__47343));
    InMux I__10423 (
            .O(N__47346),
            .I(N__47340));
    LocalMux I__10422 (
            .O(N__47343),
            .I(N__47337));
    LocalMux I__10421 (
            .O(N__47340),
            .I(N__47334));
    Span4Mux_v I__10420 (
            .O(N__47337),
            .I(N__47330));
    Span4Mux_v I__10419 (
            .O(N__47334),
            .I(N__47327));
    InMux I__10418 (
            .O(N__47333),
            .I(N__47324));
    Span4Mux_h I__10417 (
            .O(N__47330),
            .I(N__47321));
    Odrv4 I__10416 (
            .O(N__47327),
            .I(n2931));
    LocalMux I__10415 (
            .O(N__47324),
            .I(n2931));
    Odrv4 I__10414 (
            .O(N__47321),
            .I(n2931));
    CascadeMux I__10413 (
            .O(N__47314),
            .I(N__47310));
    InMux I__10412 (
            .O(N__47313),
            .I(N__47307));
    InMux I__10411 (
            .O(N__47310),
            .I(N__47304));
    LocalMux I__10410 (
            .O(N__47307),
            .I(N__47300));
    LocalMux I__10409 (
            .O(N__47304),
            .I(N__47297));
    InMux I__10408 (
            .O(N__47303),
            .I(N__47294));
    Span4Mux_h I__10407 (
            .O(N__47300),
            .I(N__47289));
    Span4Mux_h I__10406 (
            .O(N__47297),
            .I(N__47289));
    LocalMux I__10405 (
            .O(N__47294),
            .I(n2929));
    Odrv4 I__10404 (
            .O(N__47289),
            .I(n2929));
    CascadeMux I__10403 (
            .O(N__47284),
            .I(n2930_cascade_));
    InMux I__10402 (
            .O(N__47281),
            .I(N__47278));
    LocalMux I__10401 (
            .O(N__47278),
            .I(n11662));
    CascadeMux I__10400 (
            .O(N__47275),
            .I(N__47272));
    InMux I__10399 (
            .O(N__47272),
            .I(N__47269));
    LocalMux I__10398 (
            .O(N__47269),
            .I(N__47266));
    Span4Mux_h I__10397 (
            .O(N__47266),
            .I(N__47263));
    Odrv4 I__10396 (
            .O(N__47263),
            .I(n13417));
    InMux I__10395 (
            .O(N__47260),
            .I(N__47257));
    LocalMux I__10394 (
            .O(N__47257),
            .I(N__47253));
    InMux I__10393 (
            .O(N__47256),
            .I(N__47250));
    Span4Mux_v I__10392 (
            .O(N__47253),
            .I(N__47244));
    LocalMux I__10391 (
            .O(N__47250),
            .I(N__47244));
    InMux I__10390 (
            .O(N__47249),
            .I(N__47241));
    Span4Mux_h I__10389 (
            .O(N__47244),
            .I(N__47236));
    LocalMux I__10388 (
            .O(N__47241),
            .I(N__47236));
    Span4Mux_v I__10387 (
            .O(N__47236),
            .I(N__47233));
    Span4Mux_h I__10386 (
            .O(N__47233),
            .I(N__47230));
    Odrv4 I__10385 (
            .O(N__47230),
            .I(n314));
    InMux I__10384 (
            .O(N__47227),
            .I(N__47224));
    LocalMux I__10383 (
            .O(N__47224),
            .I(N__47221));
    Span4Mux_h I__10382 (
            .O(N__47221),
            .I(N__47218));
    Odrv4 I__10381 (
            .O(N__47218),
            .I(n2901));
    InMux I__10380 (
            .O(N__47215),
            .I(bfn_15_20_0_));
    InMux I__10379 (
            .O(N__47212),
            .I(N__47207));
    InMux I__10378 (
            .O(N__47211),
            .I(N__47204));
    InMux I__10377 (
            .O(N__47210),
            .I(N__47201));
    LocalMux I__10376 (
            .O(N__47207),
            .I(n31_adj_624));
    LocalMux I__10375 (
            .O(N__47204),
            .I(n31_adj_624));
    LocalMux I__10374 (
            .O(N__47201),
            .I(n31_adj_624));
    InMux I__10373 (
            .O(N__47194),
            .I(N__47191));
    LocalMux I__10372 (
            .O(N__47191),
            .I(N__47188));
    Span4Mux_s2_v I__10371 (
            .O(N__47188),
            .I(N__47185));
    Odrv4 I__10370 (
            .O(N__47185),
            .I(n14728));
    CascadeMux I__10369 (
            .O(N__47182),
            .I(n33_adj_625_cascade_));
    InMux I__10368 (
            .O(N__47179),
            .I(N__47175));
    InMux I__10367 (
            .O(N__47178),
            .I(N__47172));
    LocalMux I__10366 (
            .O(N__47175),
            .I(N__47166));
    LocalMux I__10365 (
            .O(N__47172),
            .I(N__47166));
    InMux I__10364 (
            .O(N__47171),
            .I(N__47163));
    Odrv4 I__10363 (
            .O(N__47166),
            .I(n29_adj_622));
    LocalMux I__10362 (
            .O(N__47163),
            .I(n29_adj_622));
    InMux I__10361 (
            .O(N__47158),
            .I(N__47155));
    LocalMux I__10360 (
            .O(N__47155),
            .I(n14724));
    InMux I__10359 (
            .O(N__47152),
            .I(N__47149));
    LocalMux I__10358 (
            .O(N__47149),
            .I(N__47145));
    InMux I__10357 (
            .O(N__47148),
            .I(N__47142));
    Sp12to4 I__10356 (
            .O(N__47145),
            .I(N__47137));
    LocalMux I__10355 (
            .O(N__47142),
            .I(N__47137));
    Odrv12 I__10354 (
            .O(N__47137),
            .I(duty_17));
    InMux I__10353 (
            .O(N__47134),
            .I(N__47131));
    LocalMux I__10352 (
            .O(N__47131),
            .I(N__47128));
    Odrv4 I__10351 (
            .O(N__47128),
            .I(n8_adj_574));
    InMux I__10350 (
            .O(N__47125),
            .I(N__47122));
    LocalMux I__10349 (
            .O(N__47122),
            .I(n28_adj_597));
    InMux I__10348 (
            .O(N__47119),
            .I(N__47116));
    LocalMux I__10347 (
            .O(N__47116),
            .I(n31_adj_594));
    CascadeMux I__10346 (
            .O(N__47113),
            .I(n32_adj_593_cascade_));
    InMux I__10345 (
            .O(N__47110),
            .I(N__47107));
    LocalMux I__10344 (
            .O(N__47107),
            .I(N__47104));
    Span4Mux_v I__10343 (
            .O(N__47104),
            .I(N__47099));
    InMux I__10342 (
            .O(N__47103),
            .I(N__47094));
    InMux I__10341 (
            .O(N__47102),
            .I(N__47094));
    Span4Mux_h I__10340 (
            .O(N__47099),
            .I(N__47091));
    LocalMux I__10339 (
            .O(N__47094),
            .I(N__47088));
    Span4Mux_v I__10338 (
            .O(N__47091),
            .I(N__47085));
    Span4Mux_h I__10337 (
            .O(N__47088),
            .I(N__47082));
    Odrv4 I__10336 (
            .O(N__47085),
            .I(n2910));
    Odrv4 I__10335 (
            .O(N__47082),
            .I(n2910));
    InMux I__10334 (
            .O(N__47077),
            .I(N__47074));
    LocalMux I__10333 (
            .O(N__47074),
            .I(n30_adj_595));
    InMux I__10332 (
            .O(N__47071),
            .I(N__47068));
    LocalMux I__10331 (
            .O(N__47068),
            .I(n29_adj_596));
    InMux I__10330 (
            .O(N__47065),
            .I(N__47062));
    LocalMux I__10329 (
            .O(N__47062),
            .I(N__47058));
    InMux I__10328 (
            .O(N__47061),
            .I(N__47055));
    Span4Mux_h I__10327 (
            .O(N__47058),
            .I(N__47052));
    LocalMux I__10326 (
            .O(N__47055),
            .I(N__47049));
    Odrv4 I__10325 (
            .O(N__47052),
            .I(duty_20));
    Odrv4 I__10324 (
            .O(N__47049),
            .I(duty_20));
    InMux I__10323 (
            .O(N__47044),
            .I(N__47041));
    LocalMux I__10322 (
            .O(N__47041),
            .I(n5_adj_571));
    CascadeMux I__10321 (
            .O(N__47038),
            .I(N__47035));
    InMux I__10320 (
            .O(N__47035),
            .I(N__47032));
    LocalMux I__10319 (
            .O(N__47032),
            .I(N__47026));
    InMux I__10318 (
            .O(N__47031),
            .I(N__47021));
    InMux I__10317 (
            .O(N__47030),
            .I(N__47021));
    InMux I__10316 (
            .O(N__47029),
            .I(N__47018));
    Span4Mux_h I__10315 (
            .O(N__47026),
            .I(N__47015));
    LocalMux I__10314 (
            .O(N__47021),
            .I(N__47012));
    LocalMux I__10313 (
            .O(N__47018),
            .I(pwm_counter_7));
    Odrv4 I__10312 (
            .O(N__47015),
            .I(pwm_counter_7));
    Odrv4 I__10311 (
            .O(N__47012),
            .I(pwm_counter_7));
    InMux I__10310 (
            .O(N__47005),
            .I(N__47002));
    LocalMux I__10309 (
            .O(N__47002),
            .I(N__46999));
    Span4Mux_h I__10308 (
            .O(N__46999),
            .I(N__46996));
    Odrv4 I__10307 (
            .O(N__46996),
            .I(n10_adj_609));
    CascadeMux I__10306 (
            .O(N__46993),
            .I(n14722_cascade_));
    CascadeMux I__10305 (
            .O(N__46990),
            .I(n14876_cascade_));
    InMux I__10304 (
            .O(N__46987),
            .I(N__46984));
    LocalMux I__10303 (
            .O(N__46984),
            .I(n14886));
    InMux I__10302 (
            .O(N__46981),
            .I(N__46977));
    InMux I__10301 (
            .O(N__46980),
            .I(N__46974));
    LocalMux I__10300 (
            .O(N__46977),
            .I(pwm_setpoint_15));
    LocalMux I__10299 (
            .O(N__46974),
            .I(pwm_setpoint_15));
    InMux I__10298 (
            .O(N__46969),
            .I(N__46966));
    LocalMux I__10297 (
            .O(N__46966),
            .I(n14841));
    InMux I__10296 (
            .O(N__46963),
            .I(N__46960));
    LocalMux I__10295 (
            .O(N__46960),
            .I(n14781));
    InMux I__10294 (
            .O(N__46957),
            .I(N__46954));
    LocalMux I__10293 (
            .O(N__46954),
            .I(N__46951));
    Odrv4 I__10292 (
            .O(N__46951),
            .I(pwm_setpoint_23_N_171_7));
    InMux I__10291 (
            .O(N__46948),
            .I(N__46944));
    InMux I__10290 (
            .O(N__46947),
            .I(N__46941));
    LocalMux I__10289 (
            .O(N__46944),
            .I(N__46938));
    LocalMux I__10288 (
            .O(N__46941),
            .I(N__46935));
    Span4Mux_h I__10287 (
            .O(N__46938),
            .I(N__46932));
    Odrv12 I__10286 (
            .O(N__46935),
            .I(duty_7));
    Odrv4 I__10285 (
            .O(N__46932),
            .I(duty_7));
    InMux I__10284 (
            .O(N__46927),
            .I(N__46923));
    InMux I__10283 (
            .O(N__46926),
            .I(N__46919));
    LocalMux I__10282 (
            .O(N__46923),
            .I(N__46916));
    InMux I__10281 (
            .O(N__46922),
            .I(N__46913));
    LocalMux I__10280 (
            .O(N__46919),
            .I(pwm_setpoint_7));
    Odrv4 I__10279 (
            .O(N__46916),
            .I(pwm_setpoint_7));
    LocalMux I__10278 (
            .O(N__46913),
            .I(pwm_setpoint_7));
    InMux I__10277 (
            .O(N__46906),
            .I(N__46902));
    InMux I__10276 (
            .O(N__46905),
            .I(N__46899));
    LocalMux I__10275 (
            .O(N__46902),
            .I(pwm_setpoint_17));
    LocalMux I__10274 (
            .O(N__46899),
            .I(pwm_setpoint_17));
    CascadeMux I__10273 (
            .O(N__46894),
            .I(n12_adj_611_cascade_));
    CascadeMux I__10272 (
            .O(N__46891),
            .I(N__46888));
    InMux I__10271 (
            .O(N__46888),
            .I(N__46882));
    InMux I__10270 (
            .O(N__46887),
            .I(N__46877));
    InMux I__10269 (
            .O(N__46886),
            .I(N__46877));
    InMux I__10268 (
            .O(N__46885),
            .I(N__46874));
    LocalMux I__10267 (
            .O(N__46882),
            .I(n35));
    LocalMux I__10266 (
            .O(N__46877),
            .I(n35));
    LocalMux I__10265 (
            .O(N__46874),
            .I(n35));
    InMux I__10264 (
            .O(N__46867),
            .I(N__46864));
    LocalMux I__10263 (
            .O(N__46864),
            .I(n30_adj_623));
    InMux I__10262 (
            .O(N__46861),
            .I(N__46854));
    InMux I__10261 (
            .O(N__46860),
            .I(N__46854));
    InMux I__10260 (
            .O(N__46859),
            .I(N__46851));
    LocalMux I__10259 (
            .O(N__46854),
            .I(N__46848));
    LocalMux I__10258 (
            .O(N__46851),
            .I(pwm_setpoint_16));
    Odrv4 I__10257 (
            .O(N__46848),
            .I(pwm_setpoint_16));
    CascadeMux I__10256 (
            .O(N__46843),
            .I(N__46837));
    InMux I__10255 (
            .O(N__46842),
            .I(N__46834));
    InMux I__10254 (
            .O(N__46841),
            .I(N__46829));
    InMux I__10253 (
            .O(N__46840),
            .I(N__46829));
    InMux I__10252 (
            .O(N__46837),
            .I(N__46825));
    LocalMux I__10251 (
            .O(N__46834),
            .I(N__46822));
    LocalMux I__10250 (
            .O(N__46829),
            .I(N__46819));
    InMux I__10249 (
            .O(N__46828),
            .I(N__46816));
    LocalMux I__10248 (
            .O(N__46825),
            .I(N__46809));
    Span4Mux_h I__10247 (
            .O(N__46822),
            .I(N__46809));
    Span4Mux_s1_v I__10246 (
            .O(N__46819),
            .I(N__46809));
    LocalMux I__10245 (
            .O(N__46816),
            .I(pwm_counter_16));
    Odrv4 I__10244 (
            .O(N__46809),
            .I(pwm_counter_16));
    InMux I__10243 (
            .O(N__46804),
            .I(N__46801));
    LocalMux I__10242 (
            .O(N__46801),
            .I(N__46798));
    Odrv4 I__10241 (
            .O(N__46798),
            .I(n33_adj_625));
    InMux I__10240 (
            .O(N__46795),
            .I(N__46792));
    LocalMux I__10239 (
            .O(N__46792),
            .I(N__46788));
    InMux I__10238 (
            .O(N__46791),
            .I(N__46785));
    Span4Mux_h I__10237 (
            .O(N__46788),
            .I(N__46782));
    LocalMux I__10236 (
            .O(N__46785),
            .I(N__46779));
    Odrv4 I__10235 (
            .O(N__46782),
            .I(duty_12));
    Odrv4 I__10234 (
            .O(N__46779),
            .I(duty_12));
    InMux I__10233 (
            .O(N__46774),
            .I(N__46771));
    LocalMux I__10232 (
            .O(N__46771),
            .I(n13_adj_579));
    InMux I__10231 (
            .O(N__46768),
            .I(N__46763));
    InMux I__10230 (
            .O(N__46767),
            .I(N__46760));
    InMux I__10229 (
            .O(N__46766),
            .I(N__46757));
    LocalMux I__10228 (
            .O(N__46763),
            .I(N__46754));
    LocalMux I__10227 (
            .O(N__46760),
            .I(pwm_counter_14));
    LocalMux I__10226 (
            .O(N__46757),
            .I(pwm_counter_14));
    Odrv12 I__10225 (
            .O(N__46754),
            .I(pwm_counter_14));
    InMux I__10224 (
            .O(N__46747),
            .I(N__46744));
    LocalMux I__10223 (
            .O(N__46744),
            .I(N__46739));
    InMux I__10222 (
            .O(N__46743),
            .I(N__46736));
    InMux I__10221 (
            .O(N__46742),
            .I(N__46733));
    Span4Mux_s2_v I__10220 (
            .O(N__46739),
            .I(N__46730));
    LocalMux I__10219 (
            .O(N__46736),
            .I(N__46727));
    LocalMux I__10218 (
            .O(N__46733),
            .I(pwm_counter_13));
    Odrv4 I__10217 (
            .O(N__46730),
            .I(pwm_counter_13));
    Odrv4 I__10216 (
            .O(N__46727),
            .I(pwm_counter_13));
    CascadeMux I__10215 (
            .O(N__46720),
            .I(N__46717));
    InMux I__10214 (
            .O(N__46717),
            .I(N__46714));
    LocalMux I__10213 (
            .O(N__46714),
            .I(N__46710));
    InMux I__10212 (
            .O(N__46713),
            .I(N__46707));
    Span4Mux_s2_v I__10211 (
            .O(N__46710),
            .I(N__46704));
    LocalMux I__10210 (
            .O(N__46707),
            .I(N__46701));
    Odrv4 I__10209 (
            .O(N__46704),
            .I(n27_adj_621));
    Odrv4 I__10208 (
            .O(N__46701),
            .I(n27_adj_621));
    InMux I__10207 (
            .O(N__46696),
            .I(N__46690));
    InMux I__10206 (
            .O(N__46695),
            .I(N__46690));
    LocalMux I__10205 (
            .O(N__46690),
            .I(pwm_setpoint_13));
    CascadeMux I__10204 (
            .O(N__46687),
            .I(n27_adj_621_cascade_));
    InMux I__10203 (
            .O(N__46684),
            .I(N__46681));
    LocalMux I__10202 (
            .O(N__46681),
            .I(n4_adj_605));
    InMux I__10201 (
            .O(N__46678),
            .I(N__46672));
    InMux I__10200 (
            .O(N__46677),
            .I(N__46672));
    LocalMux I__10199 (
            .O(N__46672),
            .I(pwm_setpoint_14));
    CascadeMux I__10198 (
            .O(N__46669),
            .I(n14840_cascade_));
    InMux I__10197 (
            .O(N__46666),
            .I(N__46662));
    InMux I__10196 (
            .O(N__46665),
            .I(N__46659));
    LocalMux I__10195 (
            .O(N__46662),
            .I(N__46654));
    LocalMux I__10194 (
            .O(N__46659),
            .I(N__46654));
    Odrv4 I__10193 (
            .O(N__46654),
            .I(duty_22));
    InMux I__10192 (
            .O(N__46651),
            .I(N__46648));
    LocalMux I__10191 (
            .O(N__46648),
            .I(n3_adj_569));
    InMux I__10190 (
            .O(N__46645),
            .I(N__46642));
    LocalMux I__10189 (
            .O(N__46642),
            .I(n9_adj_575));
    InMux I__10188 (
            .O(N__46639),
            .I(N__46633));
    InMux I__10187 (
            .O(N__46638),
            .I(N__46633));
    LocalMux I__10186 (
            .O(N__46633),
            .I(N__46630));
    Odrv4 I__10185 (
            .O(N__46630),
            .I(duty_16));
    InMux I__10184 (
            .O(N__46627),
            .I(N__46624));
    LocalMux I__10183 (
            .O(N__46624),
            .I(pwm_setpoint_23_N_171_16));
    InMux I__10182 (
            .O(N__46621),
            .I(N__46618));
    LocalMux I__10181 (
            .O(N__46618),
            .I(N__46615));
    Span4Mux_h I__10180 (
            .O(N__46615),
            .I(N__46612));
    Odrv4 I__10179 (
            .O(N__46612),
            .I(n3));
    InMux I__10178 (
            .O(N__46609),
            .I(n12094));
    InMux I__10177 (
            .O(N__46606),
            .I(N__46603));
    LocalMux I__10176 (
            .O(N__46603),
            .I(N__46600));
    Odrv12 I__10175 (
            .O(N__46600),
            .I(n2));
    InMux I__10174 (
            .O(N__46597),
            .I(n12095));
    InMux I__10173 (
            .O(N__46594),
            .I(N__46591));
    LocalMux I__10172 (
            .O(N__46591),
            .I(pwm_setpoint_23_N_171_13));
    InMux I__10171 (
            .O(N__46588),
            .I(N__46585));
    LocalMux I__10170 (
            .O(N__46585),
            .I(N__46581));
    InMux I__10169 (
            .O(N__46584),
            .I(N__46578));
    Span4Mux_s2_v I__10168 (
            .O(N__46581),
            .I(N__46573));
    LocalMux I__10167 (
            .O(N__46578),
            .I(N__46573));
    Odrv4 I__10166 (
            .O(N__46573),
            .I(duty_15));
    InMux I__10165 (
            .O(N__46570),
            .I(N__46567));
    LocalMux I__10164 (
            .O(N__46567),
            .I(n10_adj_576));
    InMux I__10163 (
            .O(N__46564),
            .I(N__46561));
    LocalMux I__10162 (
            .O(N__46561),
            .I(N__46557));
    InMux I__10161 (
            .O(N__46560),
            .I(N__46554));
    Odrv4 I__10160 (
            .O(N__46557),
            .I(duty_14));
    LocalMux I__10159 (
            .O(N__46554),
            .I(duty_14));
    InMux I__10158 (
            .O(N__46549),
            .I(N__46546));
    LocalMux I__10157 (
            .O(N__46546),
            .I(pwm_setpoint_23_N_171_14));
    InMux I__10156 (
            .O(N__46543),
            .I(N__46539));
    InMux I__10155 (
            .O(N__46542),
            .I(N__46536));
    LocalMux I__10154 (
            .O(N__46539),
            .I(N__46533));
    LocalMux I__10153 (
            .O(N__46536),
            .I(pwm_counter_1));
    Odrv4 I__10152 (
            .O(N__46533),
            .I(pwm_counter_1));
    CascadeMux I__10151 (
            .O(N__46528),
            .I(N__46525));
    InMux I__10150 (
            .O(N__46525),
            .I(N__46521));
    InMux I__10149 (
            .O(N__46524),
            .I(N__46518));
    LocalMux I__10148 (
            .O(N__46521),
            .I(N__46515));
    LocalMux I__10147 (
            .O(N__46518),
            .I(pwm_counter_0));
    Odrv4 I__10146 (
            .O(N__46515),
            .I(pwm_counter_0));
    InMux I__10145 (
            .O(N__46510),
            .I(N__46507));
    LocalMux I__10144 (
            .O(N__46507),
            .I(n16_adj_582));
    InMux I__10143 (
            .O(N__46504),
            .I(N__46500));
    InMux I__10142 (
            .O(N__46503),
            .I(N__46497));
    LocalMux I__10141 (
            .O(N__46500),
            .I(N__46492));
    LocalMux I__10140 (
            .O(N__46497),
            .I(N__46492));
    Odrv4 I__10139 (
            .O(N__46492),
            .I(duty_13));
    InMux I__10138 (
            .O(N__46489),
            .I(N__46486));
    LocalMux I__10137 (
            .O(N__46486),
            .I(n12_adj_578));
    InMux I__10136 (
            .O(N__46483),
            .I(N__46480));
    LocalMux I__10135 (
            .O(N__46480),
            .I(pwm_setpoint_23_N_171_0));
    InMux I__10134 (
            .O(N__46477),
            .I(N__46474));
    LocalMux I__10133 (
            .O(N__46474),
            .I(N__46470));
    InMux I__10132 (
            .O(N__46473),
            .I(N__46467));
    Odrv12 I__10131 (
            .O(N__46470),
            .I(duty_0));
    LocalMux I__10130 (
            .O(N__46467),
            .I(duty_0));
    InMux I__10129 (
            .O(N__46462),
            .I(N__46459));
    LocalMux I__10128 (
            .O(N__46459),
            .I(pwm_setpoint_0));
    CascadeMux I__10127 (
            .O(N__46456),
            .I(N__46453));
    InMux I__10126 (
            .O(N__46453),
            .I(N__46450));
    LocalMux I__10125 (
            .O(N__46450),
            .I(N__46447));
    Odrv12 I__10124 (
            .O(N__46447),
            .I(n11_adj_559));
    InMux I__10123 (
            .O(N__46444),
            .I(n12086));
    InMux I__10122 (
            .O(N__46441),
            .I(N__46438));
    LocalMux I__10121 (
            .O(N__46438),
            .I(N__46435));
    Span4Mux_h I__10120 (
            .O(N__46435),
            .I(N__46432));
    Odrv4 I__10119 (
            .O(N__46432),
            .I(n10_adj_560));
    InMux I__10118 (
            .O(N__46429),
            .I(n12087));
    CascadeMux I__10117 (
            .O(N__46426),
            .I(N__46423));
    InMux I__10116 (
            .O(N__46423),
            .I(N__46420));
    LocalMux I__10115 (
            .O(N__46420),
            .I(N__46417));
    Odrv4 I__10114 (
            .O(N__46417),
            .I(n9_adj_561));
    InMux I__10113 (
            .O(N__46414),
            .I(bfn_14_28_0_));
    InMux I__10112 (
            .O(N__46411),
            .I(N__46408));
    LocalMux I__10111 (
            .O(N__46408),
            .I(N__46405));
    Odrv12 I__10110 (
            .O(N__46405),
            .I(n8_adj_562));
    InMux I__10109 (
            .O(N__46402),
            .I(n12089));
    InMux I__10108 (
            .O(N__46399),
            .I(N__46396));
    LocalMux I__10107 (
            .O(N__46396),
            .I(N__46393));
    Odrv12 I__10106 (
            .O(N__46393),
            .I(n7_adj_563));
    InMux I__10105 (
            .O(N__46390),
            .I(n12090));
    InMux I__10104 (
            .O(N__46387),
            .I(N__46384));
    LocalMux I__10103 (
            .O(N__46384),
            .I(N__46381));
    Span4Mux_v I__10102 (
            .O(N__46381),
            .I(N__46378));
    Odrv4 I__10101 (
            .O(N__46378),
            .I(n6_adj_564));
    InMux I__10100 (
            .O(N__46375),
            .I(n12091));
    InMux I__10099 (
            .O(N__46372),
            .I(N__46369));
    LocalMux I__10098 (
            .O(N__46369),
            .I(N__46366));
    Odrv12 I__10097 (
            .O(N__46366),
            .I(n5_adj_565));
    InMux I__10096 (
            .O(N__46363),
            .I(n12092));
    InMux I__10095 (
            .O(N__46360),
            .I(N__46357));
    LocalMux I__10094 (
            .O(N__46357),
            .I(N__46354));
    Span4Mux_v I__10093 (
            .O(N__46354),
            .I(N__46351));
    Odrv4 I__10092 (
            .O(N__46351),
            .I(n4_adj_566));
    InMux I__10091 (
            .O(N__46348),
            .I(N__46344));
    InMux I__10090 (
            .O(N__46347),
            .I(N__46341));
    LocalMux I__10089 (
            .O(N__46344),
            .I(N__46338));
    LocalMux I__10088 (
            .O(N__46341),
            .I(N__46335));
    Span4Mux_h I__10087 (
            .O(N__46338),
            .I(N__46332));
    Span4Mux_h I__10086 (
            .O(N__46335),
            .I(N__46329));
    Odrv4 I__10085 (
            .O(N__46332),
            .I(duty_21));
    Odrv4 I__10084 (
            .O(N__46329),
            .I(duty_21));
    InMux I__10083 (
            .O(N__46324),
            .I(n12093));
    InMux I__10082 (
            .O(N__46321),
            .I(N__46318));
    LocalMux I__10081 (
            .O(N__46318),
            .I(N__46315));
    Span4Mux_h I__10080 (
            .O(N__46315),
            .I(N__46311));
    InMux I__10079 (
            .O(N__46314),
            .I(N__46308));
    Odrv4 I__10078 (
            .O(N__46311),
            .I(duty_6));
    LocalMux I__10077 (
            .O(N__46308),
            .I(duty_6));
    InMux I__10076 (
            .O(N__46303),
            .I(n12078));
    CascadeMux I__10075 (
            .O(N__46300),
            .I(N__46297));
    InMux I__10074 (
            .O(N__46297),
            .I(N__46294));
    LocalMux I__10073 (
            .O(N__46294),
            .I(N__46291));
    Odrv12 I__10072 (
            .O(N__46291),
            .I(n18_adj_552));
    InMux I__10071 (
            .O(N__46288),
            .I(n12079));
    CascadeMux I__10070 (
            .O(N__46285),
            .I(N__46282));
    InMux I__10069 (
            .O(N__46282),
            .I(N__46279));
    LocalMux I__10068 (
            .O(N__46279),
            .I(N__46276));
    Span4Mux_h I__10067 (
            .O(N__46276),
            .I(N__46273));
    Odrv4 I__10066 (
            .O(N__46273),
            .I(n17_adj_553));
    InMux I__10065 (
            .O(N__46270),
            .I(bfn_14_27_0_));
    CascadeMux I__10064 (
            .O(N__46267),
            .I(N__46264));
    InMux I__10063 (
            .O(N__46264),
            .I(N__46261));
    LocalMux I__10062 (
            .O(N__46261),
            .I(N__46258));
    Span4Mux_h I__10061 (
            .O(N__46258),
            .I(N__46255));
    Odrv4 I__10060 (
            .O(N__46255),
            .I(n16_adj_554));
    InMux I__10059 (
            .O(N__46252),
            .I(n12081));
    CascadeMux I__10058 (
            .O(N__46249),
            .I(N__46246));
    InMux I__10057 (
            .O(N__46246),
            .I(N__46243));
    LocalMux I__10056 (
            .O(N__46243),
            .I(N__46240));
    Span4Mux_h I__10055 (
            .O(N__46240),
            .I(N__46237));
    Odrv4 I__10054 (
            .O(N__46237),
            .I(n15_adj_555));
    InMux I__10053 (
            .O(N__46234),
            .I(N__46231));
    LocalMux I__10052 (
            .O(N__46231),
            .I(N__46228));
    Span4Mux_v I__10051 (
            .O(N__46228),
            .I(N__46224));
    InMux I__10050 (
            .O(N__46227),
            .I(N__46221));
    Odrv4 I__10049 (
            .O(N__46224),
            .I(duty_10));
    LocalMux I__10048 (
            .O(N__46221),
            .I(duty_10));
    InMux I__10047 (
            .O(N__46216),
            .I(n12082));
    CascadeMux I__10046 (
            .O(N__46213),
            .I(N__46210));
    InMux I__10045 (
            .O(N__46210),
            .I(N__46207));
    LocalMux I__10044 (
            .O(N__46207),
            .I(N__46204));
    Span4Mux_v I__10043 (
            .O(N__46204),
            .I(N__46201));
    Odrv4 I__10042 (
            .O(N__46201),
            .I(n14_adj_556));
    InMux I__10041 (
            .O(N__46198),
            .I(N__46194));
    InMux I__10040 (
            .O(N__46197),
            .I(N__46191));
    LocalMux I__10039 (
            .O(N__46194),
            .I(N__46188));
    LocalMux I__10038 (
            .O(N__46191),
            .I(N__46185));
    Span4Mux_v I__10037 (
            .O(N__46188),
            .I(N__46182));
    Span4Mux_h I__10036 (
            .O(N__46185),
            .I(N__46179));
    Odrv4 I__10035 (
            .O(N__46182),
            .I(duty_11));
    Odrv4 I__10034 (
            .O(N__46179),
            .I(duty_11));
    InMux I__10033 (
            .O(N__46174),
            .I(n12083));
    InMux I__10032 (
            .O(N__46171),
            .I(N__46168));
    LocalMux I__10031 (
            .O(N__46168),
            .I(N__46165));
    Span4Mux_h I__10030 (
            .O(N__46165),
            .I(N__46162));
    Odrv4 I__10029 (
            .O(N__46162),
            .I(n13_adj_557));
    InMux I__10028 (
            .O(N__46159),
            .I(n12084));
    CascadeMux I__10027 (
            .O(N__46156),
            .I(N__46153));
    InMux I__10026 (
            .O(N__46153),
            .I(N__46150));
    LocalMux I__10025 (
            .O(N__46150),
            .I(N__46147));
    Odrv12 I__10024 (
            .O(N__46147),
            .I(n12_adj_558));
    InMux I__10023 (
            .O(N__46144),
            .I(n12085));
    CascadeMux I__10022 (
            .O(N__46141),
            .I(N__46138));
    InMux I__10021 (
            .O(N__46138),
            .I(N__46135));
    LocalMux I__10020 (
            .O(N__46135),
            .I(N__46130));
    InMux I__10019 (
            .O(N__46134),
            .I(N__46127));
    InMux I__10018 (
            .O(N__46133),
            .I(N__46124));
    Span4Mux_h I__10017 (
            .O(N__46130),
            .I(N__46121));
    LocalMux I__10016 (
            .O(N__46127),
            .I(n3223));
    LocalMux I__10015 (
            .O(N__46124),
            .I(n3223));
    Odrv4 I__10014 (
            .O(N__46121),
            .I(n3223));
    InMux I__10013 (
            .O(N__46114),
            .I(N__46111));
    LocalMux I__10012 (
            .O(N__46111),
            .I(n14366));
    InMux I__10011 (
            .O(N__46108),
            .I(N__46103));
    InMux I__10010 (
            .O(N__46107),
            .I(N__46100));
    InMux I__10009 (
            .O(N__46106),
            .I(N__46097));
    LocalMux I__10008 (
            .O(N__46103),
            .I(n3227));
    LocalMux I__10007 (
            .O(N__46100),
            .I(n3227));
    LocalMux I__10006 (
            .O(N__46097),
            .I(n3227));
    CascadeMux I__10005 (
            .O(N__46090),
            .I(N__46087));
    InMux I__10004 (
            .O(N__46087),
            .I(N__46084));
    LocalMux I__10003 (
            .O(N__46084),
            .I(N__46081));
    Odrv12 I__10002 (
            .O(N__46081),
            .I(n25_adj_545));
    InMux I__10001 (
            .O(N__46078),
            .I(bfn_14_26_0_));
    CascadeMux I__10000 (
            .O(N__46075),
            .I(N__46072));
    InMux I__9999 (
            .O(N__46072),
            .I(N__46069));
    LocalMux I__9998 (
            .O(N__46069),
            .I(N__46066));
    Odrv12 I__9997 (
            .O(N__46066),
            .I(n24_adj_546));
    InMux I__9996 (
            .O(N__46063),
            .I(n12073));
    InMux I__9995 (
            .O(N__46060),
            .I(N__46057));
    LocalMux I__9994 (
            .O(N__46057),
            .I(N__46054));
    Span4Mux_h I__9993 (
            .O(N__46054),
            .I(N__46051));
    Odrv4 I__9992 (
            .O(N__46051),
            .I(n23_adj_547));
    InMux I__9991 (
            .O(N__46048),
            .I(N__46045));
    LocalMux I__9990 (
            .O(N__46045),
            .I(N__46042));
    Span4Mux_v I__9989 (
            .O(N__46042),
            .I(N__46038));
    InMux I__9988 (
            .O(N__46041),
            .I(N__46035));
    Odrv4 I__9987 (
            .O(N__46038),
            .I(duty_2));
    LocalMux I__9986 (
            .O(N__46035),
            .I(duty_2));
    InMux I__9985 (
            .O(N__46030),
            .I(n12074));
    CascadeMux I__9984 (
            .O(N__46027),
            .I(N__46024));
    InMux I__9983 (
            .O(N__46024),
            .I(N__46021));
    LocalMux I__9982 (
            .O(N__46021),
            .I(n22_adj_548));
    InMux I__9981 (
            .O(N__46018),
            .I(n12075));
    CascadeMux I__9980 (
            .O(N__46015),
            .I(N__46012));
    InMux I__9979 (
            .O(N__46012),
            .I(N__46009));
    LocalMux I__9978 (
            .O(N__46009),
            .I(N__46006));
    Odrv12 I__9977 (
            .O(N__46006),
            .I(n21_adj_549));
    InMux I__9976 (
            .O(N__46003),
            .I(N__45999));
    InMux I__9975 (
            .O(N__46002),
            .I(N__45996));
    LocalMux I__9974 (
            .O(N__45999),
            .I(N__45993));
    LocalMux I__9973 (
            .O(N__45996),
            .I(N__45990));
    Span4Mux_h I__9972 (
            .O(N__45993),
            .I(N__45987));
    Span4Mux_h I__9971 (
            .O(N__45990),
            .I(N__45984));
    Odrv4 I__9970 (
            .O(N__45987),
            .I(duty_4));
    Odrv4 I__9969 (
            .O(N__45984),
            .I(duty_4));
    InMux I__9968 (
            .O(N__45979),
            .I(n12076));
    CascadeMux I__9967 (
            .O(N__45976),
            .I(N__45973));
    InMux I__9966 (
            .O(N__45973),
            .I(N__45970));
    LocalMux I__9965 (
            .O(N__45970),
            .I(N__45967));
    Span4Mux_v I__9964 (
            .O(N__45967),
            .I(N__45964));
    Odrv4 I__9963 (
            .O(N__45964),
            .I(n20_adj_550));
    InMux I__9962 (
            .O(N__45961),
            .I(N__45958));
    LocalMux I__9961 (
            .O(N__45958),
            .I(N__45955));
    Span4Mux_h I__9960 (
            .O(N__45955),
            .I(N__45951));
    InMux I__9959 (
            .O(N__45954),
            .I(N__45948));
    Odrv4 I__9958 (
            .O(N__45951),
            .I(duty_5));
    LocalMux I__9957 (
            .O(N__45948),
            .I(duty_5));
    InMux I__9956 (
            .O(N__45943),
            .I(n12077));
    CascadeMux I__9955 (
            .O(N__45940),
            .I(N__45936));
    InMux I__9954 (
            .O(N__45939),
            .I(N__45933));
    InMux I__9953 (
            .O(N__45936),
            .I(N__45930));
    LocalMux I__9952 (
            .O(N__45933),
            .I(N__45927));
    LocalMux I__9951 (
            .O(N__45930),
            .I(N__45924));
    Span4Mux_h I__9950 (
            .O(N__45927),
            .I(N__45919));
    Span4Mux_v I__9949 (
            .O(N__45924),
            .I(N__45919));
    Odrv4 I__9948 (
            .O(N__45919),
            .I(n3006));
    CascadeMux I__9947 (
            .O(N__45916),
            .I(N__45912));
    InMux I__9946 (
            .O(N__45915),
            .I(N__45909));
    InMux I__9945 (
            .O(N__45912),
            .I(N__45906));
    LocalMux I__9944 (
            .O(N__45909),
            .I(N__45903));
    LocalMux I__9943 (
            .O(N__45906),
            .I(N__45900));
    Span4Mux_h I__9942 (
            .O(N__45903),
            .I(N__45897));
    Span4Mux_h I__9941 (
            .O(N__45900),
            .I(N__45894));
    Odrv4 I__9940 (
            .O(N__45897),
            .I(n15123));
    Odrv4 I__9939 (
            .O(N__45894),
            .I(n15123));
    InMux I__9938 (
            .O(N__45889),
            .I(n12491));
    InMux I__9937 (
            .O(N__45886),
            .I(N__45883));
    LocalMux I__9936 (
            .O(N__45883),
            .I(n3295));
    CascadeMux I__9935 (
            .O(N__45880),
            .I(N__45877));
    InMux I__9934 (
            .O(N__45877),
            .I(N__45874));
    LocalMux I__9933 (
            .O(N__45874),
            .I(n3294));
    InMux I__9932 (
            .O(N__45871),
            .I(N__45867));
    InMux I__9931 (
            .O(N__45870),
            .I(N__45864));
    LocalMux I__9930 (
            .O(N__45867),
            .I(N__45860));
    LocalMux I__9929 (
            .O(N__45864),
            .I(N__45857));
    InMux I__9928 (
            .O(N__45863),
            .I(N__45854));
    Span4Mux_v I__9927 (
            .O(N__45860),
            .I(N__45851));
    Span4Mux_v I__9926 (
            .O(N__45857),
            .I(N__45848));
    LocalMux I__9925 (
            .O(N__45854),
            .I(N__45845));
    Odrv4 I__9924 (
            .O(N__45851),
            .I(n3221));
    Odrv4 I__9923 (
            .O(N__45848),
            .I(n3221));
    Odrv12 I__9922 (
            .O(N__45845),
            .I(n3221));
    CascadeMux I__9921 (
            .O(N__45838),
            .I(N__45834));
    InMux I__9920 (
            .O(N__45837),
            .I(N__45830));
    InMux I__9919 (
            .O(N__45834),
            .I(N__45827));
    InMux I__9918 (
            .O(N__45833),
            .I(N__45824));
    LocalMux I__9917 (
            .O(N__45830),
            .I(N__45821));
    LocalMux I__9916 (
            .O(N__45827),
            .I(N__45816));
    LocalMux I__9915 (
            .O(N__45824),
            .I(N__45816));
    Span4Mux_v I__9914 (
            .O(N__45821),
            .I(N__45813));
    Span4Mux_v I__9913 (
            .O(N__45816),
            .I(N__45810));
    Odrv4 I__9912 (
            .O(N__45813),
            .I(n3218));
    Odrv4 I__9911 (
            .O(N__45810),
            .I(n3218));
    CascadeMux I__9910 (
            .O(N__45805),
            .I(n14368_cascade_));
    CascadeMux I__9909 (
            .O(N__45802),
            .I(N__45799));
    InMux I__9908 (
            .O(N__45799),
            .I(N__45796));
    LocalMux I__9907 (
            .O(N__45796),
            .I(N__45793));
    Span4Mux_v I__9906 (
            .O(N__45793),
            .I(N__45790));
    Odrv4 I__9905 (
            .O(N__45790),
            .I(n14374));
    CascadeMux I__9904 (
            .O(N__45787),
            .I(N__45784));
    InMux I__9903 (
            .O(N__45784),
            .I(N__45780));
    InMux I__9902 (
            .O(N__45783),
            .I(N__45777));
    LocalMux I__9901 (
            .O(N__45780),
            .I(N__45774));
    LocalMux I__9900 (
            .O(N__45777),
            .I(n3228));
    Odrv4 I__9899 (
            .O(N__45774),
            .I(n3228));
    CascadeMux I__9898 (
            .O(N__45769),
            .I(n3228_cascade_));
    InMux I__9897 (
            .O(N__45766),
            .I(N__45762));
    InMux I__9896 (
            .O(N__45765),
            .I(N__45759));
    LocalMux I__9895 (
            .O(N__45762),
            .I(N__45753));
    LocalMux I__9894 (
            .O(N__45759),
            .I(N__45753));
    InMux I__9893 (
            .O(N__45758),
            .I(N__45750));
    Odrv4 I__9892 (
            .O(N__45753),
            .I(n3224));
    LocalMux I__9891 (
            .O(N__45750),
            .I(n3224));
    CascadeMux I__9890 (
            .O(N__45745),
            .I(N__45742));
    InMux I__9889 (
            .O(N__45742),
            .I(N__45739));
    LocalMux I__9888 (
            .O(N__45739),
            .I(n14362));
    CascadeMux I__9887 (
            .O(N__45736),
            .I(N__45733));
    InMux I__9886 (
            .O(N__45733),
            .I(N__45729));
    InMux I__9885 (
            .O(N__45732),
            .I(N__45726));
    LocalMux I__9884 (
            .O(N__45729),
            .I(n3014));
    LocalMux I__9883 (
            .O(N__45726),
            .I(n3014));
    InMux I__9882 (
            .O(N__45721),
            .I(N__45718));
    LocalMux I__9881 (
            .O(N__45718),
            .I(N__45715));
    Odrv4 I__9880 (
            .O(N__45715),
            .I(n3081));
    InMux I__9879 (
            .O(N__45712),
            .I(n12483));
    InMux I__9878 (
            .O(N__45709),
            .I(N__45706));
    LocalMux I__9877 (
            .O(N__45706),
            .I(N__45701));
    InMux I__9876 (
            .O(N__45705),
            .I(N__45698));
    InMux I__9875 (
            .O(N__45704),
            .I(N__45695));
    Span4Mux_h I__9874 (
            .O(N__45701),
            .I(N__45692));
    LocalMux I__9873 (
            .O(N__45698),
            .I(N__45689));
    LocalMux I__9872 (
            .O(N__45695),
            .I(n3013));
    Odrv4 I__9871 (
            .O(N__45692),
            .I(n3013));
    Odrv4 I__9870 (
            .O(N__45689),
            .I(n3013));
    InMux I__9869 (
            .O(N__45682),
            .I(N__45679));
    LocalMux I__9868 (
            .O(N__45679),
            .I(N__45676));
    Odrv4 I__9867 (
            .O(N__45676),
            .I(n3080));
    InMux I__9866 (
            .O(N__45673),
            .I(n12484));
    InMux I__9865 (
            .O(N__45670),
            .I(N__45665));
    InMux I__9864 (
            .O(N__45669),
            .I(N__45662));
    CascadeMux I__9863 (
            .O(N__45668),
            .I(N__45659));
    LocalMux I__9862 (
            .O(N__45665),
            .I(N__45654));
    LocalMux I__9861 (
            .O(N__45662),
            .I(N__45654));
    InMux I__9860 (
            .O(N__45659),
            .I(N__45651));
    Odrv4 I__9859 (
            .O(N__45654),
            .I(n3012));
    LocalMux I__9858 (
            .O(N__45651),
            .I(n3012));
    InMux I__9857 (
            .O(N__45646),
            .I(N__45643));
    LocalMux I__9856 (
            .O(N__45643),
            .I(N__45640));
    Odrv12 I__9855 (
            .O(N__45640),
            .I(n3079));
    InMux I__9854 (
            .O(N__45637),
            .I(n12485));
    InMux I__9853 (
            .O(N__45634),
            .I(n12486));
    CascadeMux I__9852 (
            .O(N__45631),
            .I(N__45628));
    InMux I__9851 (
            .O(N__45628),
            .I(N__45625));
    LocalMux I__9850 (
            .O(N__45625),
            .I(N__45622));
    Span4Mux_v I__9849 (
            .O(N__45622),
            .I(N__45618));
    InMux I__9848 (
            .O(N__45621),
            .I(N__45615));
    Odrv4 I__9847 (
            .O(N__45618),
            .I(n3010));
    LocalMux I__9846 (
            .O(N__45615),
            .I(n3010));
    InMux I__9845 (
            .O(N__45610),
            .I(N__45607));
    LocalMux I__9844 (
            .O(N__45607),
            .I(N__45604));
    Span4Mux_v I__9843 (
            .O(N__45604),
            .I(N__45601));
    Span4Mux_h I__9842 (
            .O(N__45601),
            .I(N__45598));
    Odrv4 I__9841 (
            .O(N__45598),
            .I(n3077));
    InMux I__9840 (
            .O(N__45595),
            .I(bfn_14_24_0_));
    InMux I__9839 (
            .O(N__45592),
            .I(n12488));
    InMux I__9838 (
            .O(N__45589),
            .I(N__45585));
    InMux I__9837 (
            .O(N__45588),
            .I(N__45582));
    LocalMux I__9836 (
            .O(N__45585),
            .I(N__45579));
    LocalMux I__9835 (
            .O(N__45582),
            .I(N__45575));
    Span4Mux_v I__9834 (
            .O(N__45579),
            .I(N__45572));
    InMux I__9833 (
            .O(N__45578),
            .I(N__45569));
    Odrv4 I__9832 (
            .O(N__45575),
            .I(n3008));
    Odrv4 I__9831 (
            .O(N__45572),
            .I(n3008));
    LocalMux I__9830 (
            .O(N__45569),
            .I(n3008));
    CascadeMux I__9829 (
            .O(N__45562),
            .I(N__45559));
    InMux I__9828 (
            .O(N__45559),
            .I(N__45556));
    LocalMux I__9827 (
            .O(N__45556),
            .I(N__45553));
    Span4Mux_h I__9826 (
            .O(N__45553),
            .I(N__45550));
    Odrv4 I__9825 (
            .O(N__45550),
            .I(n3075));
    InMux I__9824 (
            .O(N__45547),
            .I(n12489));
    InMux I__9823 (
            .O(N__45544),
            .I(N__45540));
    InMux I__9822 (
            .O(N__45543),
            .I(N__45537));
    LocalMux I__9821 (
            .O(N__45540),
            .I(N__45534));
    LocalMux I__9820 (
            .O(N__45537),
            .I(N__45530));
    Span4Mux_h I__9819 (
            .O(N__45534),
            .I(N__45527));
    InMux I__9818 (
            .O(N__45533),
            .I(N__45524));
    Odrv4 I__9817 (
            .O(N__45530),
            .I(n3007));
    Odrv4 I__9816 (
            .O(N__45527),
            .I(n3007));
    LocalMux I__9815 (
            .O(N__45524),
            .I(n3007));
    CascadeMux I__9814 (
            .O(N__45517),
            .I(N__45514));
    InMux I__9813 (
            .O(N__45514),
            .I(N__45511));
    LocalMux I__9812 (
            .O(N__45511),
            .I(N__45508));
    Span4Mux_v I__9811 (
            .O(N__45508),
            .I(N__45505));
    Span4Mux_h I__9810 (
            .O(N__45505),
            .I(N__45502));
    Odrv4 I__9809 (
            .O(N__45502),
            .I(n3074));
    InMux I__9808 (
            .O(N__45499),
            .I(n12490));
    CascadeMux I__9807 (
            .O(N__45496),
            .I(N__45492));
    InMux I__9806 (
            .O(N__45495),
            .I(N__45488));
    InMux I__9805 (
            .O(N__45492),
            .I(N__45485));
    InMux I__9804 (
            .O(N__45491),
            .I(N__45482));
    LocalMux I__9803 (
            .O(N__45488),
            .I(n3022));
    LocalMux I__9802 (
            .O(N__45485),
            .I(n3022));
    LocalMux I__9801 (
            .O(N__45482),
            .I(n3022));
    CascadeMux I__9800 (
            .O(N__45475),
            .I(N__45472));
    InMux I__9799 (
            .O(N__45472),
            .I(N__45469));
    LocalMux I__9798 (
            .O(N__45469),
            .I(N__45466));
    Span4Mux_v I__9797 (
            .O(N__45466),
            .I(N__45463));
    Odrv4 I__9796 (
            .O(N__45463),
            .I(n3089));
    InMux I__9795 (
            .O(N__45460),
            .I(n12475));
    CascadeMux I__9794 (
            .O(N__45457),
            .I(N__45453));
    CascadeMux I__9793 (
            .O(N__45456),
            .I(N__45450));
    InMux I__9792 (
            .O(N__45453),
            .I(N__45447));
    InMux I__9791 (
            .O(N__45450),
            .I(N__45444));
    LocalMux I__9790 (
            .O(N__45447),
            .I(n3021));
    LocalMux I__9789 (
            .O(N__45444),
            .I(n3021));
    InMux I__9788 (
            .O(N__45439),
            .I(N__45436));
    LocalMux I__9787 (
            .O(N__45436),
            .I(n3088));
    InMux I__9786 (
            .O(N__45433),
            .I(n12476));
    CascadeMux I__9785 (
            .O(N__45430),
            .I(N__45427));
    InMux I__9784 (
            .O(N__45427),
            .I(N__45424));
    LocalMux I__9783 (
            .O(N__45424),
            .I(N__45419));
    InMux I__9782 (
            .O(N__45423),
            .I(N__45416));
    InMux I__9781 (
            .O(N__45422),
            .I(N__45413));
    Span4Mux_v I__9780 (
            .O(N__45419),
            .I(N__45408));
    LocalMux I__9779 (
            .O(N__45416),
            .I(N__45408));
    LocalMux I__9778 (
            .O(N__45413),
            .I(n3020));
    Odrv4 I__9777 (
            .O(N__45408),
            .I(n3020));
    CascadeMux I__9776 (
            .O(N__45403),
            .I(N__45400));
    InMux I__9775 (
            .O(N__45400),
            .I(N__45397));
    LocalMux I__9774 (
            .O(N__45397),
            .I(N__45394));
    Span4Mux_v I__9773 (
            .O(N__45394),
            .I(N__45391));
    Span4Mux_h I__9772 (
            .O(N__45391),
            .I(N__45388));
    Odrv4 I__9771 (
            .O(N__45388),
            .I(n3087));
    InMux I__9770 (
            .O(N__45385),
            .I(n12477));
    InMux I__9769 (
            .O(N__45382),
            .I(N__45379));
    LocalMux I__9768 (
            .O(N__45379),
            .I(N__45375));
    InMux I__9767 (
            .O(N__45378),
            .I(N__45372));
    Span4Mux_v I__9766 (
            .O(N__45375),
            .I(N__45367));
    LocalMux I__9765 (
            .O(N__45372),
            .I(N__45367));
    Odrv4 I__9764 (
            .O(N__45367),
            .I(n3019));
    InMux I__9763 (
            .O(N__45364),
            .I(N__45361));
    LocalMux I__9762 (
            .O(N__45361),
            .I(N__45358));
    Span4Mux_v I__9761 (
            .O(N__45358),
            .I(N__45355));
    Odrv4 I__9760 (
            .O(N__45355),
            .I(n3086));
    InMux I__9759 (
            .O(N__45352),
            .I(n12478));
    CascadeMux I__9758 (
            .O(N__45349),
            .I(N__45346));
    InMux I__9757 (
            .O(N__45346),
            .I(N__45342));
    InMux I__9756 (
            .O(N__45345),
            .I(N__45339));
    LocalMux I__9755 (
            .O(N__45342),
            .I(N__45333));
    LocalMux I__9754 (
            .O(N__45339),
            .I(N__45333));
    InMux I__9753 (
            .O(N__45338),
            .I(N__45330));
    Span4Mux_v I__9752 (
            .O(N__45333),
            .I(N__45327));
    LocalMux I__9751 (
            .O(N__45330),
            .I(n3018));
    Odrv4 I__9750 (
            .O(N__45327),
            .I(n3018));
    InMux I__9749 (
            .O(N__45322),
            .I(N__45319));
    LocalMux I__9748 (
            .O(N__45319),
            .I(N__45316));
    Span4Mux_h I__9747 (
            .O(N__45316),
            .I(N__45313));
    Odrv4 I__9746 (
            .O(N__45313),
            .I(n3085));
    InMux I__9745 (
            .O(N__45310),
            .I(bfn_14_23_0_));
    InMux I__9744 (
            .O(N__45307),
            .I(N__45304));
    LocalMux I__9743 (
            .O(N__45304),
            .I(N__45300));
    InMux I__9742 (
            .O(N__45303),
            .I(N__45297));
    Span4Mux_h I__9741 (
            .O(N__45300),
            .I(N__45292));
    LocalMux I__9740 (
            .O(N__45297),
            .I(N__45292));
    Odrv4 I__9739 (
            .O(N__45292),
            .I(n3017));
    InMux I__9738 (
            .O(N__45289),
            .I(N__45286));
    LocalMux I__9737 (
            .O(N__45286),
            .I(N__45283));
    Span4Mux_h I__9736 (
            .O(N__45283),
            .I(N__45280));
    Odrv4 I__9735 (
            .O(N__45280),
            .I(n3084));
    InMux I__9734 (
            .O(N__45277),
            .I(n12480));
    InMux I__9733 (
            .O(N__45274),
            .I(N__45270));
    CascadeMux I__9732 (
            .O(N__45273),
            .I(N__45266));
    LocalMux I__9731 (
            .O(N__45270),
            .I(N__45263));
    InMux I__9730 (
            .O(N__45269),
            .I(N__45260));
    InMux I__9729 (
            .O(N__45266),
            .I(N__45257));
    Span4Mux_v I__9728 (
            .O(N__45263),
            .I(N__45252));
    LocalMux I__9727 (
            .O(N__45260),
            .I(N__45252));
    LocalMux I__9726 (
            .O(N__45257),
            .I(n3016));
    Odrv4 I__9725 (
            .O(N__45252),
            .I(n3016));
    InMux I__9724 (
            .O(N__45247),
            .I(N__45244));
    LocalMux I__9723 (
            .O(N__45244),
            .I(N__45241));
    Span4Mux_v I__9722 (
            .O(N__45241),
            .I(N__45238));
    Odrv4 I__9721 (
            .O(N__45238),
            .I(n3083));
    InMux I__9720 (
            .O(N__45235),
            .I(n12481));
    InMux I__9719 (
            .O(N__45232),
            .I(n12482));
    CascadeMux I__9718 (
            .O(N__45229),
            .I(N__45226));
    InMux I__9717 (
            .O(N__45226),
            .I(N__45222));
    InMux I__9716 (
            .O(N__45225),
            .I(N__45218));
    LocalMux I__9715 (
            .O(N__45222),
            .I(N__45215));
    InMux I__9714 (
            .O(N__45221),
            .I(N__45212));
    LocalMux I__9713 (
            .O(N__45218),
            .I(n3030));
    Odrv4 I__9712 (
            .O(N__45215),
            .I(n3030));
    LocalMux I__9711 (
            .O(N__45212),
            .I(n3030));
    CascadeMux I__9710 (
            .O(N__45205),
            .I(N__45202));
    InMux I__9709 (
            .O(N__45202),
            .I(N__45199));
    LocalMux I__9708 (
            .O(N__45199),
            .I(N__45196));
    Span4Mux_v I__9707 (
            .O(N__45196),
            .I(N__45193));
    Odrv4 I__9706 (
            .O(N__45193),
            .I(n3097));
    InMux I__9705 (
            .O(N__45190),
            .I(n12467));
    InMux I__9704 (
            .O(N__45187),
            .I(N__45184));
    LocalMux I__9703 (
            .O(N__45184),
            .I(N__45181));
    Span4Mux_v I__9702 (
            .O(N__45181),
            .I(N__45177));
    InMux I__9701 (
            .O(N__45180),
            .I(N__45174));
    Odrv4 I__9700 (
            .O(N__45177),
            .I(n3029));
    LocalMux I__9699 (
            .O(N__45174),
            .I(n3029));
    InMux I__9698 (
            .O(N__45169),
            .I(N__45166));
    LocalMux I__9697 (
            .O(N__45166),
            .I(N__45163));
    Span4Mux_h I__9696 (
            .O(N__45163),
            .I(N__45160));
    Odrv4 I__9695 (
            .O(N__45160),
            .I(n3096));
    InMux I__9694 (
            .O(N__45157),
            .I(n12468));
    CascadeMux I__9693 (
            .O(N__45154),
            .I(N__45151));
    InMux I__9692 (
            .O(N__45151),
            .I(N__45147));
    InMux I__9691 (
            .O(N__45150),
            .I(N__45143));
    LocalMux I__9690 (
            .O(N__45147),
            .I(N__45140));
    InMux I__9689 (
            .O(N__45146),
            .I(N__45137));
    LocalMux I__9688 (
            .O(N__45143),
            .I(n3028));
    Odrv4 I__9687 (
            .O(N__45140),
            .I(n3028));
    LocalMux I__9686 (
            .O(N__45137),
            .I(n3028));
    InMux I__9685 (
            .O(N__45130),
            .I(N__45127));
    LocalMux I__9684 (
            .O(N__45127),
            .I(N__45124));
    Odrv12 I__9683 (
            .O(N__45124),
            .I(n3095));
    InMux I__9682 (
            .O(N__45121),
            .I(n12469));
    CascadeMux I__9681 (
            .O(N__45118),
            .I(N__45114));
    InMux I__9680 (
            .O(N__45117),
            .I(N__45110));
    InMux I__9679 (
            .O(N__45114),
            .I(N__45107));
    InMux I__9678 (
            .O(N__45113),
            .I(N__45104));
    LocalMux I__9677 (
            .O(N__45110),
            .I(n3027));
    LocalMux I__9676 (
            .O(N__45107),
            .I(n3027));
    LocalMux I__9675 (
            .O(N__45104),
            .I(n3027));
    InMux I__9674 (
            .O(N__45097),
            .I(N__45094));
    LocalMux I__9673 (
            .O(N__45094),
            .I(n3094));
    InMux I__9672 (
            .O(N__45091),
            .I(n12470));
    CascadeMux I__9671 (
            .O(N__45088),
            .I(N__45084));
    InMux I__9670 (
            .O(N__45087),
            .I(N__45080));
    InMux I__9669 (
            .O(N__45084),
            .I(N__45077));
    InMux I__9668 (
            .O(N__45083),
            .I(N__45074));
    LocalMux I__9667 (
            .O(N__45080),
            .I(n3026));
    LocalMux I__9666 (
            .O(N__45077),
            .I(n3026));
    LocalMux I__9665 (
            .O(N__45074),
            .I(n3026));
    InMux I__9664 (
            .O(N__45067),
            .I(N__45064));
    LocalMux I__9663 (
            .O(N__45064),
            .I(n3093));
    InMux I__9662 (
            .O(N__45061),
            .I(bfn_14_22_0_));
    CascadeMux I__9661 (
            .O(N__45058),
            .I(N__45055));
    InMux I__9660 (
            .O(N__45055),
            .I(N__45051));
    CascadeMux I__9659 (
            .O(N__45054),
            .I(N__45048));
    LocalMux I__9658 (
            .O(N__45051),
            .I(N__45045));
    InMux I__9657 (
            .O(N__45048),
            .I(N__45041));
    Span4Mux_h I__9656 (
            .O(N__45045),
            .I(N__45038));
    InMux I__9655 (
            .O(N__45044),
            .I(N__45035));
    LocalMux I__9654 (
            .O(N__45041),
            .I(n3025));
    Odrv4 I__9653 (
            .O(N__45038),
            .I(n3025));
    LocalMux I__9652 (
            .O(N__45035),
            .I(n3025));
    InMux I__9651 (
            .O(N__45028),
            .I(N__45025));
    LocalMux I__9650 (
            .O(N__45025),
            .I(N__45022));
    Span4Mux_v I__9649 (
            .O(N__45022),
            .I(N__45019));
    Odrv4 I__9648 (
            .O(N__45019),
            .I(n3092));
    InMux I__9647 (
            .O(N__45016),
            .I(n12472));
    CascadeMux I__9646 (
            .O(N__45013),
            .I(N__45009));
    InMux I__9645 (
            .O(N__45012),
            .I(N__45005));
    InMux I__9644 (
            .O(N__45009),
            .I(N__45002));
    InMux I__9643 (
            .O(N__45008),
            .I(N__44999));
    LocalMux I__9642 (
            .O(N__45005),
            .I(n3024));
    LocalMux I__9641 (
            .O(N__45002),
            .I(n3024));
    LocalMux I__9640 (
            .O(N__44999),
            .I(n3024));
    InMux I__9639 (
            .O(N__44992),
            .I(N__44989));
    LocalMux I__9638 (
            .O(N__44989),
            .I(N__44986));
    Odrv4 I__9637 (
            .O(N__44986),
            .I(n3091));
    InMux I__9636 (
            .O(N__44983),
            .I(n12473));
    CascadeMux I__9635 (
            .O(N__44980),
            .I(N__44976));
    InMux I__9634 (
            .O(N__44979),
            .I(N__44973));
    InMux I__9633 (
            .O(N__44976),
            .I(N__44970));
    LocalMux I__9632 (
            .O(N__44973),
            .I(n3023));
    LocalMux I__9631 (
            .O(N__44970),
            .I(n3023));
    CascadeMux I__9630 (
            .O(N__44965),
            .I(N__44962));
    InMux I__9629 (
            .O(N__44962),
            .I(N__44959));
    LocalMux I__9628 (
            .O(N__44959),
            .I(N__44956));
    Odrv4 I__9627 (
            .O(N__44956),
            .I(n3090));
    InMux I__9626 (
            .O(N__44953),
            .I(n12474));
    CascadeMux I__9625 (
            .O(N__44950),
            .I(N__44947));
    InMux I__9624 (
            .O(N__44947),
            .I(N__44944));
    LocalMux I__9623 (
            .O(N__44944),
            .I(N__44940));
    InMux I__9622 (
            .O(N__44943),
            .I(N__44936));
    Span4Mux_v I__9621 (
            .O(N__44940),
            .I(N__44933));
    InMux I__9620 (
            .O(N__44939),
            .I(N__44930));
    LocalMux I__9619 (
            .O(N__44936),
            .I(n2925));
    Odrv4 I__9618 (
            .O(N__44933),
            .I(n2925));
    LocalMux I__9617 (
            .O(N__44930),
            .I(n2925));
    CascadeMux I__9616 (
            .O(N__44923),
            .I(n3122_cascade_));
    InMux I__9615 (
            .O(N__44920),
            .I(N__44916));
    InMux I__9614 (
            .O(N__44919),
            .I(N__44913));
    LocalMux I__9613 (
            .O(N__44916),
            .I(N__44907));
    LocalMux I__9612 (
            .O(N__44913),
            .I(N__44907));
    InMux I__9611 (
            .O(N__44912),
            .I(N__44904));
    Span4Mux_v I__9610 (
            .O(N__44907),
            .I(N__44899));
    LocalMux I__9609 (
            .O(N__44904),
            .I(N__44899));
    Span4Mux_h I__9608 (
            .O(N__44899),
            .I(N__44896));
    Odrv4 I__9607 (
            .O(N__44896),
            .I(n2914));
    InMux I__9606 (
            .O(N__44893),
            .I(N__44889));
    InMux I__9605 (
            .O(N__44892),
            .I(N__44885));
    LocalMux I__9604 (
            .O(N__44889),
            .I(N__44882));
    InMux I__9603 (
            .O(N__44888),
            .I(N__44879));
    LocalMux I__9602 (
            .O(N__44885),
            .I(N__44876));
    Span4Mux_h I__9601 (
            .O(N__44882),
            .I(N__44873));
    LocalMux I__9600 (
            .O(N__44879),
            .I(N__44870));
    Span4Mux_h I__9599 (
            .O(N__44876),
            .I(N__44867));
    Span4Mux_h I__9598 (
            .O(N__44873),
            .I(N__44864));
    Span4Mux_h I__9597 (
            .O(N__44870),
            .I(N__44861));
    Odrv4 I__9596 (
            .O(N__44867),
            .I(n316));
    Odrv4 I__9595 (
            .O(N__44864),
            .I(n316));
    Odrv4 I__9594 (
            .O(N__44861),
            .I(n316));
    InMux I__9593 (
            .O(N__44854),
            .I(N__44851));
    LocalMux I__9592 (
            .O(N__44851),
            .I(N__44848));
    Span4Mux_h I__9591 (
            .O(N__44848),
            .I(N__44845));
    Span4Mux_h I__9590 (
            .O(N__44845),
            .I(N__44842));
    Odrv4 I__9589 (
            .O(N__44842),
            .I(n3101));
    InMux I__9588 (
            .O(N__44839),
            .I(bfn_14_21_0_));
    CascadeMux I__9587 (
            .O(N__44836),
            .I(N__44832));
    InMux I__9586 (
            .O(N__44835),
            .I(N__44829));
    InMux I__9585 (
            .O(N__44832),
            .I(N__44826));
    LocalMux I__9584 (
            .O(N__44829),
            .I(N__44823));
    LocalMux I__9583 (
            .O(N__44826),
            .I(N__44820));
    Span4Mux_h I__9582 (
            .O(N__44823),
            .I(N__44816));
    Span4Mux_h I__9581 (
            .O(N__44820),
            .I(N__44813));
    InMux I__9580 (
            .O(N__44819),
            .I(N__44810));
    Odrv4 I__9579 (
            .O(N__44816),
            .I(n3033));
    Odrv4 I__9578 (
            .O(N__44813),
            .I(n3033));
    LocalMux I__9577 (
            .O(N__44810),
            .I(n3033));
    InMux I__9576 (
            .O(N__44803),
            .I(N__44800));
    LocalMux I__9575 (
            .O(N__44800),
            .I(N__44797));
    Span12Mux_s11_v I__9574 (
            .O(N__44797),
            .I(N__44794));
    Odrv12 I__9573 (
            .O(N__44794),
            .I(n3100));
    InMux I__9572 (
            .O(N__44791),
            .I(n12464));
    InMux I__9571 (
            .O(N__44788),
            .I(N__44784));
    InMux I__9570 (
            .O(N__44787),
            .I(N__44781));
    LocalMux I__9569 (
            .O(N__44784),
            .I(N__44778));
    LocalMux I__9568 (
            .O(N__44781),
            .I(N__44775));
    Span4Mux_h I__9567 (
            .O(N__44778),
            .I(N__44772));
    Span4Mux_h I__9566 (
            .O(N__44775),
            .I(N__44769));
    Odrv4 I__9565 (
            .O(N__44772),
            .I(n3032));
    Odrv4 I__9564 (
            .O(N__44769),
            .I(n3032));
    CascadeMux I__9563 (
            .O(N__44764),
            .I(N__44761));
    InMux I__9562 (
            .O(N__44761),
            .I(N__44758));
    LocalMux I__9561 (
            .O(N__44758),
            .I(N__44755));
    Span4Mux_h I__9560 (
            .O(N__44755),
            .I(N__44752));
    Span4Mux_h I__9559 (
            .O(N__44752),
            .I(N__44749));
    Odrv4 I__9558 (
            .O(N__44749),
            .I(n3099));
    InMux I__9557 (
            .O(N__44746),
            .I(n12465));
    CascadeMux I__9556 (
            .O(N__44743),
            .I(N__44739));
    InMux I__9555 (
            .O(N__44742),
            .I(N__44736));
    InMux I__9554 (
            .O(N__44739),
            .I(N__44733));
    LocalMux I__9553 (
            .O(N__44736),
            .I(N__44729));
    LocalMux I__9552 (
            .O(N__44733),
            .I(N__44726));
    InMux I__9551 (
            .O(N__44732),
            .I(N__44723));
    Odrv4 I__9550 (
            .O(N__44729),
            .I(n3031));
    Odrv4 I__9549 (
            .O(N__44726),
            .I(n3031));
    LocalMux I__9548 (
            .O(N__44723),
            .I(n3031));
    InMux I__9547 (
            .O(N__44716),
            .I(N__44713));
    LocalMux I__9546 (
            .O(N__44713),
            .I(n3098));
    InMux I__9545 (
            .O(N__44710),
            .I(n12466));
    CascadeMux I__9544 (
            .O(N__44707),
            .I(n13932_cascade_));
    InMux I__9543 (
            .O(N__44704),
            .I(N__44701));
    LocalMux I__9542 (
            .O(N__44701),
            .I(n13936));
    InMux I__9541 (
            .O(N__44698),
            .I(N__44694));
    InMux I__9540 (
            .O(N__44697),
            .I(N__44691));
    LocalMux I__9539 (
            .O(N__44694),
            .I(N__44688));
    LocalMux I__9538 (
            .O(N__44691),
            .I(N__44685));
    Span4Mux_v I__9537 (
            .O(N__44688),
            .I(N__44681));
    Span4Mux_h I__9536 (
            .O(N__44685),
            .I(N__44678));
    InMux I__9535 (
            .O(N__44684),
            .I(N__44675));
    Odrv4 I__9534 (
            .O(N__44681),
            .I(n2926));
    Odrv4 I__9533 (
            .O(N__44678),
            .I(n2926));
    LocalMux I__9532 (
            .O(N__44675),
            .I(n2926));
    CascadeMux I__9531 (
            .O(N__44668),
            .I(N__44664));
    CascadeMux I__9530 (
            .O(N__44667),
            .I(N__44661));
    InMux I__9529 (
            .O(N__44664),
            .I(N__44658));
    InMux I__9528 (
            .O(N__44661),
            .I(N__44655));
    LocalMux I__9527 (
            .O(N__44658),
            .I(N__44651));
    LocalMux I__9526 (
            .O(N__44655),
            .I(N__44648));
    CascadeMux I__9525 (
            .O(N__44654),
            .I(N__44645));
    Span4Mux_v I__9524 (
            .O(N__44651),
            .I(N__44642));
    Span4Mux_h I__9523 (
            .O(N__44648),
            .I(N__44639));
    InMux I__9522 (
            .O(N__44645),
            .I(N__44636));
    Odrv4 I__9521 (
            .O(N__44642),
            .I(n2920));
    Odrv4 I__9520 (
            .O(N__44639),
            .I(n2920));
    LocalMux I__9519 (
            .O(N__44636),
            .I(n2920));
    CascadeMux I__9518 (
            .O(N__44629),
            .I(N__44626));
    InMux I__9517 (
            .O(N__44626),
            .I(N__44622));
    InMux I__9516 (
            .O(N__44625),
            .I(N__44619));
    LocalMux I__9515 (
            .O(N__44622),
            .I(N__44616));
    LocalMux I__9514 (
            .O(N__44619),
            .I(N__44610));
    Span4Mux_h I__9513 (
            .O(N__44616),
            .I(N__44610));
    InMux I__9512 (
            .O(N__44615),
            .I(N__44607));
    Odrv4 I__9511 (
            .O(N__44610),
            .I(n2927));
    LocalMux I__9510 (
            .O(N__44607),
            .I(n2927));
    InMux I__9509 (
            .O(N__44602),
            .I(N__44598));
    InMux I__9508 (
            .O(N__44601),
            .I(N__44595));
    LocalMux I__9507 (
            .O(N__44598),
            .I(N__44592));
    LocalMux I__9506 (
            .O(N__44595),
            .I(N__44589));
    Span4Mux_v I__9505 (
            .O(N__44592),
            .I(N__44585));
    Span4Mux_h I__9504 (
            .O(N__44589),
            .I(N__44582));
    InMux I__9503 (
            .O(N__44588),
            .I(N__44579));
    Odrv4 I__9502 (
            .O(N__44585),
            .I(n2919));
    Odrv4 I__9501 (
            .O(N__44582),
            .I(n2919));
    LocalMux I__9500 (
            .O(N__44579),
            .I(n2919));
    CascadeMux I__9499 (
            .O(N__44572),
            .I(N__44568));
    InMux I__9498 (
            .O(N__44571),
            .I(N__44565));
    InMux I__9497 (
            .O(N__44568),
            .I(N__44562));
    LocalMux I__9496 (
            .O(N__44565),
            .I(N__44557));
    LocalMux I__9495 (
            .O(N__44562),
            .I(N__44557));
    Span4Mux_h I__9494 (
            .O(N__44557),
            .I(N__44553));
    InMux I__9493 (
            .O(N__44556),
            .I(N__44550));
    Odrv4 I__9492 (
            .O(N__44553),
            .I(n2928));
    LocalMux I__9491 (
            .O(N__44550),
            .I(n2928));
    CascadeMux I__9490 (
            .O(N__44545),
            .I(N__44541));
    CascadeMux I__9489 (
            .O(N__44544),
            .I(N__44538));
    InMux I__9488 (
            .O(N__44541),
            .I(N__44535));
    InMux I__9487 (
            .O(N__44538),
            .I(N__44532));
    LocalMux I__9486 (
            .O(N__44535),
            .I(N__44529));
    LocalMux I__9485 (
            .O(N__44532),
            .I(N__44523));
    Span4Mux_h I__9484 (
            .O(N__44529),
            .I(N__44523));
    InMux I__9483 (
            .O(N__44528),
            .I(N__44520));
    Odrv4 I__9482 (
            .O(N__44523),
            .I(n2922));
    LocalMux I__9481 (
            .O(N__44520),
            .I(n2922));
    InMux I__9480 (
            .O(N__44515),
            .I(N__44512));
    LocalMux I__9479 (
            .O(N__44512),
            .I(N__44509));
    Span4Mux_h I__9478 (
            .O(N__44509),
            .I(N__44506));
    Odrv4 I__9477 (
            .O(N__44506),
            .I(n2793));
    CascadeMux I__9476 (
            .O(N__44503),
            .I(N__44500));
    InMux I__9475 (
            .O(N__44500),
            .I(N__44496));
    CascadeMux I__9474 (
            .O(N__44499),
            .I(N__44493));
    LocalMux I__9473 (
            .O(N__44496),
            .I(N__44490));
    InMux I__9472 (
            .O(N__44493),
            .I(N__44487));
    Span4Mux_h I__9471 (
            .O(N__44490),
            .I(N__44483));
    LocalMux I__9470 (
            .O(N__44487),
            .I(N__44480));
    InMux I__9469 (
            .O(N__44486),
            .I(N__44477));
    Odrv4 I__9468 (
            .O(N__44483),
            .I(n2726));
    Odrv4 I__9467 (
            .O(N__44480),
            .I(n2726));
    LocalMux I__9466 (
            .O(N__44477),
            .I(n2726));
    CascadeMux I__9465 (
            .O(N__44470),
            .I(n2825_cascade_));
    CascadeMux I__9464 (
            .O(N__44467),
            .I(N__44464));
    InMux I__9463 (
            .O(N__44464),
            .I(N__44461));
    LocalMux I__9462 (
            .O(N__44461),
            .I(N__44457));
    InMux I__9461 (
            .O(N__44460),
            .I(N__44453));
    Span4Mux_v I__9460 (
            .O(N__44457),
            .I(N__44450));
    InMux I__9459 (
            .O(N__44456),
            .I(N__44447));
    LocalMux I__9458 (
            .O(N__44453),
            .I(n2924));
    Odrv4 I__9457 (
            .O(N__44450),
            .I(n2924));
    LocalMux I__9456 (
            .O(N__44447),
            .I(n2924));
    InMux I__9455 (
            .O(N__44440),
            .I(N__44437));
    LocalMux I__9454 (
            .O(N__44437),
            .I(N__44434));
    Odrv4 I__9453 (
            .O(N__44434),
            .I(n2796));
    InMux I__9452 (
            .O(N__44431),
            .I(N__44427));
    CascadeMux I__9451 (
            .O(N__44430),
            .I(N__44424));
    LocalMux I__9450 (
            .O(N__44427),
            .I(N__44420));
    InMux I__9449 (
            .O(N__44424),
            .I(N__44417));
    InMux I__9448 (
            .O(N__44423),
            .I(N__44414));
    Span4Mux_h I__9447 (
            .O(N__44420),
            .I(N__44409));
    LocalMux I__9446 (
            .O(N__44417),
            .I(N__44409));
    LocalMux I__9445 (
            .O(N__44414),
            .I(n2729));
    Odrv4 I__9444 (
            .O(N__44409),
            .I(n2729));
    InMux I__9443 (
            .O(N__44404),
            .I(N__44401));
    LocalMux I__9442 (
            .O(N__44401),
            .I(N__44398));
    Span4Mux_h I__9441 (
            .O(N__44398),
            .I(N__44395));
    Odrv4 I__9440 (
            .O(N__44395),
            .I(n2800));
    CascadeMux I__9439 (
            .O(N__44392),
            .I(N__44389));
    InMux I__9438 (
            .O(N__44389),
            .I(N__44386));
    LocalMux I__9437 (
            .O(N__44386),
            .I(N__44382));
    CascadeMux I__9436 (
            .O(N__44385),
            .I(N__44378));
    Span4Mux_v I__9435 (
            .O(N__44382),
            .I(N__44375));
    InMux I__9434 (
            .O(N__44381),
            .I(N__44372));
    InMux I__9433 (
            .O(N__44378),
            .I(N__44369));
    Odrv4 I__9432 (
            .O(N__44375),
            .I(n2733));
    LocalMux I__9431 (
            .O(N__44372),
            .I(n2733));
    LocalMux I__9430 (
            .O(N__44369),
            .I(n2733));
    InMux I__9429 (
            .O(N__44362),
            .I(N__44359));
    LocalMux I__9428 (
            .O(N__44359),
            .I(N__44356));
    Span4Mux_h I__9427 (
            .O(N__44356),
            .I(N__44353));
    Odrv4 I__9426 (
            .O(N__44353),
            .I(n2799));
    InMux I__9425 (
            .O(N__44350),
            .I(N__44347));
    LocalMux I__9424 (
            .O(N__44347),
            .I(N__44343));
    CascadeMux I__9423 (
            .O(N__44346),
            .I(N__44340));
    Span4Mux_h I__9422 (
            .O(N__44343),
            .I(N__44337));
    InMux I__9421 (
            .O(N__44340),
            .I(N__44334));
    Odrv4 I__9420 (
            .O(N__44337),
            .I(n2732));
    LocalMux I__9419 (
            .O(N__44334),
            .I(n2732));
    InMux I__9418 (
            .O(N__44329),
            .I(N__44326));
    LocalMux I__9417 (
            .O(N__44326),
            .I(n14246));
    CascadeMux I__9416 (
            .O(N__44323),
            .I(n14248_cascade_));
    CascadeMux I__9415 (
            .O(N__44320),
            .I(n14254_cascade_));
    InMux I__9414 (
            .O(N__44317),
            .I(N__44314));
    LocalMux I__9413 (
            .O(N__44314),
            .I(n14266));
    CascadeMux I__9412 (
            .O(N__44311),
            .I(n2841_cascade_));
    CascadeMux I__9411 (
            .O(N__44308),
            .I(N__44305));
    InMux I__9410 (
            .O(N__44305),
            .I(N__44301));
    CascadeMux I__9409 (
            .O(N__44304),
            .I(N__44298));
    LocalMux I__9408 (
            .O(N__44301),
            .I(N__44295));
    InMux I__9407 (
            .O(N__44298),
            .I(N__44292));
    Span4Mux_h I__9406 (
            .O(N__44295),
            .I(N__44287));
    LocalMux I__9405 (
            .O(N__44292),
            .I(N__44287));
    Span4Mux_v I__9404 (
            .O(N__44287),
            .I(N__44283));
    InMux I__9403 (
            .O(N__44286),
            .I(N__44280));
    Odrv4 I__9402 (
            .O(N__44283),
            .I(n2923));
    LocalMux I__9401 (
            .O(N__44280),
            .I(n2923));
    InMux I__9400 (
            .O(N__44275),
            .I(N__44271));
    InMux I__9399 (
            .O(N__44274),
            .I(N__44267));
    LocalMux I__9398 (
            .O(N__44271),
            .I(N__44264));
    InMux I__9397 (
            .O(N__44270),
            .I(N__44261));
    LocalMux I__9396 (
            .O(N__44267),
            .I(N__44256));
    Span4Mux_s1_v I__9395 (
            .O(N__44264),
            .I(N__44256));
    LocalMux I__9394 (
            .O(N__44261),
            .I(pwm_counter_17));
    Odrv4 I__9393 (
            .O(N__44256),
            .I(pwm_counter_17));
    InMux I__9392 (
            .O(N__44251),
            .I(N__44247));
    InMux I__9391 (
            .O(N__44250),
            .I(N__44243));
    LocalMux I__9390 (
            .O(N__44247),
            .I(N__44240));
    InMux I__9389 (
            .O(N__44246),
            .I(N__44237));
    LocalMux I__9388 (
            .O(N__44243),
            .I(N__44234));
    Span4Mux_h I__9387 (
            .O(N__44240),
            .I(N__44229));
    LocalMux I__9386 (
            .O(N__44237),
            .I(N__44229));
    Odrv4 I__9385 (
            .O(N__44234),
            .I(n2712));
    Odrv4 I__9384 (
            .O(N__44229),
            .I(n2712));
    CascadeMux I__9383 (
            .O(N__44224),
            .I(N__44221));
    InMux I__9382 (
            .O(N__44221),
            .I(N__44218));
    LocalMux I__9381 (
            .O(N__44218),
            .I(N__44215));
    Span4Mux_h I__9380 (
            .O(N__44215),
            .I(N__44212));
    Odrv4 I__9379 (
            .O(N__44212),
            .I(n2779));
    CascadeMux I__9378 (
            .O(N__44209),
            .I(n2811_cascade_));
    InMux I__9377 (
            .O(N__44206),
            .I(N__44203));
    LocalMux I__9376 (
            .O(N__44203),
            .I(N__44200));
    Odrv12 I__9375 (
            .O(N__44200),
            .I(n2794));
    CascadeMux I__9374 (
            .O(N__44197),
            .I(N__44194));
    InMux I__9373 (
            .O(N__44194),
            .I(N__44190));
    CascadeMux I__9372 (
            .O(N__44193),
            .I(N__44186));
    LocalMux I__9371 (
            .O(N__44190),
            .I(N__44183));
    InMux I__9370 (
            .O(N__44189),
            .I(N__44180));
    InMux I__9369 (
            .O(N__44186),
            .I(N__44177));
    Span4Mux_h I__9368 (
            .O(N__44183),
            .I(N__44170));
    LocalMux I__9367 (
            .O(N__44180),
            .I(N__44170));
    LocalMux I__9366 (
            .O(N__44177),
            .I(N__44170));
    Odrv4 I__9365 (
            .O(N__44170),
            .I(n2727));
    InMux I__9364 (
            .O(N__44167),
            .I(N__44162));
    InMux I__9363 (
            .O(N__44166),
            .I(N__44159));
    InMux I__9362 (
            .O(N__44165),
            .I(N__44156));
    LocalMux I__9361 (
            .O(N__44162),
            .I(N__44153));
    LocalMux I__9360 (
            .O(N__44159),
            .I(N__44148));
    LocalMux I__9359 (
            .O(N__44156),
            .I(N__44148));
    Odrv4 I__9358 (
            .O(N__44153),
            .I(n2716));
    Odrv12 I__9357 (
            .O(N__44148),
            .I(n2716));
    CascadeMux I__9356 (
            .O(N__44143),
            .I(N__44140));
    InMux I__9355 (
            .O(N__44140),
            .I(N__44137));
    LocalMux I__9354 (
            .O(N__44137),
            .I(N__44134));
    Span4Mux_v I__9353 (
            .O(N__44134),
            .I(N__44131));
    Odrv4 I__9352 (
            .O(N__44131),
            .I(n2783));
    InMux I__9351 (
            .O(N__44128),
            .I(N__44125));
    LocalMux I__9350 (
            .O(N__44125),
            .I(N__44122));
    Span4Mux_v I__9349 (
            .O(N__44122),
            .I(N__44119));
    Odrv4 I__9348 (
            .O(N__44119),
            .I(n2782));
    CascadeMux I__9347 (
            .O(N__44116),
            .I(N__44112));
    InMux I__9346 (
            .O(N__44115),
            .I(N__44108));
    InMux I__9345 (
            .O(N__44112),
            .I(N__44105));
    InMux I__9344 (
            .O(N__44111),
            .I(N__44102));
    LocalMux I__9343 (
            .O(N__44108),
            .I(N__44097));
    LocalMux I__9342 (
            .O(N__44105),
            .I(N__44097));
    LocalMux I__9341 (
            .O(N__44102),
            .I(N__44094));
    Span4Mux_h I__9340 (
            .O(N__44097),
            .I(N__44091));
    Odrv4 I__9339 (
            .O(N__44094),
            .I(n2715));
    Odrv4 I__9338 (
            .O(N__44091),
            .I(n2715));
    CascadeMux I__9337 (
            .O(N__44086),
            .I(n2814_cascade_));
    InMux I__9336 (
            .O(N__44083),
            .I(N__44080));
    LocalMux I__9335 (
            .O(N__44080),
            .I(n14260));
    InMux I__9334 (
            .O(N__44077),
            .I(N__44074));
    LocalMux I__9333 (
            .O(N__44074),
            .I(N__44071));
    Odrv4 I__9332 (
            .O(N__44071),
            .I(pwm_setpoint_23_N_171_15));
    InMux I__9331 (
            .O(N__44068),
            .I(N__44065));
    LocalMux I__9330 (
            .O(N__44065),
            .I(pwm_setpoint_23_N_171_18));
    InMux I__9329 (
            .O(N__44062),
            .I(N__44057));
    InMux I__9328 (
            .O(N__44061),
            .I(N__44054));
    InMux I__9327 (
            .O(N__44060),
            .I(N__44051));
    LocalMux I__9326 (
            .O(N__44057),
            .I(N__44046));
    LocalMux I__9325 (
            .O(N__44054),
            .I(N__44046));
    LocalMux I__9324 (
            .O(N__44051),
            .I(pwm_counter_23));
    Odrv4 I__9323 (
            .O(N__44046),
            .I(pwm_counter_23));
    InMux I__9322 (
            .O(N__44041),
            .I(N__44038));
    LocalMux I__9321 (
            .O(N__44038),
            .I(\PWM.n28 ));
    CascadeMux I__9320 (
            .O(N__44035),
            .I(N__44032));
    InMux I__9319 (
            .O(N__44032),
            .I(N__44027));
    InMux I__9318 (
            .O(N__44031),
            .I(N__44024));
    InMux I__9317 (
            .O(N__44030),
            .I(N__44021));
    LocalMux I__9316 (
            .O(N__44027),
            .I(N__44018));
    LocalMux I__9315 (
            .O(N__44024),
            .I(N__44015));
    LocalMux I__9314 (
            .O(N__44021),
            .I(N__44008));
    Span4Mux_h I__9313 (
            .O(N__44018),
            .I(N__44008));
    Span4Mux_s2_v I__9312 (
            .O(N__44015),
            .I(N__44008));
    Odrv4 I__9311 (
            .O(N__44008),
            .I(pwm_counter_15));
    InMux I__9310 (
            .O(N__44005),
            .I(N__44001));
    InMux I__9309 (
            .O(N__44004),
            .I(N__43997));
    LocalMux I__9308 (
            .O(N__44001),
            .I(N__43994));
    InMux I__9307 (
            .O(N__44000),
            .I(N__43991));
    LocalMux I__9306 (
            .O(N__43997),
            .I(N__43984));
    Span4Mux_v I__9305 (
            .O(N__43994),
            .I(N__43984));
    LocalMux I__9304 (
            .O(N__43991),
            .I(N__43984));
    Odrv4 I__9303 (
            .O(N__43984),
            .I(pwm_counter_18));
    InMux I__9302 (
            .O(N__43981),
            .I(N__43978));
    LocalMux I__9301 (
            .O(N__43978),
            .I(n37));
    InMux I__9300 (
            .O(N__43975),
            .I(N__43969));
    InMux I__9299 (
            .O(N__43974),
            .I(N__43969));
    LocalMux I__9298 (
            .O(N__43969),
            .I(pwm_setpoint_18));
    CascadeMux I__9297 (
            .O(N__43966),
            .I(n37_cascade_));
    InMux I__9296 (
            .O(N__43963),
            .I(N__43960));
    LocalMux I__9295 (
            .O(N__43960),
            .I(n14887));
    InMux I__9294 (
            .O(N__43957),
            .I(N__43954));
    LocalMux I__9293 (
            .O(N__43954),
            .I(pwm_setpoint_23_N_171_22));
    InMux I__9292 (
            .O(N__43951),
            .I(N__43945));
    InMux I__9291 (
            .O(N__43950),
            .I(N__43945));
    LocalMux I__9290 (
            .O(N__43945),
            .I(N__43942));
    Odrv12 I__9289 (
            .O(N__43942),
            .I(pwm_setpoint_22));
    InMux I__9288 (
            .O(N__43939),
            .I(N__43936));
    LocalMux I__9287 (
            .O(N__43936),
            .I(N__43933));
    Odrv4 I__9286 (
            .O(N__43933),
            .I(pwm_setpoint_23_N_171_17));
    InMux I__9285 (
            .O(N__43930),
            .I(N__43927));
    LocalMux I__9284 (
            .O(N__43927),
            .I(n14870));
    InMux I__9283 (
            .O(N__43924),
            .I(N__43921));
    LocalMux I__9282 (
            .O(N__43921),
            .I(n14832));
    InMux I__9281 (
            .O(N__43918),
            .I(n12064));
    InMux I__9280 (
            .O(N__43915),
            .I(bfn_13_30_0_));
    InMux I__9279 (
            .O(N__43912),
            .I(n12066));
    InMux I__9278 (
            .O(N__43909),
            .I(n12067));
    InMux I__9277 (
            .O(N__43906),
            .I(N__43903));
    LocalMux I__9276 (
            .O(N__43903),
            .I(pwm_setpoint_23_N_171_19));
    InMux I__9275 (
            .O(N__43900),
            .I(n12068));
    InMux I__9274 (
            .O(N__43897),
            .I(N__43894));
    LocalMux I__9273 (
            .O(N__43894),
            .I(pwm_setpoint_23_N_171_20));
    InMux I__9272 (
            .O(N__43891),
            .I(n12069));
    InMux I__9271 (
            .O(N__43888),
            .I(N__43885));
    LocalMux I__9270 (
            .O(N__43885),
            .I(N__43882));
    Span4Mux_v I__9269 (
            .O(N__43882),
            .I(N__43879));
    Odrv4 I__9268 (
            .O(N__43879),
            .I(n4_adj_570));
    InMux I__9267 (
            .O(N__43876),
            .I(N__43873));
    LocalMux I__9266 (
            .O(N__43873),
            .I(N__43870));
    Span4Mux_v I__9265 (
            .O(N__43870),
            .I(N__43867));
    Odrv4 I__9264 (
            .O(N__43867),
            .I(pwm_setpoint_23_N_171_21));
    InMux I__9263 (
            .O(N__43864),
            .I(n12070));
    InMux I__9262 (
            .O(N__43861),
            .I(n12071));
    InMux I__9261 (
            .O(N__43858),
            .I(n12072));
    InMux I__9260 (
            .O(N__43855),
            .I(N__43852));
    LocalMux I__9259 (
            .O(N__43852),
            .I(N__43849));
    Odrv4 I__9258 (
            .O(N__43849),
            .I(pwm_setpoint_23));
    InMux I__9257 (
            .O(N__43846),
            .I(N__43843));
    LocalMux I__9256 (
            .O(N__43843),
            .I(n18_adj_584));
    InMux I__9255 (
            .O(N__43840),
            .I(n12056));
    InMux I__9254 (
            .O(N__43837),
            .I(N__43834));
    LocalMux I__9253 (
            .O(N__43834),
            .I(pwm_setpoint_23_N_171_8));
    InMux I__9252 (
            .O(N__43831),
            .I(bfn_13_29_0_));
    InMux I__9251 (
            .O(N__43828),
            .I(n12058));
    InMux I__9250 (
            .O(N__43825),
            .I(N__43822));
    LocalMux I__9249 (
            .O(N__43822),
            .I(N__43819));
    Odrv4 I__9248 (
            .O(N__43819),
            .I(n15_adj_581));
    InMux I__9247 (
            .O(N__43816),
            .I(N__43813));
    LocalMux I__9246 (
            .O(N__43813),
            .I(pwm_setpoint_23_N_171_10));
    InMux I__9245 (
            .O(N__43810),
            .I(n12059));
    InMux I__9244 (
            .O(N__43807),
            .I(N__43804));
    LocalMux I__9243 (
            .O(N__43804),
            .I(N__43801));
    Odrv4 I__9242 (
            .O(N__43801),
            .I(n14_adj_580));
    InMux I__9241 (
            .O(N__43798),
            .I(N__43795));
    LocalMux I__9240 (
            .O(N__43795),
            .I(pwm_setpoint_23_N_171_11));
    InMux I__9239 (
            .O(N__43792),
            .I(n12060));
    CascadeMux I__9238 (
            .O(N__43789),
            .I(N__43786));
    InMux I__9237 (
            .O(N__43786),
            .I(N__43783));
    LocalMux I__9236 (
            .O(N__43783),
            .I(pwm_setpoint_23_N_171_12));
    InMux I__9235 (
            .O(N__43780),
            .I(n12061));
    InMux I__9234 (
            .O(N__43777),
            .I(n12062));
    InMux I__9233 (
            .O(N__43774),
            .I(N__43771));
    LocalMux I__9232 (
            .O(N__43771),
            .I(N__43768));
    Odrv4 I__9231 (
            .O(N__43768),
            .I(n11_adj_577));
    InMux I__9230 (
            .O(N__43765),
            .I(n12063));
    InMux I__9229 (
            .O(N__43762),
            .I(N__43759));
    LocalMux I__9228 (
            .O(N__43759),
            .I(n25_adj_591));
    InMux I__9227 (
            .O(N__43756),
            .I(bfn_13_28_0_));
    InMux I__9226 (
            .O(N__43753),
            .I(n12050));
    InMux I__9225 (
            .O(N__43750),
            .I(N__43747));
    LocalMux I__9224 (
            .O(N__43747),
            .I(n23_adj_589));
    InMux I__9223 (
            .O(N__43744),
            .I(N__43741));
    LocalMux I__9222 (
            .O(N__43741),
            .I(pwm_setpoint_23_N_171_2));
    InMux I__9221 (
            .O(N__43738),
            .I(n12051));
    InMux I__9220 (
            .O(N__43735),
            .I(N__43732));
    LocalMux I__9219 (
            .O(N__43732),
            .I(pwm_setpoint_23_N_171_3));
    InMux I__9218 (
            .O(N__43729),
            .I(n12052));
    InMux I__9217 (
            .O(N__43726),
            .I(N__43723));
    LocalMux I__9216 (
            .O(N__43723),
            .I(N__43720));
    Span4Mux_v I__9215 (
            .O(N__43720),
            .I(N__43717));
    Odrv4 I__9214 (
            .O(N__43717),
            .I(n21_adj_587));
    InMux I__9213 (
            .O(N__43714),
            .I(N__43711));
    LocalMux I__9212 (
            .O(N__43711),
            .I(pwm_setpoint_23_N_171_4));
    InMux I__9211 (
            .O(N__43708),
            .I(n12053));
    InMux I__9210 (
            .O(N__43705),
            .I(N__43702));
    LocalMux I__9209 (
            .O(N__43702),
            .I(n20_adj_586));
    InMux I__9208 (
            .O(N__43699),
            .I(N__43696));
    LocalMux I__9207 (
            .O(N__43696),
            .I(N__43693));
    Odrv4 I__9206 (
            .O(N__43693),
            .I(pwm_setpoint_23_N_171_5));
    InMux I__9205 (
            .O(N__43690),
            .I(n12054));
    InMux I__9204 (
            .O(N__43687),
            .I(N__43684));
    LocalMux I__9203 (
            .O(N__43684),
            .I(n19_adj_585));
    InMux I__9202 (
            .O(N__43681),
            .I(N__43678));
    LocalMux I__9201 (
            .O(N__43678),
            .I(pwm_setpoint_23_N_171_6));
    InMux I__9200 (
            .O(N__43675),
            .I(n12055));
    InMux I__9199 (
            .O(N__43672),
            .I(N__43669));
    LocalMux I__9198 (
            .O(N__43669),
            .I(N__43665));
    CascadeMux I__9197 (
            .O(N__43668),
            .I(N__43662));
    Span4Mux_v I__9196 (
            .O(N__43665),
            .I(N__43658));
    InMux I__9195 (
            .O(N__43662),
            .I(N__43655));
    InMux I__9194 (
            .O(N__43661),
            .I(N__43652));
    Sp12to4 I__9193 (
            .O(N__43658),
            .I(N__43647));
    LocalMux I__9192 (
            .O(N__43655),
            .I(N__43647));
    LocalMux I__9191 (
            .O(N__43652),
            .I(n3206));
    Odrv12 I__9190 (
            .O(N__43647),
            .I(n3206));
    InMux I__9189 (
            .O(N__43642),
            .I(N__43639));
    LocalMux I__9188 (
            .O(N__43639),
            .I(N__43636));
    Span4Mux_h I__9187 (
            .O(N__43636),
            .I(N__43633));
    Odrv4 I__9186 (
            .O(N__43633),
            .I(n3273));
    InMux I__9185 (
            .O(N__43630),
            .I(n12549));
    InMux I__9184 (
            .O(N__43627),
            .I(N__43624));
    LocalMux I__9183 (
            .O(N__43624),
            .I(N__43621));
    Span4Mux_h I__9182 (
            .O(N__43621),
            .I(N__43616));
    InMux I__9181 (
            .O(N__43620),
            .I(N__43611));
    InMux I__9180 (
            .O(N__43619),
            .I(N__43611));
    Odrv4 I__9179 (
            .O(N__43616),
            .I(n3205));
    LocalMux I__9178 (
            .O(N__43611),
            .I(n3205));
    InMux I__9177 (
            .O(N__43606),
            .I(N__43603));
    LocalMux I__9176 (
            .O(N__43603),
            .I(N__43600));
    Span4Mux_v I__9175 (
            .O(N__43600),
            .I(N__43597));
    Odrv4 I__9174 (
            .O(N__43597),
            .I(n3272));
    InMux I__9173 (
            .O(N__43594),
            .I(n12550));
    InMux I__9172 (
            .O(N__43591),
            .I(N__43588));
    LocalMux I__9171 (
            .O(N__43588),
            .I(N__43584));
    InMux I__9170 (
            .O(N__43587),
            .I(N__43581));
    Span12Mux_s7_v I__9169 (
            .O(N__43584),
            .I(N__43578));
    LocalMux I__9168 (
            .O(N__43581),
            .I(n15163));
    Odrv12 I__9167 (
            .O(N__43578),
            .I(n15163));
    InMux I__9166 (
            .O(N__43573),
            .I(n12551));
    InMux I__9165 (
            .O(N__43570),
            .I(N__43567));
    LocalMux I__9164 (
            .O(N__43567),
            .I(N__43564));
    Span4Mux_h I__9163 (
            .O(N__43564),
            .I(N__43561));
    Odrv4 I__9162 (
            .O(N__43561),
            .I(n14461));
    InMux I__9161 (
            .O(N__43558),
            .I(N__43555));
    LocalMux I__9160 (
            .O(N__43555),
            .I(N__43552));
    Span4Mux_v I__9159 (
            .O(N__43552),
            .I(N__43549));
    Odrv4 I__9158 (
            .O(N__43549),
            .I(encoder0_position_scaled_3));
    InMux I__9157 (
            .O(N__43546),
            .I(N__43541));
    InMux I__9156 (
            .O(N__43545),
            .I(N__43538));
    InMux I__9155 (
            .O(N__43544),
            .I(N__43535));
    LocalMux I__9154 (
            .O(N__43541),
            .I(dti_counter_2));
    LocalMux I__9153 (
            .O(N__43538),
            .I(dti_counter_2));
    LocalMux I__9152 (
            .O(N__43535),
            .I(dti_counter_2));
    CascadeMux I__9151 (
            .O(N__43528),
            .I(N__43524));
    InMux I__9150 (
            .O(N__43527),
            .I(N__43520));
    InMux I__9149 (
            .O(N__43524),
            .I(N__43517));
    InMux I__9148 (
            .O(N__43523),
            .I(N__43514));
    LocalMux I__9147 (
            .O(N__43520),
            .I(dti_counter_1));
    LocalMux I__9146 (
            .O(N__43517),
            .I(dti_counter_1));
    LocalMux I__9145 (
            .O(N__43514),
            .I(dti_counter_1));
    InMux I__9144 (
            .O(N__43507),
            .I(N__43504));
    LocalMux I__9143 (
            .O(N__43504),
            .I(n10_adj_680));
    InMux I__9142 (
            .O(N__43501),
            .I(N__43498));
    LocalMux I__9141 (
            .O(N__43498),
            .I(n3281));
    InMux I__9140 (
            .O(N__43495),
            .I(n12541));
    InMux I__9139 (
            .O(N__43492),
            .I(N__43489));
    LocalMux I__9138 (
            .O(N__43489),
            .I(n3280));
    InMux I__9137 (
            .O(N__43486),
            .I(n12542));
    InMux I__9136 (
            .O(N__43483),
            .I(N__43479));
    InMux I__9135 (
            .O(N__43482),
            .I(N__43475));
    LocalMux I__9134 (
            .O(N__43479),
            .I(N__43472));
    InMux I__9133 (
            .O(N__43478),
            .I(N__43469));
    LocalMux I__9132 (
            .O(N__43475),
            .I(N__43466));
    Span4Mux_v I__9131 (
            .O(N__43472),
            .I(N__43463));
    LocalMux I__9130 (
            .O(N__43469),
            .I(N__43460));
    Odrv4 I__9129 (
            .O(N__43466),
            .I(n3212));
    Odrv4 I__9128 (
            .O(N__43463),
            .I(n3212));
    Odrv4 I__9127 (
            .O(N__43460),
            .I(n3212));
    InMux I__9126 (
            .O(N__43453),
            .I(N__43450));
    LocalMux I__9125 (
            .O(N__43450),
            .I(N__43447));
    Odrv4 I__9124 (
            .O(N__43447),
            .I(n3279));
    InMux I__9123 (
            .O(N__43444),
            .I(n12543));
    InMux I__9122 (
            .O(N__43441),
            .I(N__43437));
    InMux I__9121 (
            .O(N__43440),
            .I(N__43434));
    LocalMux I__9120 (
            .O(N__43437),
            .I(N__43430));
    LocalMux I__9119 (
            .O(N__43434),
            .I(N__43427));
    InMux I__9118 (
            .O(N__43433),
            .I(N__43424));
    Odrv4 I__9117 (
            .O(N__43430),
            .I(n3211));
    Odrv4 I__9116 (
            .O(N__43427),
            .I(n3211));
    LocalMux I__9115 (
            .O(N__43424),
            .I(n3211));
    InMux I__9114 (
            .O(N__43417),
            .I(N__43414));
    LocalMux I__9113 (
            .O(N__43414),
            .I(N__43411));
    Span4Mux_v I__9112 (
            .O(N__43411),
            .I(N__43408));
    Odrv4 I__9111 (
            .O(N__43408),
            .I(n3278));
    InMux I__9110 (
            .O(N__43405),
            .I(bfn_13_26_0_));
    InMux I__9109 (
            .O(N__43402),
            .I(N__43398));
    CascadeMux I__9108 (
            .O(N__43401),
            .I(N__43395));
    LocalMux I__9107 (
            .O(N__43398),
            .I(N__43391));
    InMux I__9106 (
            .O(N__43395),
            .I(N__43388));
    InMux I__9105 (
            .O(N__43394),
            .I(N__43385));
    Span4Mux_v I__9104 (
            .O(N__43391),
            .I(N__43380));
    LocalMux I__9103 (
            .O(N__43388),
            .I(N__43380));
    LocalMux I__9102 (
            .O(N__43385),
            .I(n3210));
    Odrv4 I__9101 (
            .O(N__43380),
            .I(n3210));
    InMux I__9100 (
            .O(N__43375),
            .I(N__43372));
    LocalMux I__9099 (
            .O(N__43372),
            .I(N__43369));
    Span4Mux_v I__9098 (
            .O(N__43369),
            .I(N__43366));
    Odrv4 I__9097 (
            .O(N__43366),
            .I(n3277));
    InMux I__9096 (
            .O(N__43363),
            .I(n12545));
    InMux I__9095 (
            .O(N__43360),
            .I(N__43357));
    LocalMux I__9094 (
            .O(N__43357),
            .I(N__43354));
    Span4Mux_h I__9093 (
            .O(N__43354),
            .I(N__43351));
    Odrv4 I__9092 (
            .O(N__43351),
            .I(n3276));
    InMux I__9091 (
            .O(N__43348),
            .I(n12546));
    InMux I__9090 (
            .O(N__43345),
            .I(N__43342));
    LocalMux I__9089 (
            .O(N__43342),
            .I(N__43338));
    InMux I__9088 (
            .O(N__43341),
            .I(N__43334));
    Span4Mux_h I__9087 (
            .O(N__43338),
            .I(N__43331));
    InMux I__9086 (
            .O(N__43337),
            .I(N__43328));
    LocalMux I__9085 (
            .O(N__43334),
            .I(n3208));
    Odrv4 I__9084 (
            .O(N__43331),
            .I(n3208));
    LocalMux I__9083 (
            .O(N__43328),
            .I(n3208));
    InMux I__9082 (
            .O(N__43321),
            .I(N__43318));
    LocalMux I__9081 (
            .O(N__43318),
            .I(N__43315));
    Span4Mux_h I__9080 (
            .O(N__43315),
            .I(N__43312));
    Odrv4 I__9079 (
            .O(N__43312),
            .I(n3275));
    InMux I__9078 (
            .O(N__43309),
            .I(n12547));
    InMux I__9077 (
            .O(N__43306),
            .I(N__43303));
    LocalMux I__9076 (
            .O(N__43303),
            .I(N__43299));
    InMux I__9075 (
            .O(N__43302),
            .I(N__43295));
    Span4Mux_h I__9074 (
            .O(N__43299),
            .I(N__43292));
    InMux I__9073 (
            .O(N__43298),
            .I(N__43289));
    LocalMux I__9072 (
            .O(N__43295),
            .I(n3207));
    Odrv4 I__9071 (
            .O(N__43292),
            .I(n3207));
    LocalMux I__9070 (
            .O(N__43289),
            .I(n3207));
    InMux I__9069 (
            .O(N__43282),
            .I(N__43279));
    LocalMux I__9068 (
            .O(N__43279),
            .I(N__43276));
    Span4Mux_h I__9067 (
            .O(N__43276),
            .I(N__43273));
    Odrv4 I__9066 (
            .O(N__43273),
            .I(n3274));
    InMux I__9065 (
            .O(N__43270),
            .I(n12548));
    InMux I__9064 (
            .O(N__43267),
            .I(n12533));
    InMux I__9063 (
            .O(N__43264),
            .I(N__43261));
    LocalMux I__9062 (
            .O(N__43261),
            .I(n3288));
    InMux I__9061 (
            .O(N__43258),
            .I(n12534));
    InMux I__9060 (
            .O(N__43255),
            .I(n12535));
    InMux I__9059 (
            .O(N__43252),
            .I(bfn_13_25_0_));
    InMux I__9058 (
            .O(N__43249),
            .I(N__43246));
    LocalMux I__9057 (
            .O(N__43246),
            .I(n3285));
    InMux I__9056 (
            .O(N__43243),
            .I(n12537));
    CascadeMux I__9055 (
            .O(N__43240),
            .I(N__43237));
    InMux I__9054 (
            .O(N__43237),
            .I(N__43233));
    InMux I__9053 (
            .O(N__43236),
            .I(N__43230));
    LocalMux I__9052 (
            .O(N__43233),
            .I(N__43224));
    LocalMux I__9051 (
            .O(N__43230),
            .I(N__43224));
    InMux I__9050 (
            .O(N__43229),
            .I(N__43221));
    Odrv4 I__9049 (
            .O(N__43224),
            .I(n3217));
    LocalMux I__9048 (
            .O(N__43221),
            .I(n3217));
    InMux I__9047 (
            .O(N__43216),
            .I(N__43213));
    LocalMux I__9046 (
            .O(N__43213),
            .I(n3284));
    InMux I__9045 (
            .O(N__43210),
            .I(n12538));
    InMux I__9044 (
            .O(N__43207),
            .I(N__43204));
    LocalMux I__9043 (
            .O(N__43204),
            .I(N__43200));
    InMux I__9042 (
            .O(N__43203),
            .I(N__43196));
    Span4Mux_v I__9041 (
            .O(N__43200),
            .I(N__43193));
    InMux I__9040 (
            .O(N__43199),
            .I(N__43190));
    LocalMux I__9039 (
            .O(N__43196),
            .I(n3216));
    Odrv4 I__9038 (
            .O(N__43193),
            .I(n3216));
    LocalMux I__9037 (
            .O(N__43190),
            .I(n3216));
    InMux I__9036 (
            .O(N__43183),
            .I(N__43180));
    LocalMux I__9035 (
            .O(N__43180),
            .I(N__43177));
    Odrv4 I__9034 (
            .O(N__43177),
            .I(n3283));
    InMux I__9033 (
            .O(N__43174),
            .I(n12539));
    InMux I__9032 (
            .O(N__43171),
            .I(N__43168));
    LocalMux I__9031 (
            .O(N__43168),
            .I(N__43163));
    InMux I__9030 (
            .O(N__43167),
            .I(N__43160));
    InMux I__9029 (
            .O(N__43166),
            .I(N__43157));
    Span4Mux_v I__9028 (
            .O(N__43163),
            .I(N__43152));
    LocalMux I__9027 (
            .O(N__43160),
            .I(N__43152));
    LocalMux I__9026 (
            .O(N__43157),
            .I(N__43149));
    Span4Mux_v I__9025 (
            .O(N__43152),
            .I(N__43146));
    Odrv12 I__9024 (
            .O(N__43149),
            .I(n3215));
    Odrv4 I__9023 (
            .O(N__43146),
            .I(n3215));
    InMux I__9022 (
            .O(N__43141),
            .I(N__43138));
    LocalMux I__9021 (
            .O(N__43138),
            .I(n3282));
    InMux I__9020 (
            .O(N__43135),
            .I(n12540));
    InMux I__9019 (
            .O(N__43132),
            .I(N__43127));
    InMux I__9018 (
            .O(N__43131),
            .I(N__43124));
    InMux I__9017 (
            .O(N__43130),
            .I(N__43121));
    LocalMux I__9016 (
            .O(N__43127),
            .I(N__43118));
    LocalMux I__9015 (
            .O(N__43124),
            .I(n3214));
    LocalMux I__9014 (
            .O(N__43121),
            .I(n3214));
    Odrv4 I__9013 (
            .O(N__43118),
            .I(n3214));
    InMux I__9012 (
            .O(N__43111),
            .I(N__43108));
    LocalMux I__9011 (
            .O(N__43108),
            .I(n3298));
    CascadeMux I__9010 (
            .O(N__43105),
            .I(N__43101));
    InMux I__9009 (
            .O(N__43104),
            .I(N__43098));
    InMux I__9008 (
            .O(N__43101),
            .I(N__43095));
    LocalMux I__9007 (
            .O(N__43098),
            .I(N__43091));
    LocalMux I__9006 (
            .O(N__43095),
            .I(N__43088));
    InMux I__9005 (
            .O(N__43094),
            .I(N__43085));
    Odrv4 I__9004 (
            .O(N__43091),
            .I(n3230));
    Odrv12 I__9003 (
            .O(N__43088),
            .I(n3230));
    LocalMux I__9002 (
            .O(N__43085),
            .I(n3230));
    InMux I__9001 (
            .O(N__43078),
            .I(N__43075));
    LocalMux I__9000 (
            .O(N__43075),
            .I(N__43072));
    Span4Mux_h I__8999 (
            .O(N__43072),
            .I(N__43069));
    Odrv4 I__8998 (
            .O(N__43069),
            .I(n14697));
    InMux I__8997 (
            .O(N__43066),
            .I(n12525));
    InMux I__8996 (
            .O(N__43063),
            .I(n12526));
    InMux I__8995 (
            .O(N__43060),
            .I(n12527));
    InMux I__8994 (
            .O(N__43057),
            .I(bfn_13_24_0_));
    InMux I__8993 (
            .O(N__43054),
            .I(N__43051));
    LocalMux I__8992 (
            .O(N__43051),
            .I(n3293));
    InMux I__8991 (
            .O(N__43048),
            .I(n12529));
    InMux I__8990 (
            .O(N__43045),
            .I(n12530));
    CascadeMux I__8989 (
            .O(N__43042),
            .I(N__43039));
    InMux I__8988 (
            .O(N__43039),
            .I(N__43036));
    LocalMux I__8987 (
            .O(N__43036),
            .I(n3291));
    InMux I__8986 (
            .O(N__43033),
            .I(n12531));
    CascadeMux I__8985 (
            .O(N__43030),
            .I(N__43027));
    InMux I__8984 (
            .O(N__43027),
            .I(N__43024));
    LocalMux I__8983 (
            .O(N__43024),
            .I(n3290));
    InMux I__8982 (
            .O(N__43021),
            .I(n12532));
    CascadeMux I__8981 (
            .O(N__43018),
            .I(n3014_cascade_));
    InMux I__8980 (
            .O(N__43015),
            .I(N__43012));
    LocalMux I__8979 (
            .O(N__43012),
            .I(n14408));
    InMux I__8978 (
            .O(N__43009),
            .I(N__43006));
    LocalMux I__8977 (
            .O(N__43006),
            .I(N__42990));
    InMux I__8976 (
            .O(N__43005),
            .I(N__42981));
    InMux I__8975 (
            .O(N__43004),
            .I(N__42981));
    InMux I__8974 (
            .O(N__43003),
            .I(N__42981));
    InMux I__8973 (
            .O(N__43002),
            .I(N__42981));
    CascadeMux I__8972 (
            .O(N__43001),
            .I(N__42976));
    CascadeMux I__8971 (
            .O(N__43000),
            .I(N__42972));
    CascadeMux I__8970 (
            .O(N__42999),
            .I(N__42968));
    CascadeMux I__8969 (
            .O(N__42998),
            .I(N__42965));
    CascadeMux I__8968 (
            .O(N__42997),
            .I(N__42957));
    CascadeMux I__8967 (
            .O(N__42996),
            .I(N__42954));
    CascadeMux I__8966 (
            .O(N__42995),
            .I(N__42950));
    CascadeMux I__8965 (
            .O(N__42994),
            .I(N__42947));
    CascadeMux I__8964 (
            .O(N__42993),
            .I(N__42942));
    Span4Mux_v I__8963 (
            .O(N__42990),
            .I(N__42937));
    LocalMux I__8962 (
            .O(N__42981),
            .I(N__42934));
    InMux I__8961 (
            .O(N__42980),
            .I(N__42931));
    InMux I__8960 (
            .O(N__42979),
            .I(N__42920));
    InMux I__8959 (
            .O(N__42976),
            .I(N__42920));
    InMux I__8958 (
            .O(N__42975),
            .I(N__42920));
    InMux I__8957 (
            .O(N__42972),
            .I(N__42920));
    InMux I__8956 (
            .O(N__42971),
            .I(N__42920));
    InMux I__8955 (
            .O(N__42968),
            .I(N__42913));
    InMux I__8954 (
            .O(N__42965),
            .I(N__42913));
    InMux I__8953 (
            .O(N__42964),
            .I(N__42913));
    InMux I__8952 (
            .O(N__42963),
            .I(N__42906));
    InMux I__8951 (
            .O(N__42962),
            .I(N__42906));
    InMux I__8950 (
            .O(N__42961),
            .I(N__42906));
    InMux I__8949 (
            .O(N__42960),
            .I(N__42897));
    InMux I__8948 (
            .O(N__42957),
            .I(N__42897));
    InMux I__8947 (
            .O(N__42954),
            .I(N__42897));
    InMux I__8946 (
            .O(N__42953),
            .I(N__42897));
    InMux I__8945 (
            .O(N__42950),
            .I(N__42888));
    InMux I__8944 (
            .O(N__42947),
            .I(N__42888));
    InMux I__8943 (
            .O(N__42946),
            .I(N__42888));
    InMux I__8942 (
            .O(N__42945),
            .I(N__42888));
    InMux I__8941 (
            .O(N__42942),
            .I(N__42881));
    InMux I__8940 (
            .O(N__42941),
            .I(N__42881));
    InMux I__8939 (
            .O(N__42940),
            .I(N__42881));
    Odrv4 I__8938 (
            .O(N__42937),
            .I(n2940));
    Odrv4 I__8937 (
            .O(N__42934),
            .I(n2940));
    LocalMux I__8936 (
            .O(N__42931),
            .I(n2940));
    LocalMux I__8935 (
            .O(N__42920),
            .I(n2940));
    LocalMux I__8934 (
            .O(N__42913),
            .I(n2940));
    LocalMux I__8933 (
            .O(N__42906),
            .I(n2940));
    LocalMux I__8932 (
            .O(N__42897),
            .I(n2940));
    LocalMux I__8931 (
            .O(N__42888),
            .I(n2940));
    LocalMux I__8930 (
            .O(N__42881),
            .I(n2940));
    InMux I__8929 (
            .O(N__42862),
            .I(N__42859));
    LocalMux I__8928 (
            .O(N__42859),
            .I(N__42856));
    Odrv4 I__8927 (
            .O(N__42856),
            .I(n2989));
    CascadeMux I__8926 (
            .O(N__42853),
            .I(n3021_cascade_));
    InMux I__8925 (
            .O(N__42850),
            .I(N__42846));
    InMux I__8924 (
            .O(N__42849),
            .I(N__42843));
    LocalMux I__8923 (
            .O(N__42846),
            .I(N__42840));
    LocalMux I__8922 (
            .O(N__42843),
            .I(N__42837));
    Span4Mux_v I__8921 (
            .O(N__42840),
            .I(N__42834));
    Span4Mux_v I__8920 (
            .O(N__42837),
            .I(N__42829));
    Span4Mux_h I__8919 (
            .O(N__42834),
            .I(N__42829));
    Span4Mux_h I__8918 (
            .O(N__42829),
            .I(N__42826));
    Odrv4 I__8917 (
            .O(N__42826),
            .I(n319));
    InMux I__8916 (
            .O(N__42823),
            .I(N__42819));
    InMux I__8915 (
            .O(N__42822),
            .I(N__42815));
    LocalMux I__8914 (
            .O(N__42819),
            .I(N__42812));
    InMux I__8913 (
            .O(N__42818),
            .I(N__42809));
    LocalMux I__8912 (
            .O(N__42815),
            .I(N__42806));
    Span4Mux_v I__8911 (
            .O(N__42812),
            .I(N__42803));
    LocalMux I__8910 (
            .O(N__42809),
            .I(N__42800));
    Span4Mux_h I__8909 (
            .O(N__42806),
            .I(N__42797));
    Span4Mux_h I__8908 (
            .O(N__42803),
            .I(N__42792));
    Span4Mux_v I__8907 (
            .O(N__42800),
            .I(N__42792));
    Odrv4 I__8906 (
            .O(N__42797),
            .I(n318));
    Odrv4 I__8905 (
            .O(N__42792),
            .I(n318));
    CascadeMux I__8904 (
            .O(N__42787),
            .I(N__42784));
    InMux I__8903 (
            .O(N__42784),
            .I(N__42781));
    LocalMux I__8902 (
            .O(N__42781),
            .I(N__42778));
    Span4Mux_h I__8901 (
            .O(N__42778),
            .I(N__42775));
    Odrv4 I__8900 (
            .O(N__42775),
            .I(n3301));
    InMux I__8899 (
            .O(N__42772),
            .I(n12521));
    InMux I__8898 (
            .O(N__42769),
            .I(N__42766));
    LocalMux I__8897 (
            .O(N__42766),
            .I(N__42762));
    InMux I__8896 (
            .O(N__42765),
            .I(N__42758));
    Span4Mux_h I__8895 (
            .O(N__42762),
            .I(N__42755));
    InMux I__8894 (
            .O(N__42761),
            .I(N__42752));
    LocalMux I__8893 (
            .O(N__42758),
            .I(n3233));
    Odrv4 I__8892 (
            .O(N__42755),
            .I(n3233));
    LocalMux I__8891 (
            .O(N__42752),
            .I(n3233));
    InMux I__8890 (
            .O(N__42745),
            .I(N__42742));
    LocalMux I__8889 (
            .O(N__42742),
            .I(N__42739));
    Span4Mux_v I__8888 (
            .O(N__42739),
            .I(N__42736));
    Span4Mux_h I__8887 (
            .O(N__42736),
            .I(N__42733));
    Odrv4 I__8886 (
            .O(N__42733),
            .I(n3300));
    InMux I__8885 (
            .O(N__42730),
            .I(n12522));
    InMux I__8884 (
            .O(N__42727),
            .I(N__42724));
    LocalMux I__8883 (
            .O(N__42724),
            .I(N__42720));
    InMux I__8882 (
            .O(N__42723),
            .I(N__42717));
    Span4Mux_v I__8881 (
            .O(N__42720),
            .I(N__42714));
    LocalMux I__8880 (
            .O(N__42717),
            .I(N__42711));
    Odrv4 I__8879 (
            .O(N__42714),
            .I(n3232));
    Odrv12 I__8878 (
            .O(N__42711),
            .I(n3232));
    InMux I__8877 (
            .O(N__42706),
            .I(N__42703));
    LocalMux I__8876 (
            .O(N__42703),
            .I(N__42700));
    Span4Mux_v I__8875 (
            .O(N__42700),
            .I(N__42697));
    Odrv4 I__8874 (
            .O(N__42697),
            .I(n3299));
    InMux I__8873 (
            .O(N__42694),
            .I(n12523));
    InMux I__8872 (
            .O(N__42691),
            .I(N__42688));
    LocalMux I__8871 (
            .O(N__42688),
            .I(N__42684));
    InMux I__8870 (
            .O(N__42687),
            .I(N__42680));
    Span4Mux_h I__8869 (
            .O(N__42684),
            .I(N__42677));
    InMux I__8868 (
            .O(N__42683),
            .I(N__42674));
    LocalMux I__8867 (
            .O(N__42680),
            .I(n3231));
    Odrv4 I__8866 (
            .O(N__42677),
            .I(n3231));
    LocalMux I__8865 (
            .O(N__42674),
            .I(n3231));
    InMux I__8864 (
            .O(N__42667),
            .I(n12524));
    InMux I__8863 (
            .O(N__42664),
            .I(N__42661));
    LocalMux I__8862 (
            .O(N__42661),
            .I(N__42658));
    Span4Mux_v I__8861 (
            .O(N__42658),
            .I(N__42655));
    Odrv4 I__8860 (
            .O(N__42655),
            .I(n2992));
    InMux I__8859 (
            .O(N__42652),
            .I(N__42649));
    LocalMux I__8858 (
            .O(N__42649),
            .I(N__42646));
    Span4Mux_v I__8857 (
            .O(N__42646),
            .I(N__42643));
    Odrv4 I__8856 (
            .O(N__42643),
            .I(n2991));
    CascadeMux I__8855 (
            .O(N__42640),
            .I(n3023_cascade_));
    InMux I__8854 (
            .O(N__42637),
            .I(N__42634));
    LocalMux I__8853 (
            .O(N__42634),
            .I(n14320));
    InMux I__8852 (
            .O(N__42631),
            .I(N__42628));
    LocalMux I__8851 (
            .O(N__42628),
            .I(N__42625));
    Odrv12 I__8850 (
            .O(N__42625),
            .I(n2995));
    CascadeMux I__8849 (
            .O(N__42622),
            .I(N__42619));
    InMux I__8848 (
            .O(N__42619),
            .I(N__42616));
    LocalMux I__8847 (
            .O(N__42616),
            .I(N__42613));
    Span4Mux_h I__8846 (
            .O(N__42613),
            .I(N__42610));
    Odrv4 I__8845 (
            .O(N__42610),
            .I(n2994));
    InMux I__8844 (
            .O(N__42607),
            .I(N__42603));
    InMux I__8843 (
            .O(N__42606),
            .I(N__42600));
    LocalMux I__8842 (
            .O(N__42603),
            .I(N__42595));
    LocalMux I__8841 (
            .O(N__42600),
            .I(N__42595));
    Span4Mux_h I__8840 (
            .O(N__42595),
            .I(N__42591));
    InMux I__8839 (
            .O(N__42594),
            .I(N__42588));
    Odrv4 I__8838 (
            .O(N__42591),
            .I(n2913));
    LocalMux I__8837 (
            .O(N__42588),
            .I(n2913));
    InMux I__8836 (
            .O(N__42583),
            .I(N__42580));
    LocalMux I__8835 (
            .O(N__42580),
            .I(N__42577));
    Odrv12 I__8834 (
            .O(N__42577),
            .I(n2990));
    CascadeMux I__8833 (
            .O(N__42574),
            .I(N__42571));
    InMux I__8832 (
            .O(N__42571),
            .I(N__42568));
    LocalMux I__8831 (
            .O(N__42568),
            .I(N__42565));
    Span4Mux_h I__8830 (
            .O(N__42565),
            .I(N__42562));
    Odrv4 I__8829 (
            .O(N__42562),
            .I(n2982));
    InMux I__8828 (
            .O(N__42559),
            .I(N__42555));
    InMux I__8827 (
            .O(N__42558),
            .I(N__42552));
    LocalMux I__8826 (
            .O(N__42555),
            .I(N__42549));
    LocalMux I__8825 (
            .O(N__42552),
            .I(N__42545));
    Span4Mux_v I__8824 (
            .O(N__42549),
            .I(N__42542));
    InMux I__8823 (
            .O(N__42548),
            .I(N__42539));
    Odrv4 I__8822 (
            .O(N__42545),
            .I(n2915));
    Odrv4 I__8821 (
            .O(N__42542),
            .I(n2915));
    LocalMux I__8820 (
            .O(N__42539),
            .I(n2915));
    InMux I__8819 (
            .O(N__42532),
            .I(N__42528));
    InMux I__8818 (
            .O(N__42531),
            .I(N__42525));
    LocalMux I__8817 (
            .O(N__42528),
            .I(N__42519));
    LocalMux I__8816 (
            .O(N__42525),
            .I(N__42519));
    InMux I__8815 (
            .O(N__42524),
            .I(N__42516));
    Span4Mux_v I__8814 (
            .O(N__42519),
            .I(N__42511));
    LocalMux I__8813 (
            .O(N__42516),
            .I(N__42511));
    Odrv4 I__8812 (
            .O(N__42511),
            .I(n2916));
    CascadeMux I__8811 (
            .O(N__42508),
            .I(n13934_cascade_));
    InMux I__8810 (
            .O(N__42505),
            .I(N__42502));
    LocalMux I__8809 (
            .O(N__42502),
            .I(N__42499));
    Odrv4 I__8808 (
            .O(N__42499),
            .I(n13942));
    InMux I__8807 (
            .O(N__42496),
            .I(N__42493));
    LocalMux I__8806 (
            .O(N__42493),
            .I(N__42490));
    Span4Mux_h I__8805 (
            .O(N__42490),
            .I(N__42487));
    Odrv4 I__8804 (
            .O(N__42487),
            .I(n2679));
    CascadeMux I__8803 (
            .O(N__42484),
            .I(N__42481));
    InMux I__8802 (
            .O(N__42481),
            .I(N__42478));
    LocalMux I__8801 (
            .O(N__42478),
            .I(N__42475));
    Span4Mux_v I__8800 (
            .O(N__42475),
            .I(N__42470));
    InMux I__8799 (
            .O(N__42474),
            .I(N__42467));
    InMux I__8798 (
            .O(N__42473),
            .I(N__42464));
    Span4Mux_h I__8797 (
            .O(N__42470),
            .I(N__42461));
    LocalMux I__8796 (
            .O(N__42467),
            .I(N__42458));
    LocalMux I__8795 (
            .O(N__42464),
            .I(N__42455));
    Odrv4 I__8794 (
            .O(N__42461),
            .I(n2612));
    Odrv4 I__8793 (
            .O(N__42458),
            .I(n2612));
    Odrv4 I__8792 (
            .O(N__42455),
            .I(n2612));
    InMux I__8791 (
            .O(N__42448),
            .I(N__42445));
    LocalMux I__8790 (
            .O(N__42445),
            .I(N__42439));
    InMux I__8789 (
            .O(N__42444),
            .I(N__42436));
    InMux I__8788 (
            .O(N__42443),
            .I(N__42433));
    CascadeMux I__8787 (
            .O(N__42442),
            .I(N__42424));
    Span4Mux_v I__8786 (
            .O(N__42439),
            .I(N__42419));
    LocalMux I__8785 (
            .O(N__42436),
            .I(N__42416));
    LocalMux I__8784 (
            .O(N__42433),
            .I(N__42413));
    CascadeMux I__8783 (
            .O(N__42432),
            .I(N__42409));
    CascadeMux I__8782 (
            .O(N__42431),
            .I(N__42406));
    CascadeMux I__8781 (
            .O(N__42430),
            .I(N__42399));
    CascadeMux I__8780 (
            .O(N__42429),
            .I(N__42392));
    CascadeMux I__8779 (
            .O(N__42428),
            .I(N__42387));
    CascadeMux I__8778 (
            .O(N__42427),
            .I(N__42384));
    InMux I__8777 (
            .O(N__42424),
            .I(N__42375));
    InMux I__8776 (
            .O(N__42423),
            .I(N__42375));
    InMux I__8775 (
            .O(N__42422),
            .I(N__42375));
    Span4Mux_v I__8774 (
            .O(N__42419),
            .I(N__42368));
    Span4Mux_v I__8773 (
            .O(N__42416),
            .I(N__42368));
    Span4Mux_v I__8772 (
            .O(N__42413),
            .I(N__42368));
    InMux I__8771 (
            .O(N__42412),
            .I(N__42357));
    InMux I__8770 (
            .O(N__42409),
            .I(N__42357));
    InMux I__8769 (
            .O(N__42406),
            .I(N__42357));
    InMux I__8768 (
            .O(N__42405),
            .I(N__42357));
    InMux I__8767 (
            .O(N__42404),
            .I(N__42357));
    InMux I__8766 (
            .O(N__42403),
            .I(N__42346));
    InMux I__8765 (
            .O(N__42402),
            .I(N__42346));
    InMux I__8764 (
            .O(N__42399),
            .I(N__42346));
    InMux I__8763 (
            .O(N__42398),
            .I(N__42346));
    InMux I__8762 (
            .O(N__42397),
            .I(N__42346));
    InMux I__8761 (
            .O(N__42396),
            .I(N__42341));
    InMux I__8760 (
            .O(N__42395),
            .I(N__42341));
    InMux I__8759 (
            .O(N__42392),
            .I(N__42336));
    InMux I__8758 (
            .O(N__42391),
            .I(N__42336));
    InMux I__8757 (
            .O(N__42390),
            .I(N__42325));
    InMux I__8756 (
            .O(N__42387),
            .I(N__42325));
    InMux I__8755 (
            .O(N__42384),
            .I(N__42325));
    InMux I__8754 (
            .O(N__42383),
            .I(N__42325));
    InMux I__8753 (
            .O(N__42382),
            .I(N__42325));
    LocalMux I__8752 (
            .O(N__42375),
            .I(n2643));
    Odrv4 I__8751 (
            .O(N__42368),
            .I(n2643));
    LocalMux I__8750 (
            .O(N__42357),
            .I(n2643));
    LocalMux I__8749 (
            .O(N__42346),
            .I(n2643));
    LocalMux I__8748 (
            .O(N__42341),
            .I(n2643));
    LocalMux I__8747 (
            .O(N__42336),
            .I(n2643));
    LocalMux I__8746 (
            .O(N__42325),
            .I(n2643));
    CascadeMux I__8745 (
            .O(N__42310),
            .I(N__42306));
    CascadeMux I__8744 (
            .O(N__42309),
            .I(N__42302));
    InMux I__8743 (
            .O(N__42306),
            .I(N__42299));
    InMux I__8742 (
            .O(N__42305),
            .I(N__42296));
    InMux I__8741 (
            .O(N__42302),
            .I(N__42293));
    LocalMux I__8740 (
            .O(N__42299),
            .I(N__42288));
    LocalMux I__8739 (
            .O(N__42296),
            .I(N__42288));
    LocalMux I__8738 (
            .O(N__42293),
            .I(n2711));
    Odrv4 I__8737 (
            .O(N__42288),
            .I(n2711));
    InMux I__8736 (
            .O(N__42283),
            .I(N__42280));
    LocalMux I__8735 (
            .O(N__42280),
            .I(N__42277));
    Span4Mux_v I__8734 (
            .O(N__42277),
            .I(N__42274));
    Span4Mux_h I__8733 (
            .O(N__42274),
            .I(N__42270));
    InMux I__8732 (
            .O(N__42273),
            .I(N__42267));
    Odrv4 I__8731 (
            .O(N__42270),
            .I(n15467));
    LocalMux I__8730 (
            .O(N__42267),
            .I(n15467));
    InMux I__8729 (
            .O(N__42262),
            .I(N__42258));
    InMux I__8728 (
            .O(N__42261),
            .I(N__42255));
    LocalMux I__8727 (
            .O(N__42258),
            .I(N__42252));
    LocalMux I__8726 (
            .O(N__42255),
            .I(N__42249));
    Span4Mux_v I__8725 (
            .O(N__42252),
            .I(N__42245));
    Span4Mux_v I__8724 (
            .O(N__42249),
            .I(N__42242));
    InMux I__8723 (
            .O(N__42248),
            .I(N__42239));
    Odrv4 I__8722 (
            .O(N__42245),
            .I(n2909));
    Odrv4 I__8721 (
            .O(N__42242),
            .I(n2909));
    LocalMux I__8720 (
            .O(N__42239),
            .I(n2909));
    InMux I__8719 (
            .O(N__42232),
            .I(N__42228));
    InMux I__8718 (
            .O(N__42231),
            .I(N__42224));
    LocalMux I__8717 (
            .O(N__42228),
            .I(N__42221));
    InMux I__8716 (
            .O(N__42227),
            .I(N__42218));
    LocalMux I__8715 (
            .O(N__42224),
            .I(N__42215));
    Span4Mux_v I__8714 (
            .O(N__42221),
            .I(N__42212));
    LocalMux I__8713 (
            .O(N__42218),
            .I(N__42207));
    Span4Mux_v I__8712 (
            .O(N__42215),
            .I(N__42207));
    Odrv4 I__8711 (
            .O(N__42212),
            .I(n2713));
    Odrv4 I__8710 (
            .O(N__42207),
            .I(n2713));
    InMux I__8709 (
            .O(N__42202),
            .I(N__42199));
    LocalMux I__8708 (
            .O(N__42199),
            .I(n2780));
    CascadeMux I__8707 (
            .O(N__42196),
            .I(n14322_cascade_));
    CascadeMux I__8706 (
            .O(N__42193),
            .I(N__42190));
    InMux I__8705 (
            .O(N__42190),
            .I(N__42187));
    LocalMux I__8704 (
            .O(N__42187),
            .I(n14328));
    CascadeMux I__8703 (
            .O(N__42184),
            .I(N__42180));
    InMux I__8702 (
            .O(N__42183),
            .I(N__42177));
    InMux I__8701 (
            .O(N__42180),
            .I(N__42174));
    LocalMux I__8700 (
            .O(N__42177),
            .I(N__42168));
    LocalMux I__8699 (
            .O(N__42174),
            .I(N__42168));
    InMux I__8698 (
            .O(N__42173),
            .I(N__42165));
    Odrv12 I__8697 (
            .O(N__42168),
            .I(n2724));
    LocalMux I__8696 (
            .O(N__42165),
            .I(n2724));
    CascadeMux I__8695 (
            .O(N__42160),
            .I(N__42157));
    InMux I__8694 (
            .O(N__42157),
            .I(N__42154));
    LocalMux I__8693 (
            .O(N__42154),
            .I(N__42151));
    Odrv4 I__8692 (
            .O(N__42151),
            .I(n2791));
    InMux I__8691 (
            .O(N__42148),
            .I(N__42145));
    LocalMux I__8690 (
            .O(N__42145),
            .I(n2786));
    InMux I__8689 (
            .O(N__42142),
            .I(N__42139));
    LocalMux I__8688 (
            .O(N__42139),
            .I(N__42135));
    InMux I__8687 (
            .O(N__42138),
            .I(N__42132));
    Span4Mux_h I__8686 (
            .O(N__42135),
            .I(N__42126));
    LocalMux I__8685 (
            .O(N__42132),
            .I(N__42126));
    InMux I__8684 (
            .O(N__42131),
            .I(N__42123));
    Odrv4 I__8683 (
            .O(N__42126),
            .I(n2719));
    LocalMux I__8682 (
            .O(N__42123),
            .I(n2719));
    InMux I__8681 (
            .O(N__42118),
            .I(N__42114));
    InMux I__8680 (
            .O(N__42117),
            .I(N__42111));
    LocalMux I__8679 (
            .O(N__42114),
            .I(N__42106));
    LocalMux I__8678 (
            .O(N__42111),
            .I(N__42106));
    Span4Mux_v I__8677 (
            .O(N__42106),
            .I(N__42103));
    Odrv4 I__8676 (
            .O(N__42103),
            .I(n2921));
    CascadeMux I__8675 (
            .O(N__42100),
            .I(n2921_cascade_));
    InMux I__8674 (
            .O(N__42097),
            .I(N__42094));
    LocalMux I__8673 (
            .O(N__42094),
            .I(n2778));
    CascadeMux I__8672 (
            .O(N__42091),
            .I(N__42087));
    InMux I__8671 (
            .O(N__42090),
            .I(N__42084));
    InMux I__8670 (
            .O(N__42087),
            .I(N__42081));
    LocalMux I__8669 (
            .O(N__42084),
            .I(N__42078));
    LocalMux I__8668 (
            .O(N__42081),
            .I(N__42075));
    Span4Mux_h I__8667 (
            .O(N__42078),
            .I(N__42072));
    Span4Mux_v I__8666 (
            .O(N__42075),
            .I(N__42069));
    Odrv4 I__8665 (
            .O(N__42072),
            .I(n2917));
    Odrv4 I__8664 (
            .O(N__42069),
            .I(n2917));
    InMux I__8663 (
            .O(N__42064),
            .I(N__42060));
    CascadeMux I__8662 (
            .O(N__42063),
            .I(N__42057));
    LocalMux I__8661 (
            .O(N__42060),
            .I(N__42054));
    InMux I__8660 (
            .O(N__42057),
            .I(N__42050));
    Span4Mux_v I__8659 (
            .O(N__42054),
            .I(N__42047));
    InMux I__8658 (
            .O(N__42053),
            .I(N__42044));
    LocalMux I__8657 (
            .O(N__42050),
            .I(n2918));
    Odrv4 I__8656 (
            .O(N__42047),
            .I(n2918));
    LocalMux I__8655 (
            .O(N__42044),
            .I(n2918));
    InMux I__8654 (
            .O(N__42037),
            .I(N__42034));
    LocalMux I__8653 (
            .O(N__42034),
            .I(n13926));
    CascadeMux I__8652 (
            .O(N__42031),
            .I(n2917_cascade_));
    CascadeMux I__8651 (
            .O(N__42028),
            .I(N__42024));
    InMux I__8650 (
            .O(N__42027),
            .I(N__42021));
    InMux I__8649 (
            .O(N__42024),
            .I(N__42018));
    LocalMux I__8648 (
            .O(N__42021),
            .I(N__42015));
    LocalMux I__8647 (
            .O(N__42018),
            .I(N__42012));
    Span4Mux_v I__8646 (
            .O(N__42015),
            .I(N__42009));
    Span4Mux_h I__8645 (
            .O(N__42012),
            .I(N__42006));
    Span4Mux_h I__8644 (
            .O(N__42009),
            .I(N__42003));
    Odrv4 I__8643 (
            .O(N__42006),
            .I(n2709));
    Odrv4 I__8642 (
            .O(N__42003),
            .I(n2709));
    InMux I__8641 (
            .O(N__41998),
            .I(N__41995));
    LocalMux I__8640 (
            .O(N__41995),
            .I(n2798));
    CascadeMux I__8639 (
            .O(N__41992),
            .I(n2742_cascade_));
    InMux I__8638 (
            .O(N__41989),
            .I(N__41986));
    LocalMux I__8637 (
            .O(N__41986),
            .I(N__41982));
    CascadeMux I__8636 (
            .O(N__41985),
            .I(N__41978));
    Span4Mux_v I__8635 (
            .O(N__41982),
            .I(N__41975));
    InMux I__8634 (
            .O(N__41981),
            .I(N__41972));
    InMux I__8633 (
            .O(N__41978),
            .I(N__41969));
    Odrv4 I__8632 (
            .O(N__41975),
            .I(n2731));
    LocalMux I__8631 (
            .O(N__41972),
            .I(n2731));
    LocalMux I__8630 (
            .O(N__41969),
            .I(n2731));
    CascadeMux I__8629 (
            .O(N__41962),
            .I(N__41958));
    InMux I__8628 (
            .O(N__41961),
            .I(N__41955));
    InMux I__8627 (
            .O(N__41958),
            .I(N__41952));
    LocalMux I__8626 (
            .O(N__41955),
            .I(N__41946));
    LocalMux I__8625 (
            .O(N__41952),
            .I(N__41946));
    InMux I__8624 (
            .O(N__41951),
            .I(N__41943));
    Odrv4 I__8623 (
            .O(N__41946),
            .I(n2728));
    LocalMux I__8622 (
            .O(N__41943),
            .I(n2728));
    CascadeMux I__8621 (
            .O(N__41938),
            .I(N__41935));
    InMux I__8620 (
            .O(N__41935),
            .I(N__41932));
    LocalMux I__8619 (
            .O(N__41932),
            .I(n2795));
    CascadeMux I__8618 (
            .O(N__41929),
            .I(n14238_cascade_));
    CascadeMux I__8617 (
            .O(N__41926),
            .I(n14240_cascade_));
    CascadeMux I__8616 (
            .O(N__41923),
            .I(N__41920));
    InMux I__8615 (
            .O(N__41920),
            .I(N__41916));
    InMux I__8614 (
            .O(N__41919),
            .I(N__41913));
    LocalMux I__8613 (
            .O(N__41916),
            .I(N__41908));
    LocalMux I__8612 (
            .O(N__41913),
            .I(N__41908));
    Odrv4 I__8611 (
            .O(N__41908),
            .I(n2720));
    InMux I__8610 (
            .O(N__41905),
            .I(N__41902));
    LocalMux I__8609 (
            .O(N__41902),
            .I(N__41899));
    Odrv4 I__8608 (
            .O(N__41899),
            .I(n2787));
    InMux I__8607 (
            .O(N__41896),
            .I(N__41893));
    LocalMux I__8606 (
            .O(N__41893),
            .I(n2789));
    CascadeMux I__8605 (
            .O(N__41890),
            .I(N__41887));
    InMux I__8604 (
            .O(N__41887),
            .I(N__41883));
    CascadeMux I__8603 (
            .O(N__41886),
            .I(N__41880));
    LocalMux I__8602 (
            .O(N__41883),
            .I(N__41876));
    InMux I__8601 (
            .O(N__41880),
            .I(N__41873));
    InMux I__8600 (
            .O(N__41879),
            .I(N__41870));
    Odrv4 I__8599 (
            .O(N__41876),
            .I(n2722));
    LocalMux I__8598 (
            .O(N__41873),
            .I(n2722));
    LocalMux I__8597 (
            .O(N__41870),
            .I(n2722));
    InMux I__8596 (
            .O(N__41863),
            .I(N__41860));
    LocalMux I__8595 (
            .O(N__41860),
            .I(n2797));
    InMux I__8594 (
            .O(N__41857),
            .I(N__41853));
    CascadeMux I__8593 (
            .O(N__41856),
            .I(N__41849));
    LocalMux I__8592 (
            .O(N__41853),
            .I(N__41846));
    InMux I__8591 (
            .O(N__41852),
            .I(N__41843));
    InMux I__8590 (
            .O(N__41849),
            .I(N__41840));
    Odrv4 I__8589 (
            .O(N__41846),
            .I(n2730));
    LocalMux I__8588 (
            .O(N__41843),
            .I(n2730));
    LocalMux I__8587 (
            .O(N__41840),
            .I(n2730));
    CascadeMux I__8586 (
            .O(N__41833),
            .I(N__41829));
    InMux I__8585 (
            .O(N__41832),
            .I(N__41825));
    InMux I__8584 (
            .O(N__41829),
            .I(N__41820));
    InMux I__8583 (
            .O(N__41828),
            .I(N__41820));
    LocalMux I__8582 (
            .O(N__41825),
            .I(N__41817));
    LocalMux I__8581 (
            .O(N__41820),
            .I(N__41812));
    Span4Mux_h I__8580 (
            .O(N__41817),
            .I(N__41812));
    Odrv4 I__8579 (
            .O(N__41812),
            .I(n23_adj_618));
    CascadeMux I__8578 (
            .O(N__41809),
            .I(n14800_cascade_));
    InMux I__8577 (
            .O(N__41806),
            .I(N__41803));
    LocalMux I__8576 (
            .O(N__41803),
            .I(n19_adj_616));
    InMux I__8575 (
            .O(N__41800),
            .I(N__41794));
    InMux I__8574 (
            .O(N__41799),
            .I(N__41794));
    LocalMux I__8573 (
            .O(N__41794),
            .I(N__41791));
    Span4Mux_h I__8572 (
            .O(N__41791),
            .I(N__41788));
    Odrv4 I__8571 (
            .O(N__41788),
            .I(n17_adj_615));
    CascadeMux I__8570 (
            .O(N__41785),
            .I(N__41782));
    InMux I__8569 (
            .O(N__41782),
            .I(N__41779));
    LocalMux I__8568 (
            .O(N__41779),
            .I(N__41775));
    InMux I__8567 (
            .O(N__41778),
            .I(N__41772));
    Span4Mux_s2_v I__8566 (
            .O(N__41775),
            .I(N__41767));
    LocalMux I__8565 (
            .O(N__41772),
            .I(N__41767));
    Odrv4 I__8564 (
            .O(N__41767),
            .I(n9_adj_608));
    InMux I__8563 (
            .O(N__41764),
            .I(N__41758));
    InMux I__8562 (
            .O(N__41763),
            .I(N__41758));
    LocalMux I__8561 (
            .O(N__41758),
            .I(N__41755));
    Odrv4 I__8560 (
            .O(N__41755),
            .I(n21_adj_617));
    InMux I__8559 (
            .O(N__41752),
            .I(N__41749));
    LocalMux I__8558 (
            .O(N__41749),
            .I(N__41746));
    Odrv4 I__8557 (
            .O(N__41746),
            .I(n14734));
    InMux I__8556 (
            .O(N__41743),
            .I(N__41740));
    LocalMux I__8555 (
            .O(N__41740),
            .I(N__41737));
    Span4Mux_h I__8554 (
            .O(N__41737),
            .I(N__41734));
    Odrv4 I__8553 (
            .O(N__41734),
            .I(n14874));
    InMux I__8552 (
            .O(N__41731),
            .I(N__41728));
    LocalMux I__8551 (
            .O(N__41728),
            .I(N__41724));
    InMux I__8550 (
            .O(N__41727),
            .I(N__41721));
    Span4Mux_h I__8549 (
            .O(N__41724),
            .I(N__41716));
    LocalMux I__8548 (
            .O(N__41721),
            .I(N__41716));
    Odrv4 I__8547 (
            .O(N__41716),
            .I(pwm_setpoint_12));
    InMux I__8546 (
            .O(N__41713),
            .I(N__41708));
    InMux I__8545 (
            .O(N__41712),
            .I(N__41705));
    InMux I__8544 (
            .O(N__41711),
            .I(N__41702));
    LocalMux I__8543 (
            .O(N__41708),
            .I(N__41699));
    LocalMux I__8542 (
            .O(N__41705),
            .I(pwm_counter_12));
    LocalMux I__8541 (
            .O(N__41702),
            .I(pwm_counter_12));
    Odrv4 I__8540 (
            .O(N__41699),
            .I(pwm_counter_12));
    InMux I__8539 (
            .O(N__41692),
            .I(N__41686));
    InMux I__8538 (
            .O(N__41691),
            .I(N__41686));
    LocalMux I__8537 (
            .O(N__41686),
            .I(N__41682));
    InMux I__8536 (
            .O(N__41685),
            .I(N__41679));
    Odrv4 I__8535 (
            .O(N__41682),
            .I(n25_adj_620));
    LocalMux I__8534 (
            .O(N__41679),
            .I(n25_adj_620));
    InMux I__8533 (
            .O(N__41674),
            .I(N__41670));
    CascadeMux I__8532 (
            .O(N__41673),
            .I(N__41667));
    LocalMux I__8531 (
            .O(N__41670),
            .I(N__41663));
    InMux I__8530 (
            .O(N__41667),
            .I(N__41660));
    InMux I__8529 (
            .O(N__41666),
            .I(N__41657));
    Odrv4 I__8528 (
            .O(N__41663),
            .I(n2723));
    LocalMux I__8527 (
            .O(N__41660),
            .I(n2723));
    LocalMux I__8526 (
            .O(N__41657),
            .I(n2723));
    CascadeMux I__8525 (
            .O(N__41650),
            .I(N__41647));
    InMux I__8524 (
            .O(N__41647),
            .I(N__41644));
    LocalMux I__8523 (
            .O(N__41644),
            .I(n2790));
    CascadeMux I__8522 (
            .O(N__41641),
            .I(N__41638));
    InMux I__8521 (
            .O(N__41638),
            .I(N__41634));
    InMux I__8520 (
            .O(N__41637),
            .I(N__41631));
    LocalMux I__8519 (
            .O(N__41634),
            .I(N__41628));
    LocalMux I__8518 (
            .O(N__41631),
            .I(N__41625));
    Span4Mux_h I__8517 (
            .O(N__41628),
            .I(N__41622));
    Odrv4 I__8516 (
            .O(N__41625),
            .I(n2725));
    Odrv4 I__8515 (
            .O(N__41622),
            .I(n2725));
    InMux I__8514 (
            .O(N__41617),
            .I(N__41614));
    LocalMux I__8513 (
            .O(N__41614),
            .I(n2792));
    InMux I__8512 (
            .O(N__41611),
            .I(N__41608));
    LocalMux I__8511 (
            .O(N__41608),
            .I(N__41605));
    Odrv4 I__8510 (
            .O(N__41605),
            .I(n13403));
    InMux I__8509 (
            .O(N__41602),
            .I(N__41599));
    LocalMux I__8508 (
            .O(N__41599),
            .I(N__41596));
    Odrv4 I__8507 (
            .O(N__41596),
            .I(n14048));
    InMux I__8506 (
            .O(N__41593),
            .I(N__41590));
    LocalMux I__8505 (
            .O(N__41590),
            .I(N__41586));
    InMux I__8504 (
            .O(N__41589),
            .I(N__41583));
    Span4Mux_h I__8503 (
            .O(N__41586),
            .I(N__41580));
    LocalMux I__8502 (
            .O(N__41583),
            .I(n2714));
    Odrv4 I__8501 (
            .O(N__41580),
            .I(n2714));
    CascadeMux I__8500 (
            .O(N__41575),
            .I(n14054_cascade_));
    CascadeMux I__8499 (
            .O(N__41572),
            .I(N__41569));
    InMux I__8498 (
            .O(N__41569),
            .I(N__41564));
    InMux I__8497 (
            .O(N__41568),
            .I(N__41561));
    InMux I__8496 (
            .O(N__41567),
            .I(N__41558));
    LocalMux I__8495 (
            .O(N__41564),
            .I(N__41555));
    LocalMux I__8494 (
            .O(N__41561),
            .I(N__41552));
    LocalMux I__8493 (
            .O(N__41558),
            .I(N__41549));
    Span4Mux_v I__8492 (
            .O(N__41555),
            .I(N__41544));
    Span4Mux_v I__8491 (
            .O(N__41552),
            .I(N__41544));
    Odrv4 I__8490 (
            .O(N__41549),
            .I(n2710));
    Odrv4 I__8489 (
            .O(N__41544),
            .I(n2710));
    CascadeMux I__8488 (
            .O(N__41539),
            .I(n14060_cascade_));
    CascadeMux I__8487 (
            .O(N__41536),
            .I(\PWM.n13596_cascade_ ));
    InMux I__8486 (
            .O(N__41533),
            .I(N__41527));
    InMux I__8485 (
            .O(N__41532),
            .I(N__41524));
    InMux I__8484 (
            .O(N__41531),
            .I(N__41519));
    InMux I__8483 (
            .O(N__41530),
            .I(N__41519));
    LocalMux I__8482 (
            .O(N__41527),
            .I(pwm_counter_8));
    LocalMux I__8481 (
            .O(N__41524),
            .I(pwm_counter_8));
    LocalMux I__8480 (
            .O(N__41519),
            .I(pwm_counter_8));
    InMux I__8479 (
            .O(N__41512),
            .I(N__41509));
    LocalMux I__8478 (
            .O(N__41509),
            .I(N__41506));
    Span4Mux_h I__8477 (
            .O(N__41506),
            .I(N__41503));
    Odrv4 I__8476 (
            .O(N__41503),
            .I(\PWM.n26 ));
    InMux I__8475 (
            .O(N__41500),
            .I(N__41497));
    LocalMux I__8474 (
            .O(N__41497),
            .I(N__41493));
    InMux I__8473 (
            .O(N__41496),
            .I(N__41490));
    Span4Mux_h I__8472 (
            .O(N__41493),
            .I(N__41487));
    LocalMux I__8471 (
            .O(N__41490),
            .I(N__41484));
    Odrv4 I__8470 (
            .O(N__41487),
            .I(n4823));
    Odrv4 I__8469 (
            .O(N__41484),
            .I(n4823));
    CascadeMux I__8468 (
            .O(N__41479),
            .I(\PWM.n17_cascade_ ));
    InMux I__8467 (
            .O(N__41476),
            .I(N__41471));
    InMux I__8466 (
            .O(N__41475),
            .I(N__41468));
    InMux I__8465 (
            .O(N__41474),
            .I(N__41465));
    LocalMux I__8464 (
            .O(N__41471),
            .I(N__41462));
    LocalMux I__8463 (
            .O(N__41468),
            .I(pwm_counter_31));
    LocalMux I__8462 (
            .O(N__41465),
            .I(pwm_counter_31));
    Odrv4 I__8461 (
            .O(N__41462),
            .I(pwm_counter_31));
    CascadeMux I__8460 (
            .O(N__41455),
            .I(\PWM.n29_cascade_ ));
    InMux I__8459 (
            .O(N__41452),
            .I(N__41449));
    LocalMux I__8458 (
            .O(N__41449),
            .I(N__41446));
    Span4Mux_s2_v I__8457 (
            .O(N__41446),
            .I(N__41443));
    Odrv4 I__8456 (
            .O(N__41443),
            .I(\PWM.n27 ));
    SRMux I__8455 (
            .O(N__41440),
            .I(N__41437));
    LocalMux I__8454 (
            .O(N__41437),
            .I(N__41433));
    SRMux I__8453 (
            .O(N__41436),
            .I(N__41430));
    Span4Mux_v I__8452 (
            .O(N__41433),
            .I(N__41424));
    LocalMux I__8451 (
            .O(N__41430),
            .I(N__41424));
    SRMux I__8450 (
            .O(N__41429),
            .I(N__41420));
    Span4Mux_s1_v I__8449 (
            .O(N__41424),
            .I(N__41417));
    SRMux I__8448 (
            .O(N__41423),
            .I(N__41414));
    LocalMux I__8447 (
            .O(N__41420),
            .I(N__41407));
    Span4Mux_h I__8446 (
            .O(N__41417),
            .I(N__41407));
    LocalMux I__8445 (
            .O(N__41414),
            .I(N__41407));
    Span4Mux_v I__8444 (
            .O(N__41407),
            .I(N__41404));
    Odrv4 I__8443 (
            .O(N__41404),
            .I(\PWM.pwm_counter_31__N_401 ));
    InMux I__8442 (
            .O(N__41401),
            .I(N__41396));
    InMux I__8441 (
            .O(N__41400),
            .I(N__41391));
    InMux I__8440 (
            .O(N__41399),
            .I(N__41391));
    LocalMux I__8439 (
            .O(N__41396),
            .I(pwm_counter_19));
    LocalMux I__8438 (
            .O(N__41391),
            .I(pwm_counter_19));
    InMux I__8437 (
            .O(N__41386),
            .I(N__41383));
    LocalMux I__8436 (
            .O(N__41383),
            .I(N__41380));
    Span4Mux_h I__8435 (
            .O(N__41380),
            .I(N__41377));
    Odrv4 I__8434 (
            .O(N__41377),
            .I(n39));
    InMux I__8433 (
            .O(N__41374),
            .I(N__41368));
    InMux I__8432 (
            .O(N__41373),
            .I(N__41368));
    LocalMux I__8431 (
            .O(N__41368),
            .I(pwm_setpoint_19));
    CascadeMux I__8430 (
            .O(N__41365),
            .I(n39_cascade_));
    InMux I__8429 (
            .O(N__41362),
            .I(N__41359));
    LocalMux I__8428 (
            .O(N__41359),
            .I(N__41356));
    Span4Mux_h I__8427 (
            .O(N__41356),
            .I(N__41353));
    Odrv4 I__8426 (
            .O(N__41353),
            .I(n14883));
    CascadeMux I__8425 (
            .O(N__41350),
            .I(N__41347));
    InMux I__8424 (
            .O(N__41347),
            .I(N__41344));
    LocalMux I__8423 (
            .O(N__41344),
            .I(N__41338));
    InMux I__8422 (
            .O(N__41343),
            .I(N__41335));
    InMux I__8421 (
            .O(N__41342),
            .I(N__41332));
    InMux I__8420 (
            .O(N__41341),
            .I(N__41329));
    Span4Mux_h I__8419 (
            .O(N__41338),
            .I(N__41324));
    LocalMux I__8418 (
            .O(N__41335),
            .I(N__41324));
    LocalMux I__8417 (
            .O(N__41332),
            .I(pwm_counter_9));
    LocalMux I__8416 (
            .O(N__41329),
            .I(pwm_counter_9));
    Odrv4 I__8415 (
            .O(N__41324),
            .I(pwm_counter_9));
    InMux I__8414 (
            .O(N__41317),
            .I(N__41314));
    LocalMux I__8413 (
            .O(N__41314),
            .I(N__41311));
    Odrv4 I__8412 (
            .O(N__41311),
            .I(n14804));
    CascadeMux I__8411 (
            .O(N__41308),
            .I(n19_adj_616_cascade_));
    InMux I__8410 (
            .O(N__41305),
            .I(N__41301));
    InMux I__8409 (
            .O(N__41304),
            .I(N__41298));
    LocalMux I__8408 (
            .O(N__41301),
            .I(n15_adj_613));
    LocalMux I__8407 (
            .O(N__41298),
            .I(n15_adj_613));
    InMux I__8406 (
            .O(N__41293),
            .I(N__41287));
    InMux I__8405 (
            .O(N__41292),
            .I(N__41287));
    LocalMux I__8404 (
            .O(N__41287),
            .I(pwm_setpoint_10));
    CascadeMux I__8403 (
            .O(N__41284),
            .I(n11_adj_610_cascade_));
    InMux I__8402 (
            .O(N__41281),
            .I(N__41275));
    InMux I__8401 (
            .O(N__41280),
            .I(N__41275));
    LocalMux I__8400 (
            .O(N__41275),
            .I(pwm_setpoint_5));
    InMux I__8399 (
            .O(N__41272),
            .I(N__41268));
    InMux I__8398 (
            .O(N__41271),
            .I(N__41265));
    LocalMux I__8397 (
            .O(N__41268),
            .I(N__41262));
    LocalMux I__8396 (
            .O(N__41265),
            .I(N__41259));
    Span4Mux_h I__8395 (
            .O(N__41262),
            .I(N__41256));
    Odrv4 I__8394 (
            .O(N__41259),
            .I(pwm_setpoint_6));
    Odrv4 I__8393 (
            .O(N__41256),
            .I(pwm_setpoint_6));
    SRMux I__8392 (
            .O(N__41251),
            .I(N__41248));
    LocalMux I__8391 (
            .O(N__41248),
            .I(N__41245));
    Span4Mux_h I__8390 (
            .O(N__41245),
            .I(N__41242));
    Span4Mux_s2_v I__8389 (
            .O(N__41242),
            .I(N__41239));
    Odrv4 I__8388 (
            .O(N__41239),
            .I(n4825));
    InMux I__8387 (
            .O(N__41236),
            .I(N__41230));
    InMux I__8386 (
            .O(N__41235),
            .I(N__41230));
    LocalMux I__8385 (
            .O(N__41230),
            .I(N__41227));
    Span4Mux_s3_v I__8384 (
            .O(N__41227),
            .I(N__41224));
    Odrv4 I__8383 (
            .O(N__41224),
            .I(n13_adj_612));
    CascadeMux I__8382 (
            .O(N__41221),
            .I(N__41218));
    InMux I__8381 (
            .O(N__41218),
            .I(N__41215));
    LocalMux I__8380 (
            .O(N__41215),
            .I(n11_adj_610));
    InMux I__8379 (
            .O(N__41212),
            .I(N__41209));
    LocalMux I__8378 (
            .O(N__41209),
            .I(N__41206));
    Odrv4 I__8377 (
            .O(N__41206),
            .I(n14745));
    InMux I__8376 (
            .O(N__41203),
            .I(N__41197));
    InMux I__8375 (
            .O(N__41202),
            .I(N__41197));
    LocalMux I__8374 (
            .O(N__41197),
            .I(N__41194));
    Odrv4 I__8373 (
            .O(N__41194),
            .I(pwm_setpoint_20));
    InMux I__8372 (
            .O(N__41191),
            .I(N__41187));
    InMux I__8371 (
            .O(N__41190),
            .I(N__41183));
    LocalMux I__8370 (
            .O(N__41187),
            .I(N__41180));
    InMux I__8369 (
            .O(N__41186),
            .I(N__41177));
    LocalMux I__8368 (
            .O(N__41183),
            .I(pwm_counter_5));
    Odrv4 I__8367 (
            .O(N__41180),
            .I(pwm_counter_5));
    LocalMux I__8366 (
            .O(N__41177),
            .I(pwm_counter_5));
    InMux I__8365 (
            .O(N__41170),
            .I(N__41166));
    InMux I__8364 (
            .O(N__41169),
            .I(N__41161));
    LocalMux I__8363 (
            .O(N__41166),
            .I(N__41158));
    InMux I__8362 (
            .O(N__41165),
            .I(N__41155));
    InMux I__8361 (
            .O(N__41164),
            .I(N__41152));
    LocalMux I__8360 (
            .O(N__41161),
            .I(pwm_counter_6));
    Odrv4 I__8359 (
            .O(N__41158),
            .I(pwm_counter_6));
    LocalMux I__8358 (
            .O(N__41155),
            .I(pwm_counter_6));
    LocalMux I__8357 (
            .O(N__41152),
            .I(pwm_counter_6));
    CascadeMux I__8356 (
            .O(N__41143),
            .I(N__41136));
    CascadeMux I__8355 (
            .O(N__41142),
            .I(N__41133));
    CascadeMux I__8354 (
            .O(N__41141),
            .I(N__41128));
    CascadeMux I__8353 (
            .O(N__41140),
            .I(N__41125));
    InMux I__8352 (
            .O(N__41139),
            .I(N__41121));
    InMux I__8351 (
            .O(N__41136),
            .I(N__41116));
    InMux I__8350 (
            .O(N__41133),
            .I(N__41116));
    InMux I__8349 (
            .O(N__41132),
            .I(N__41107));
    InMux I__8348 (
            .O(N__41131),
            .I(N__41107));
    InMux I__8347 (
            .O(N__41128),
            .I(N__41107));
    InMux I__8346 (
            .O(N__41125),
            .I(N__41107));
    InMux I__8345 (
            .O(N__41124),
            .I(N__41104));
    LocalMux I__8344 (
            .O(N__41121),
            .I(n4_adj_698));
    LocalMux I__8343 (
            .O(N__41116),
            .I(n4_adj_698));
    LocalMux I__8342 (
            .O(N__41107),
            .I(n4_adj_698));
    LocalMux I__8341 (
            .O(N__41104),
            .I(n4_adj_698));
    CascadeMux I__8340 (
            .O(N__41095),
            .I(N__41091));
    CascadeMux I__8339 (
            .O(N__41094),
            .I(N__41088));
    InMux I__8338 (
            .O(N__41091),
            .I(N__41085));
    InMux I__8337 (
            .O(N__41088),
            .I(N__41081));
    LocalMux I__8336 (
            .O(N__41085),
            .I(N__41078));
    InMux I__8335 (
            .O(N__41084),
            .I(N__41075));
    LocalMux I__8334 (
            .O(N__41081),
            .I(dti_counter_5));
    Odrv4 I__8333 (
            .O(N__41078),
            .I(dti_counter_5));
    LocalMux I__8332 (
            .O(N__41075),
            .I(dti_counter_5));
    InMux I__8331 (
            .O(N__41068),
            .I(N__41061));
    InMux I__8330 (
            .O(N__41067),
            .I(N__41061));
    InMux I__8329 (
            .O(N__41066),
            .I(N__41052));
    LocalMux I__8328 (
            .O(N__41061),
            .I(N__41049));
    InMux I__8327 (
            .O(N__41060),
            .I(N__41046));
    InMux I__8326 (
            .O(N__41059),
            .I(N__41035));
    InMux I__8325 (
            .O(N__41058),
            .I(N__41035));
    InMux I__8324 (
            .O(N__41057),
            .I(N__41035));
    InMux I__8323 (
            .O(N__41056),
            .I(N__41035));
    InMux I__8322 (
            .O(N__41055),
            .I(N__41035));
    LocalMux I__8321 (
            .O(N__41052),
            .I(commutation_state_prev_0));
    Odrv4 I__8320 (
            .O(N__41049),
            .I(commutation_state_prev_0));
    LocalMux I__8319 (
            .O(N__41046),
            .I(commutation_state_prev_0));
    LocalMux I__8318 (
            .O(N__41035),
            .I(commutation_state_prev_0));
    InMux I__8317 (
            .O(N__41026),
            .I(N__41023));
    LocalMux I__8316 (
            .O(N__41023),
            .I(n14689));
    InMux I__8315 (
            .O(N__41020),
            .I(N__41014));
    InMux I__8314 (
            .O(N__41019),
            .I(N__41014));
    LocalMux I__8313 (
            .O(N__41014),
            .I(pwm_setpoint_2));
    InMux I__8312 (
            .O(N__41011),
            .I(N__41008));
    LocalMux I__8311 (
            .O(N__41008),
            .I(N__41004));
    InMux I__8310 (
            .O(N__41007),
            .I(N__41001));
    Span4Mux_s3_v I__8309 (
            .O(N__41004),
            .I(N__40996));
    LocalMux I__8308 (
            .O(N__41001),
            .I(N__40996));
    Odrv4 I__8307 (
            .O(N__40996),
            .I(pwm_setpoint_11));
    InMux I__8306 (
            .O(N__40993),
            .I(N__40989));
    InMux I__8305 (
            .O(N__40992),
            .I(N__40986));
    LocalMux I__8304 (
            .O(N__40989),
            .I(N__40981));
    LocalMux I__8303 (
            .O(N__40986),
            .I(N__40981));
    Span4Mux_s3_v I__8302 (
            .O(N__40981),
            .I(N__40978));
    Odrv4 I__8301 (
            .O(N__40978),
            .I(pwm_setpoint_8));
    InMux I__8300 (
            .O(N__40975),
            .I(N__40970));
    InMux I__8299 (
            .O(N__40974),
            .I(N__40967));
    InMux I__8298 (
            .O(N__40973),
            .I(N__40964));
    LocalMux I__8297 (
            .O(N__40970),
            .I(pwm_counter_10));
    LocalMux I__8296 (
            .O(N__40967),
            .I(pwm_counter_10));
    LocalMux I__8295 (
            .O(N__40964),
            .I(pwm_counter_10));
    CascadeMux I__8294 (
            .O(N__40957),
            .I(n21_adj_617_cascade_));
    InMux I__8293 (
            .O(N__40954),
            .I(N__40951));
    LocalMux I__8292 (
            .O(N__40951),
            .I(n6_adj_606));
    InMux I__8291 (
            .O(N__40948),
            .I(N__40945));
    LocalMux I__8290 (
            .O(N__40945),
            .I(N__40942));
    Span4Mux_h I__8289 (
            .O(N__40942),
            .I(N__40939));
    Odrv4 I__8288 (
            .O(N__40939),
            .I(n14842));
    InMux I__8287 (
            .O(N__40936),
            .I(N__40933));
    LocalMux I__8286 (
            .O(N__40933),
            .I(N__40930));
    Odrv4 I__8285 (
            .O(N__40930),
            .I(n14690));
    CascadeMux I__8284 (
            .O(N__40927),
            .I(N__40922));
    InMux I__8283 (
            .O(N__40926),
            .I(N__40919));
    InMux I__8282 (
            .O(N__40925),
            .I(N__40916));
    InMux I__8281 (
            .O(N__40922),
            .I(N__40913));
    LocalMux I__8280 (
            .O(N__40919),
            .I(dti_counter_4));
    LocalMux I__8279 (
            .O(N__40916),
            .I(dti_counter_4));
    LocalMux I__8278 (
            .O(N__40913),
            .I(dti_counter_4));
    InMux I__8277 (
            .O(N__40906),
            .I(n12745));
    InMux I__8276 (
            .O(N__40903),
            .I(n12746));
    InMux I__8275 (
            .O(N__40900),
            .I(N__40897));
    LocalMux I__8274 (
            .O(N__40897),
            .I(n14688));
    InMux I__8273 (
            .O(N__40894),
            .I(N__40889));
    InMux I__8272 (
            .O(N__40893),
            .I(N__40884));
    InMux I__8271 (
            .O(N__40892),
            .I(N__40884));
    LocalMux I__8270 (
            .O(N__40889),
            .I(dti_counter_6));
    LocalMux I__8269 (
            .O(N__40884),
            .I(dti_counter_6));
    InMux I__8268 (
            .O(N__40879),
            .I(n12747));
    InMux I__8267 (
            .O(N__40876),
            .I(N__40873));
    LocalMux I__8266 (
            .O(N__40873),
            .I(n14687));
    CascadeMux I__8265 (
            .O(N__40870),
            .I(N__40864));
    CascadeMux I__8264 (
            .O(N__40869),
            .I(N__40860));
    CascadeMux I__8263 (
            .O(N__40868),
            .I(N__40856));
    InMux I__8262 (
            .O(N__40867),
            .I(N__40840));
    InMux I__8261 (
            .O(N__40864),
            .I(N__40840));
    InMux I__8260 (
            .O(N__40863),
            .I(N__40840));
    InMux I__8259 (
            .O(N__40860),
            .I(N__40840));
    InMux I__8258 (
            .O(N__40859),
            .I(N__40840));
    InMux I__8257 (
            .O(N__40856),
            .I(N__40840));
    InMux I__8256 (
            .O(N__40855),
            .I(N__40840));
    LocalMux I__8255 (
            .O(N__40840),
            .I(N__40837));
    Odrv4 I__8254 (
            .O(N__40837),
            .I(n11202));
    InMux I__8253 (
            .O(N__40834),
            .I(n12748));
    CascadeMux I__8252 (
            .O(N__40831),
            .I(N__40827));
    CascadeMux I__8251 (
            .O(N__40830),
            .I(N__40824));
    InMux I__8250 (
            .O(N__40827),
            .I(N__40821));
    InMux I__8249 (
            .O(N__40824),
            .I(N__40817));
    LocalMux I__8248 (
            .O(N__40821),
            .I(N__40814));
    InMux I__8247 (
            .O(N__40820),
            .I(N__40811));
    LocalMux I__8246 (
            .O(N__40817),
            .I(dti_counter_7));
    Odrv4 I__8245 (
            .O(N__40814),
            .I(dti_counter_7));
    LocalMux I__8244 (
            .O(N__40811),
            .I(dti_counter_7));
    InMux I__8243 (
            .O(N__40804),
            .I(N__40801));
    LocalMux I__8242 (
            .O(N__40801),
            .I(N__40798));
    Span4Mux_v I__8241 (
            .O(N__40798),
            .I(N__40794));
    InMux I__8240 (
            .O(N__40797),
            .I(N__40791));
    Odrv4 I__8239 (
            .O(N__40794),
            .I(pwm_setpoint_4));
    LocalMux I__8238 (
            .O(N__40791),
            .I(pwm_setpoint_4));
    CascadeMux I__8237 (
            .O(N__40786),
            .I(N__40783));
    InMux I__8236 (
            .O(N__40783),
            .I(N__40779));
    InMux I__8235 (
            .O(N__40782),
            .I(N__40776));
    LocalMux I__8234 (
            .O(N__40779),
            .I(N__40773));
    LocalMux I__8233 (
            .O(N__40776),
            .I(pwm_counter_2));
    Odrv4 I__8232 (
            .O(N__40773),
            .I(pwm_counter_2));
    InMux I__8231 (
            .O(N__40768),
            .I(N__40763));
    InMux I__8230 (
            .O(N__40767),
            .I(N__40758));
    InMux I__8229 (
            .O(N__40766),
            .I(N__40758));
    LocalMux I__8228 (
            .O(N__40763),
            .I(pwm_counter_3));
    LocalMux I__8227 (
            .O(N__40758),
            .I(pwm_counter_3));
    CascadeMux I__8226 (
            .O(N__40753),
            .I(N__40750));
    InMux I__8225 (
            .O(N__40750),
            .I(N__40744));
    InMux I__8224 (
            .O(N__40749),
            .I(N__40744));
    LocalMux I__8223 (
            .O(N__40744),
            .I(pwm_setpoint_3));
    CascadeMux I__8222 (
            .O(N__40741),
            .I(n14_adj_679_cascade_));
    CascadeMux I__8221 (
            .O(N__40738),
            .I(n4781_cascade_));
    InMux I__8220 (
            .O(N__40735),
            .I(N__40732));
    LocalMux I__8219 (
            .O(N__40732),
            .I(n14700));
    InMux I__8218 (
            .O(N__40729),
            .I(N__40726));
    LocalMux I__8217 (
            .O(N__40726),
            .I(n1259));
    CascadeMux I__8216 (
            .O(N__40723),
            .I(N__40719));
    InMux I__8215 (
            .O(N__40722),
            .I(N__40715));
    InMux I__8214 (
            .O(N__40719),
            .I(N__40712));
    InMux I__8213 (
            .O(N__40718),
            .I(N__40709));
    LocalMux I__8212 (
            .O(N__40715),
            .I(dti_counter_0));
    LocalMux I__8211 (
            .O(N__40712),
            .I(dti_counter_0));
    LocalMux I__8210 (
            .O(N__40709),
            .I(dti_counter_0));
    InMux I__8209 (
            .O(N__40702),
            .I(bfn_12_27_0_));
    InMux I__8208 (
            .O(N__40699),
            .I(N__40696));
    LocalMux I__8207 (
            .O(N__40696),
            .I(n14693));
    InMux I__8206 (
            .O(N__40693),
            .I(n12742));
    InMux I__8205 (
            .O(N__40690),
            .I(N__40687));
    LocalMux I__8204 (
            .O(N__40687),
            .I(n14692));
    InMux I__8203 (
            .O(N__40684),
            .I(n12743));
    InMux I__8202 (
            .O(N__40681),
            .I(N__40678));
    LocalMux I__8201 (
            .O(N__40678),
            .I(n14691));
    CascadeMux I__8200 (
            .O(N__40675),
            .I(N__40671));
    CascadeMux I__8199 (
            .O(N__40674),
            .I(N__40668));
    InMux I__8198 (
            .O(N__40671),
            .I(N__40665));
    InMux I__8197 (
            .O(N__40668),
            .I(N__40661));
    LocalMux I__8196 (
            .O(N__40665),
            .I(N__40658));
    InMux I__8195 (
            .O(N__40664),
            .I(N__40655));
    LocalMux I__8194 (
            .O(N__40661),
            .I(dti_counter_3));
    Odrv12 I__8193 (
            .O(N__40658),
            .I(dti_counter_3));
    LocalMux I__8192 (
            .O(N__40655),
            .I(dti_counter_3));
    InMux I__8191 (
            .O(N__40648),
            .I(n12744));
    CascadeMux I__8190 (
            .O(N__40645),
            .I(n13848_cascade_));
    InMux I__8189 (
            .O(N__40642),
            .I(N__40639));
    LocalMux I__8188 (
            .O(N__40639),
            .I(N__40636));
    Odrv4 I__8187 (
            .O(N__40636),
            .I(n5_adj_713));
    CascadeMux I__8186 (
            .O(N__40633),
            .I(n13850_cascade_));
    InMux I__8185 (
            .O(N__40630),
            .I(N__40627));
    LocalMux I__8184 (
            .O(N__40627),
            .I(N__40624));
    Odrv4 I__8183 (
            .O(N__40624),
            .I(n11656));
    CascadeMux I__8182 (
            .O(N__40621),
            .I(n13852_cascade_));
    InMux I__8181 (
            .O(N__40618),
            .I(N__40615));
    LocalMux I__8180 (
            .O(N__40615),
            .I(n13854));
    InMux I__8179 (
            .O(N__40612),
            .I(N__40609));
    LocalMux I__8178 (
            .O(N__40609),
            .I(n37_adj_710));
    InMux I__8177 (
            .O(N__40606),
            .I(N__40603));
    LocalMux I__8176 (
            .O(N__40603),
            .I(n7_adj_703));
    CascadeMux I__8175 (
            .O(N__40600),
            .I(n23_adj_707_cascade_));
    CascadeMux I__8174 (
            .O(N__40597),
            .I(n25_adj_708_cascade_));
    CascadeMux I__8173 (
            .O(N__40594),
            .I(n13832_cascade_));
    InMux I__8172 (
            .O(N__40591),
            .I(N__40588));
    LocalMux I__8171 (
            .O(N__40588),
            .I(n13828));
    InMux I__8170 (
            .O(N__40585),
            .I(N__40582));
    LocalMux I__8169 (
            .O(N__40582),
            .I(n13826));
    CascadeMux I__8168 (
            .O(N__40579),
            .I(n13840_cascade_));
    InMux I__8167 (
            .O(N__40576),
            .I(N__40573));
    LocalMux I__8166 (
            .O(N__40573),
            .I(n13846));
    InMux I__8165 (
            .O(N__40570),
            .I(N__40567));
    LocalMux I__8164 (
            .O(N__40567),
            .I(N__40564));
    Odrv4 I__8163 (
            .O(N__40564),
            .I(n13466));
    InMux I__8162 (
            .O(N__40561),
            .I(N__40558));
    LocalMux I__8161 (
            .O(N__40558),
            .I(n14334));
    CascadeMux I__8160 (
            .O(N__40555),
            .I(n3121_cascade_));
    CascadeMux I__8159 (
            .O(N__40552),
            .I(n3112_cascade_));
    CascadeMux I__8158 (
            .O(N__40549),
            .I(N__40546));
    InMux I__8157 (
            .O(N__40546),
            .I(N__40542));
    InMux I__8156 (
            .O(N__40545),
            .I(N__40539));
    LocalMux I__8155 (
            .O(N__40542),
            .I(N__40534));
    LocalMux I__8154 (
            .O(N__40539),
            .I(N__40534));
    Span4Mux_h I__8153 (
            .O(N__40534),
            .I(N__40530));
    InMux I__8152 (
            .O(N__40533),
            .I(N__40527));
    Odrv4 I__8151 (
            .O(N__40530),
            .I(n2911));
    LocalMux I__8150 (
            .O(N__40527),
            .I(n2911));
    CascadeMux I__8149 (
            .O(N__40522),
            .I(N__40519));
    InMux I__8148 (
            .O(N__40519),
            .I(N__40515));
    InMux I__8147 (
            .O(N__40518),
            .I(N__40512));
    LocalMux I__8146 (
            .O(N__40515),
            .I(n2912));
    LocalMux I__8145 (
            .O(N__40512),
            .I(n2912));
    CascadeMux I__8144 (
            .O(N__40507),
            .I(n13948_cascade_));
    CascadeMux I__8143 (
            .O(N__40504),
            .I(n13954_cascade_));
    InMux I__8142 (
            .O(N__40501),
            .I(N__40498));
    LocalMux I__8141 (
            .O(N__40498),
            .I(N__40495));
    Odrv4 I__8140 (
            .O(N__40495),
            .I(n2999));
    CascadeMux I__8139 (
            .O(N__40492),
            .I(n2940_cascade_));
    CascadeMux I__8138 (
            .O(N__40489),
            .I(N__40486));
    InMux I__8137 (
            .O(N__40486),
            .I(N__40483));
    LocalMux I__8136 (
            .O(N__40483),
            .I(N__40480));
    Odrv4 I__8135 (
            .O(N__40480),
            .I(n2996));
    CascadeMux I__8134 (
            .O(N__40477),
            .I(n14340_cascade_));
    InMux I__8133 (
            .O(N__40474),
            .I(N__40471));
    LocalMux I__8132 (
            .O(N__40471),
            .I(N__40467));
    InMux I__8131 (
            .O(N__40470),
            .I(N__40463));
    Span4Mux_v I__8130 (
            .O(N__40467),
            .I(N__40460));
    InMux I__8129 (
            .O(N__40466),
            .I(N__40457));
    LocalMux I__8128 (
            .O(N__40463),
            .I(n2908));
    Odrv4 I__8127 (
            .O(N__40460),
            .I(n2908));
    LocalMux I__8126 (
            .O(N__40457),
            .I(n2908));
    InMux I__8125 (
            .O(N__40450),
            .I(N__40447));
    LocalMux I__8124 (
            .O(N__40447),
            .I(n14344));
    CascadeMux I__8123 (
            .O(N__40444),
            .I(n3039_cascade_));
    InMux I__8122 (
            .O(N__40441),
            .I(N__40438));
    LocalMux I__8121 (
            .O(N__40438),
            .I(N__40435));
    Span4Mux_h I__8120 (
            .O(N__40435),
            .I(N__40432));
    Odrv4 I__8119 (
            .O(N__40432),
            .I(n2777));
    InMux I__8118 (
            .O(N__40429),
            .I(bfn_12_20_0_));
    InMux I__8117 (
            .O(N__40426),
            .I(n12410));
    InMux I__8116 (
            .O(N__40423),
            .I(N__40420));
    LocalMux I__8115 (
            .O(N__40420),
            .I(N__40417));
    Span4Mux_h I__8114 (
            .O(N__40417),
            .I(N__40414));
    Odrv4 I__8113 (
            .O(N__40414),
            .I(n2985));
    CascadeMux I__8112 (
            .O(N__40411),
            .I(n3017_cascade_));
    InMux I__8111 (
            .O(N__40408),
            .I(N__40405));
    LocalMux I__8110 (
            .O(N__40405),
            .I(N__40402));
    Span4Mux_v I__8109 (
            .O(N__40402),
            .I(N__40399));
    Odrv4 I__8108 (
            .O(N__40399),
            .I(n2977));
    CascadeMux I__8107 (
            .O(N__40396),
            .I(N__40393));
    InMux I__8106 (
            .O(N__40393),
            .I(N__40390));
    LocalMux I__8105 (
            .O(N__40390),
            .I(N__40387));
    Span4Mux_v I__8104 (
            .O(N__40387),
            .I(N__40384));
    Odrv4 I__8103 (
            .O(N__40384),
            .I(n2993));
    InMux I__8102 (
            .O(N__40381),
            .I(n12400));
    InMux I__8101 (
            .O(N__40378),
            .I(N__40374));
    InMux I__8100 (
            .O(N__40377),
            .I(N__40371));
    LocalMux I__8099 (
            .O(N__40374),
            .I(N__40366));
    LocalMux I__8098 (
            .O(N__40371),
            .I(N__40366));
    Span4Mux_h I__8097 (
            .O(N__40366),
            .I(N__40362));
    InMux I__8096 (
            .O(N__40365),
            .I(N__40359));
    Odrv4 I__8095 (
            .O(N__40362),
            .I(n2718));
    LocalMux I__8094 (
            .O(N__40359),
            .I(n2718));
    CascadeMux I__8093 (
            .O(N__40354),
            .I(N__40351));
    InMux I__8092 (
            .O(N__40351),
            .I(N__40348));
    LocalMux I__8091 (
            .O(N__40348),
            .I(n2785));
    InMux I__8090 (
            .O(N__40345),
            .I(bfn_12_19_0_));
    InMux I__8089 (
            .O(N__40342),
            .I(N__40337));
    InMux I__8088 (
            .O(N__40341),
            .I(N__40334));
    InMux I__8087 (
            .O(N__40340),
            .I(N__40331));
    LocalMux I__8086 (
            .O(N__40337),
            .I(N__40328));
    LocalMux I__8085 (
            .O(N__40334),
            .I(N__40325));
    LocalMux I__8084 (
            .O(N__40331),
            .I(n2717));
    Odrv4 I__8083 (
            .O(N__40328),
            .I(n2717));
    Odrv4 I__8082 (
            .O(N__40325),
            .I(n2717));
    CascadeMux I__8081 (
            .O(N__40318),
            .I(N__40315));
    InMux I__8080 (
            .O(N__40315),
            .I(N__40312));
    LocalMux I__8079 (
            .O(N__40312),
            .I(n2784));
    InMux I__8078 (
            .O(N__40309),
            .I(n12402));
    InMux I__8077 (
            .O(N__40306),
            .I(n12403));
    InMux I__8076 (
            .O(N__40303),
            .I(n12404));
    InMux I__8075 (
            .O(N__40300),
            .I(N__40297));
    LocalMux I__8074 (
            .O(N__40297),
            .I(n2781));
    InMux I__8073 (
            .O(N__40294),
            .I(n12405));
    InMux I__8072 (
            .O(N__40291),
            .I(n12406));
    InMux I__8071 (
            .O(N__40288),
            .I(n12407));
    InMux I__8070 (
            .O(N__40285),
            .I(n12408));
    InMux I__8069 (
            .O(N__40282),
            .I(n12391));
    InMux I__8068 (
            .O(N__40279),
            .I(n12392));
    InMux I__8067 (
            .O(N__40276),
            .I(bfn_12_18_0_));
    InMux I__8066 (
            .O(N__40273),
            .I(n12394));
    InMux I__8065 (
            .O(N__40270),
            .I(n12395));
    InMux I__8064 (
            .O(N__40267),
            .I(n12396));
    InMux I__8063 (
            .O(N__40264),
            .I(n12397));
    CascadeMux I__8062 (
            .O(N__40261),
            .I(N__40258));
    InMux I__8061 (
            .O(N__40258),
            .I(N__40255));
    LocalMux I__8060 (
            .O(N__40255),
            .I(N__40251));
    InMux I__8059 (
            .O(N__40254),
            .I(N__40248));
    Odrv4 I__8058 (
            .O(N__40251),
            .I(n2721));
    LocalMux I__8057 (
            .O(N__40248),
            .I(n2721));
    InMux I__8056 (
            .O(N__40243),
            .I(N__40240));
    LocalMux I__8055 (
            .O(N__40240),
            .I(N__40237));
    Odrv4 I__8054 (
            .O(N__40237),
            .I(n2788));
    InMux I__8053 (
            .O(N__40234),
            .I(n12398));
    InMux I__8052 (
            .O(N__40231),
            .I(n12399));
    InMux I__8051 (
            .O(N__40228),
            .I(N__40224));
    InMux I__8050 (
            .O(N__40227),
            .I(N__40221));
    LocalMux I__8049 (
            .O(N__40224),
            .I(pwm_counter_29));
    LocalMux I__8048 (
            .O(N__40221),
            .I(pwm_counter_29));
    InMux I__8047 (
            .O(N__40216),
            .I(\PWM.n12714 ));
    InMux I__8046 (
            .O(N__40213),
            .I(N__40209));
    InMux I__8045 (
            .O(N__40212),
            .I(N__40206));
    LocalMux I__8044 (
            .O(N__40209),
            .I(pwm_counter_30));
    LocalMux I__8043 (
            .O(N__40206),
            .I(pwm_counter_30));
    InMux I__8042 (
            .O(N__40201),
            .I(\PWM.n12715 ));
    InMux I__8041 (
            .O(N__40198),
            .I(\PWM.n12716 ));
    InMux I__8040 (
            .O(N__40195),
            .I(bfn_12_17_0_));
    InMux I__8039 (
            .O(N__40192),
            .I(n12386));
    InMux I__8038 (
            .O(N__40189),
            .I(n12387));
    InMux I__8037 (
            .O(N__40186),
            .I(n12388));
    InMux I__8036 (
            .O(N__40183),
            .I(n12389));
    InMux I__8035 (
            .O(N__40180),
            .I(n12390));
    InMux I__8034 (
            .O(N__40177),
            .I(N__40170));
    InMux I__8033 (
            .O(N__40176),
            .I(N__40170));
    InMux I__8032 (
            .O(N__40175),
            .I(N__40165));
    LocalMux I__8031 (
            .O(N__40170),
            .I(N__40162));
    InMux I__8030 (
            .O(N__40169),
            .I(N__40159));
    InMux I__8029 (
            .O(N__40168),
            .I(N__40156));
    LocalMux I__8028 (
            .O(N__40165),
            .I(N__40153));
    Span4Mux_h I__8027 (
            .O(N__40162),
            .I(N__40150));
    LocalMux I__8026 (
            .O(N__40159),
            .I(pwm_counter_21));
    LocalMux I__8025 (
            .O(N__40156),
            .I(pwm_counter_21));
    Odrv4 I__8024 (
            .O(N__40153),
            .I(pwm_counter_21));
    Odrv4 I__8023 (
            .O(N__40150),
            .I(pwm_counter_21));
    InMux I__8022 (
            .O(N__40141),
            .I(\PWM.n12706 ));
    InMux I__8021 (
            .O(N__40138),
            .I(N__40135));
    LocalMux I__8020 (
            .O(N__40135),
            .I(N__40131));
    InMux I__8019 (
            .O(N__40134),
            .I(N__40127));
    Span4Mux_h I__8018 (
            .O(N__40131),
            .I(N__40124));
    InMux I__8017 (
            .O(N__40130),
            .I(N__40121));
    LocalMux I__8016 (
            .O(N__40127),
            .I(pwm_counter_22));
    Odrv4 I__8015 (
            .O(N__40124),
            .I(pwm_counter_22));
    LocalMux I__8014 (
            .O(N__40121),
            .I(pwm_counter_22));
    InMux I__8013 (
            .O(N__40114),
            .I(\PWM.n12707 ));
    InMux I__8012 (
            .O(N__40111),
            .I(\PWM.n12708 ));
    InMux I__8011 (
            .O(N__40108),
            .I(N__40104));
    InMux I__8010 (
            .O(N__40107),
            .I(N__40101));
    LocalMux I__8009 (
            .O(N__40104),
            .I(pwm_counter_24));
    LocalMux I__8008 (
            .O(N__40101),
            .I(pwm_counter_24));
    InMux I__8007 (
            .O(N__40096),
            .I(bfn_11_32_0_));
    InMux I__8006 (
            .O(N__40093),
            .I(N__40089));
    InMux I__8005 (
            .O(N__40092),
            .I(N__40086));
    LocalMux I__8004 (
            .O(N__40089),
            .I(pwm_counter_25));
    LocalMux I__8003 (
            .O(N__40086),
            .I(pwm_counter_25));
    InMux I__8002 (
            .O(N__40081),
            .I(\PWM.n12710 ));
    InMux I__8001 (
            .O(N__40078),
            .I(N__40074));
    InMux I__8000 (
            .O(N__40077),
            .I(N__40071));
    LocalMux I__7999 (
            .O(N__40074),
            .I(pwm_counter_26));
    LocalMux I__7998 (
            .O(N__40071),
            .I(pwm_counter_26));
    InMux I__7997 (
            .O(N__40066),
            .I(\PWM.n12711 ));
    CascadeMux I__7996 (
            .O(N__40063),
            .I(N__40059));
    InMux I__7995 (
            .O(N__40062),
            .I(N__40056));
    InMux I__7994 (
            .O(N__40059),
            .I(N__40053));
    LocalMux I__7993 (
            .O(N__40056),
            .I(pwm_counter_27));
    LocalMux I__7992 (
            .O(N__40053),
            .I(pwm_counter_27));
    InMux I__7991 (
            .O(N__40048),
            .I(\PWM.n12712 ));
    InMux I__7990 (
            .O(N__40045),
            .I(N__40041));
    InMux I__7989 (
            .O(N__40044),
            .I(N__40038));
    LocalMux I__7988 (
            .O(N__40041),
            .I(pwm_counter_28));
    LocalMux I__7987 (
            .O(N__40038),
            .I(pwm_counter_28));
    InMux I__7986 (
            .O(N__40033),
            .I(\PWM.n12713 ));
    InMux I__7985 (
            .O(N__40030),
            .I(\PWM.n12697 ));
    InMux I__7984 (
            .O(N__40027),
            .I(\PWM.n12698 ));
    InMux I__7983 (
            .O(N__40024),
            .I(\PWM.n12699 ));
    InMux I__7982 (
            .O(N__40021),
            .I(\PWM.n12700 ));
    InMux I__7981 (
            .O(N__40018),
            .I(bfn_11_31_0_));
    InMux I__7980 (
            .O(N__40015),
            .I(\PWM.n12702 ));
    InMux I__7979 (
            .O(N__40012),
            .I(\PWM.n12703 ));
    InMux I__7978 (
            .O(N__40009),
            .I(\PWM.n12704 ));
    InMux I__7977 (
            .O(N__40006),
            .I(N__40001));
    InMux I__7976 (
            .O(N__40005),
            .I(N__39996));
    InMux I__7975 (
            .O(N__40004),
            .I(N__39996));
    LocalMux I__7974 (
            .O(N__40001),
            .I(pwm_counter_20));
    LocalMux I__7973 (
            .O(N__39996),
            .I(pwm_counter_20));
    InMux I__7972 (
            .O(N__39991),
            .I(\PWM.n12705 ));
    InMux I__7971 (
            .O(N__39988),
            .I(\PWM.n12688 ));
    InMux I__7970 (
            .O(N__39985),
            .I(N__39981));
    InMux I__7969 (
            .O(N__39984),
            .I(N__39978));
    LocalMux I__7968 (
            .O(N__39981),
            .I(pwm_counter_4));
    LocalMux I__7967 (
            .O(N__39978),
            .I(pwm_counter_4));
    InMux I__7966 (
            .O(N__39973),
            .I(\PWM.n12689 ));
    InMux I__7965 (
            .O(N__39970),
            .I(\PWM.n12690 ));
    InMux I__7964 (
            .O(N__39967),
            .I(\PWM.n12691 ));
    InMux I__7963 (
            .O(N__39964),
            .I(\PWM.n12692 ));
    InMux I__7962 (
            .O(N__39961),
            .I(bfn_11_30_0_));
    InMux I__7961 (
            .O(N__39958),
            .I(\PWM.n12694 ));
    InMux I__7960 (
            .O(N__39955),
            .I(\PWM.n12695 ));
    CascadeMux I__7959 (
            .O(N__39952),
            .I(N__39948));
    InMux I__7958 (
            .O(N__39951),
            .I(N__39944));
    InMux I__7957 (
            .O(N__39948),
            .I(N__39941));
    InMux I__7956 (
            .O(N__39947),
            .I(N__39938));
    LocalMux I__7955 (
            .O(N__39944),
            .I(pwm_counter_11));
    LocalMux I__7954 (
            .O(N__39941),
            .I(pwm_counter_11));
    LocalMux I__7953 (
            .O(N__39938),
            .I(pwm_counter_11));
    InMux I__7952 (
            .O(N__39931),
            .I(\PWM.n12696 ));
    InMux I__7951 (
            .O(N__39928),
            .I(N__39925));
    LocalMux I__7950 (
            .O(N__39925),
            .I(N__39922));
    Span4Mux_h I__7949 (
            .O(N__39922),
            .I(N__39919));
    Odrv4 I__7948 (
            .O(N__39919),
            .I(encoder0_position_scaled_14));
    InMux I__7947 (
            .O(N__39916),
            .I(N__39913));
    LocalMux I__7946 (
            .O(N__39913),
            .I(N__39910));
    Span4Mux_h I__7945 (
            .O(N__39910),
            .I(N__39907));
    Odrv4 I__7944 (
            .O(N__39907),
            .I(encoder0_position_scaled_16));
    InMux I__7943 (
            .O(N__39904),
            .I(N__39901));
    LocalMux I__7942 (
            .O(N__39901),
            .I(N__39898));
    Span4Mux_h I__7941 (
            .O(N__39898),
            .I(N__39895));
    Odrv4 I__7940 (
            .O(N__39895),
            .I(encoder0_position_scaled_18));
    InMux I__7939 (
            .O(N__39892),
            .I(N__39889));
    LocalMux I__7938 (
            .O(N__39889),
            .I(commutation_state_prev_2));
    InMux I__7937 (
            .O(N__39886),
            .I(bfn_11_29_0_));
    InMux I__7936 (
            .O(N__39883),
            .I(\PWM.n12686 ));
    InMux I__7935 (
            .O(N__39880),
            .I(\PWM.n12687 ));
    InMux I__7934 (
            .O(N__39877),
            .I(N__39874));
    LocalMux I__7933 (
            .O(N__39874),
            .I(N__39871));
    Span4Mux_v I__7932 (
            .O(N__39871),
            .I(N__39868));
    Odrv4 I__7931 (
            .O(N__39868),
            .I(encoder0_position_scaled_7));
    InMux I__7930 (
            .O(N__39865),
            .I(N__39862));
    LocalMux I__7929 (
            .O(N__39862),
            .I(N__39859));
    Span4Mux_v I__7928 (
            .O(N__39859),
            .I(N__39856));
    Odrv4 I__7927 (
            .O(N__39856),
            .I(encoder0_position_scaled_1));
    CascadeMux I__7926 (
            .O(N__39853),
            .I(n4_adj_698_cascade_));
    InMux I__7925 (
            .O(N__39850),
            .I(N__39845));
    InMux I__7924 (
            .O(N__39849),
            .I(N__39842));
    InMux I__7923 (
            .O(N__39848),
            .I(N__39839));
    LocalMux I__7922 (
            .O(N__39845),
            .I(N__39836));
    LocalMux I__7921 (
            .O(N__39842),
            .I(N__39833));
    LocalMux I__7920 (
            .O(N__39839),
            .I(N__39830));
    Span4Mux_s3_v I__7919 (
            .O(N__39836),
            .I(N__39827));
    Span4Mux_s2_v I__7918 (
            .O(N__39833),
            .I(N__39822));
    Span4Mux_h I__7917 (
            .O(N__39830),
            .I(N__39822));
    Odrv4 I__7916 (
            .O(N__39827),
            .I(pwm_setpoint_21));
    Odrv4 I__7915 (
            .O(N__39822),
            .I(pwm_setpoint_21));
    CascadeMux I__7914 (
            .O(N__39817),
            .I(n13856_cascade_));
    CascadeMux I__7913 (
            .O(N__39814),
            .I(n13858_cascade_));
    CascadeMux I__7912 (
            .O(N__39811),
            .I(n13860_cascade_));
    CascadeMux I__7911 (
            .O(N__39808),
            .I(n13862_cascade_));
    CascadeMux I__7910 (
            .O(N__39805),
            .I(n13864_cascade_));
    InMux I__7909 (
            .O(N__39802),
            .I(N__39799));
    LocalMux I__7908 (
            .O(N__39799),
            .I(n13866));
    InMux I__7907 (
            .O(N__39796),
            .I(N__39793));
    LocalMux I__7906 (
            .O(N__39793),
            .I(N__39790));
    Span4Mux_h I__7905 (
            .O(N__39790),
            .I(N__39787));
    Odrv4 I__7904 (
            .O(N__39787),
            .I(encoder0_position_scaled_5));
    InMux I__7903 (
            .O(N__39784),
            .I(N__39781));
    LocalMux I__7902 (
            .O(N__39781),
            .I(N__39778));
    Odrv4 I__7901 (
            .O(N__39778),
            .I(encoder0_position_scaled_8));
    InMux I__7900 (
            .O(N__39775),
            .I(N__39772));
    LocalMux I__7899 (
            .O(N__39772),
            .I(N__39769));
    Odrv4 I__7898 (
            .O(N__39769),
            .I(encoder0_position_scaled_11));
    CascadeMux I__7897 (
            .O(N__39766),
            .I(n3010_cascade_));
    InMux I__7896 (
            .O(N__39763),
            .I(N__39760));
    LocalMux I__7895 (
            .O(N__39760),
            .I(N__39757));
    Span4Mux_h I__7894 (
            .O(N__39757),
            .I(N__39753));
    InMux I__7893 (
            .O(N__39756),
            .I(N__39750));
    Odrv4 I__7892 (
            .O(N__39753),
            .I(n15090));
    LocalMux I__7891 (
            .O(N__39750),
            .I(n15090));
    CascadeMux I__7890 (
            .O(N__39745),
            .I(n14392_cascade_));
    InMux I__7889 (
            .O(N__39742),
            .I(N__39739));
    LocalMux I__7888 (
            .O(N__39739),
            .I(N__39736));
    Odrv4 I__7887 (
            .O(N__39736),
            .I(n13470));
    CascadeMux I__7886 (
            .O(N__39733),
            .I(n14380_cascade_));
    InMux I__7885 (
            .O(N__39730),
            .I(N__39727));
    LocalMux I__7884 (
            .O(N__39727),
            .I(n14386));
    InMux I__7883 (
            .O(N__39724),
            .I(N__39721));
    LocalMux I__7882 (
            .O(N__39721),
            .I(n14398));
    CascadeMux I__7881 (
            .O(N__39718),
            .I(n3237_cascade_));
    InMux I__7880 (
            .O(N__39715),
            .I(N__39712));
    LocalMux I__7879 (
            .O(N__39712),
            .I(n61));
    InMux I__7878 (
            .O(N__39709),
            .I(N__39706));
    LocalMux I__7877 (
            .O(N__39706),
            .I(n2981));
    InMux I__7876 (
            .O(N__39703),
            .I(N__39700));
    LocalMux I__7875 (
            .O(N__39700),
            .I(n2984));
    CascadeMux I__7874 (
            .O(N__39697),
            .I(n2912_cascade_));
    InMux I__7873 (
            .O(N__39694),
            .I(N__39691));
    LocalMux I__7872 (
            .O(N__39691),
            .I(n2979));
    CascadeMux I__7871 (
            .O(N__39688),
            .I(N__39685));
    InMux I__7870 (
            .O(N__39685),
            .I(N__39682));
    LocalMux I__7869 (
            .O(N__39682),
            .I(N__39679));
    Odrv4 I__7868 (
            .O(N__39679),
            .I(n2975));
    CascadeMux I__7867 (
            .O(N__39676),
            .I(N__39673));
    InMux I__7866 (
            .O(N__39673),
            .I(N__39670));
    LocalMux I__7865 (
            .O(N__39670),
            .I(n2980));
    CascadeMux I__7864 (
            .O(N__39667),
            .I(N__39664));
    InMux I__7863 (
            .O(N__39664),
            .I(N__39661));
    LocalMux I__7862 (
            .O(N__39661),
            .I(n2976));
    InMux I__7861 (
            .O(N__39658),
            .I(N__39655));
    LocalMux I__7860 (
            .O(N__39655),
            .I(n2978));
    InMux I__7859 (
            .O(N__39652),
            .I(N__39649));
    LocalMux I__7858 (
            .O(N__39649),
            .I(n2998));
    CascadeMux I__7857 (
            .O(N__39646),
            .I(n3115_cascade_));
    InMux I__7856 (
            .O(N__39643),
            .I(N__39640));
    LocalMux I__7855 (
            .O(N__39640),
            .I(n13894));
    InMux I__7854 (
            .O(N__39637),
            .I(N__39634));
    LocalMux I__7853 (
            .O(N__39634),
            .I(N__39631));
    Span4Mux_v I__7852 (
            .O(N__39631),
            .I(N__39628));
    Odrv4 I__7851 (
            .O(N__39628),
            .I(n13898));
    InMux I__7850 (
            .O(N__39625),
            .I(N__39622));
    LocalMux I__7849 (
            .O(N__39622),
            .I(n2988));
    InMux I__7848 (
            .O(N__39619),
            .I(N__39616));
    LocalMux I__7847 (
            .O(N__39616),
            .I(n2987));
    CascadeMux I__7846 (
            .O(N__39613),
            .I(n3019_cascade_));
    CascadeMux I__7845 (
            .O(N__39610),
            .I(N__39607));
    InMux I__7844 (
            .O(N__39607),
            .I(N__39604));
    LocalMux I__7843 (
            .O(N__39604),
            .I(n2983));
    CascadeMux I__7842 (
            .O(N__39601),
            .I(n2817_cascade_));
    InMux I__7841 (
            .O(N__39598),
            .I(N__39595));
    LocalMux I__7840 (
            .O(N__39595),
            .I(n3000));
    CascadeMux I__7839 (
            .O(N__39592),
            .I(n3032_cascade_));
    CascadeMux I__7838 (
            .O(N__39589),
            .I(n11660_cascade_));
    CascadeMux I__7837 (
            .O(N__39586),
            .I(N__39583));
    InMux I__7836 (
            .O(N__39583),
            .I(N__39580));
    LocalMux I__7835 (
            .O(N__39580),
            .I(N__39577));
    Odrv4 I__7834 (
            .O(N__39577),
            .I(n2986));
    InMux I__7833 (
            .O(N__39574),
            .I(N__39571));
    LocalMux I__7832 (
            .O(N__39571),
            .I(n2997));
    CascadeMux I__7831 (
            .O(N__39568),
            .I(n3029_cascade_));
    InMux I__7830 (
            .O(N__39565),
            .I(N__39559));
    InMux I__7829 (
            .O(N__39564),
            .I(N__39551));
    InMux I__7828 (
            .O(N__39563),
            .I(N__39551));
    InMux I__7827 (
            .O(N__39562),
            .I(N__39551));
    LocalMux I__7826 (
            .O(N__39559),
            .I(N__39543));
    InMux I__7825 (
            .O(N__39558),
            .I(N__39539));
    LocalMux I__7824 (
            .O(N__39551),
            .I(N__39536));
    InMux I__7823 (
            .O(N__39550),
            .I(N__39519));
    InMux I__7822 (
            .O(N__39549),
            .I(N__39519));
    InMux I__7821 (
            .O(N__39548),
            .I(N__39519));
    InMux I__7820 (
            .O(N__39547),
            .I(N__39519));
    InMux I__7819 (
            .O(N__39546),
            .I(N__39513));
    Span4Mux_h I__7818 (
            .O(N__39543),
            .I(N__39510));
    InMux I__7817 (
            .O(N__39542),
            .I(N__39507));
    LocalMux I__7816 (
            .O(N__39539),
            .I(N__39504));
    Span4Mux_v I__7815 (
            .O(N__39536),
            .I(N__39501));
    InMux I__7814 (
            .O(N__39535),
            .I(N__39498));
    InMux I__7813 (
            .O(N__39534),
            .I(N__39493));
    InMux I__7812 (
            .O(N__39533),
            .I(N__39490));
    InMux I__7811 (
            .O(N__39532),
            .I(N__39487));
    CascadeMux I__7810 (
            .O(N__39531),
            .I(N__39482));
    CascadeMux I__7809 (
            .O(N__39530),
            .I(N__39477));
    CascadeMux I__7808 (
            .O(N__39529),
            .I(N__39472));
    CascadeMux I__7807 (
            .O(N__39528),
            .I(N__39468));
    LocalMux I__7806 (
            .O(N__39519),
            .I(N__39462));
    InMux I__7805 (
            .O(N__39518),
            .I(N__39455));
    InMux I__7804 (
            .O(N__39517),
            .I(N__39455));
    InMux I__7803 (
            .O(N__39516),
            .I(N__39455));
    LocalMux I__7802 (
            .O(N__39513),
            .I(N__39452));
    Span4Mux_v I__7801 (
            .O(N__39510),
            .I(N__39449));
    LocalMux I__7800 (
            .O(N__39507),
            .I(N__39446));
    Span4Mux_v I__7799 (
            .O(N__39504),
            .I(N__39437));
    Span4Mux_v I__7798 (
            .O(N__39501),
            .I(N__39437));
    LocalMux I__7797 (
            .O(N__39498),
            .I(N__39434));
    InMux I__7796 (
            .O(N__39497),
            .I(N__39429));
    InMux I__7795 (
            .O(N__39496),
            .I(N__39429));
    LocalMux I__7794 (
            .O(N__39493),
            .I(N__39422));
    LocalMux I__7793 (
            .O(N__39490),
            .I(N__39422));
    LocalMux I__7792 (
            .O(N__39487),
            .I(N__39422));
    InMux I__7791 (
            .O(N__39486),
            .I(N__39419));
    InMux I__7790 (
            .O(N__39485),
            .I(N__39408));
    InMux I__7789 (
            .O(N__39482),
            .I(N__39408));
    InMux I__7788 (
            .O(N__39481),
            .I(N__39408));
    InMux I__7787 (
            .O(N__39480),
            .I(N__39408));
    InMux I__7786 (
            .O(N__39477),
            .I(N__39408));
    InMux I__7785 (
            .O(N__39476),
            .I(N__39397));
    InMux I__7784 (
            .O(N__39475),
            .I(N__39397));
    InMux I__7783 (
            .O(N__39472),
            .I(N__39397));
    InMux I__7782 (
            .O(N__39471),
            .I(N__39397));
    InMux I__7781 (
            .O(N__39468),
            .I(N__39397));
    InMux I__7780 (
            .O(N__39467),
            .I(N__39391));
    InMux I__7779 (
            .O(N__39466),
            .I(N__39386));
    InMux I__7778 (
            .O(N__39465),
            .I(N__39386));
    Span4Mux_v I__7777 (
            .O(N__39462),
            .I(N__39379));
    LocalMux I__7776 (
            .O(N__39455),
            .I(N__39379));
    Span4Mux_h I__7775 (
            .O(N__39452),
            .I(N__39379));
    Span4Mux_h I__7774 (
            .O(N__39449),
            .I(N__39374));
    Span4Mux_h I__7773 (
            .O(N__39446),
            .I(N__39374));
    InMux I__7772 (
            .O(N__39445),
            .I(N__39367));
    InMux I__7771 (
            .O(N__39444),
            .I(N__39367));
    InMux I__7770 (
            .O(N__39443),
            .I(N__39367));
    InMux I__7769 (
            .O(N__39442),
            .I(N__39364));
    Span4Mux_h I__7768 (
            .O(N__39437),
            .I(N__39349));
    Span4Mux_h I__7767 (
            .O(N__39434),
            .I(N__39349));
    LocalMux I__7766 (
            .O(N__39429),
            .I(N__39349));
    Span4Mux_s3_v I__7765 (
            .O(N__39422),
            .I(N__39349));
    LocalMux I__7764 (
            .O(N__39419),
            .I(N__39349));
    LocalMux I__7763 (
            .O(N__39408),
            .I(N__39349));
    LocalMux I__7762 (
            .O(N__39397),
            .I(N__39349));
    InMux I__7761 (
            .O(N__39396),
            .I(N__39342));
    InMux I__7760 (
            .O(N__39395),
            .I(N__39342));
    InMux I__7759 (
            .O(N__39394),
            .I(N__39342));
    LocalMux I__7758 (
            .O(N__39391),
            .I(encoder0_position_31));
    LocalMux I__7757 (
            .O(N__39386),
            .I(encoder0_position_31));
    Odrv4 I__7756 (
            .O(N__39379),
            .I(encoder0_position_31));
    Odrv4 I__7755 (
            .O(N__39374),
            .I(encoder0_position_31));
    LocalMux I__7754 (
            .O(N__39367),
            .I(encoder0_position_31));
    LocalMux I__7753 (
            .O(N__39364),
            .I(encoder0_position_31));
    Odrv4 I__7752 (
            .O(N__39349),
            .I(encoder0_position_31));
    LocalMux I__7751 (
            .O(N__39342),
            .I(encoder0_position_31));
    InMux I__7750 (
            .O(N__39325),
            .I(N__39322));
    LocalMux I__7749 (
            .O(N__39322),
            .I(N__39319));
    Span12Mux_v I__7748 (
            .O(N__39319),
            .I(N__39316));
    Odrv12 I__7747 (
            .O(N__39316),
            .I(n29));
    InMux I__7746 (
            .O(N__39313),
            .I(N__39310));
    LocalMux I__7745 (
            .O(N__39310),
            .I(N__39306));
    CascadeMux I__7744 (
            .O(N__39309),
            .I(N__39303));
    Span4Mux_v I__7743 (
            .O(N__39306),
            .I(N__39299));
    InMux I__7742 (
            .O(N__39303),
            .I(N__39296));
    InMux I__7741 (
            .O(N__39302),
            .I(N__39293));
    Span4Mux_h I__7740 (
            .O(N__39299),
            .I(N__39290));
    LocalMux I__7739 (
            .O(N__39296),
            .I(N__39287));
    LocalMux I__7738 (
            .O(N__39293),
            .I(encoder0_position_4));
    Odrv4 I__7737 (
            .O(N__39290),
            .I(encoder0_position_4));
    Odrv4 I__7736 (
            .O(N__39287),
            .I(encoder0_position_4));
    InMux I__7735 (
            .O(N__39280),
            .I(N__39277));
    LocalMux I__7734 (
            .O(N__39277),
            .I(n3001));
    CascadeMux I__7733 (
            .O(N__39274),
            .I(n315_cascade_));
    CascadeMux I__7732 (
            .O(N__39271),
            .I(n2714_cascade_));
    CascadeMux I__7731 (
            .O(N__39268),
            .I(N__39265));
    InMux I__7730 (
            .O(N__39265),
            .I(N__39261));
    InMux I__7729 (
            .O(N__39264),
            .I(N__39258));
    LocalMux I__7728 (
            .O(N__39261),
            .I(N__39255));
    LocalMux I__7727 (
            .O(N__39258),
            .I(N__39251));
    Span4Mux_h I__7726 (
            .O(N__39255),
            .I(N__39248));
    InMux I__7725 (
            .O(N__39254),
            .I(N__39245));
    Odrv12 I__7724 (
            .O(N__39251),
            .I(n2623));
    Odrv4 I__7723 (
            .O(N__39248),
            .I(n2623));
    LocalMux I__7722 (
            .O(N__39245),
            .I(n2623));
    CascadeMux I__7721 (
            .O(N__39238),
            .I(N__39235));
    InMux I__7720 (
            .O(N__39235),
            .I(N__39232));
    LocalMux I__7719 (
            .O(N__39232),
            .I(N__39229));
    Span4Mux_v I__7718 (
            .O(N__39229),
            .I(N__39226));
    Odrv4 I__7717 (
            .O(N__39226),
            .I(n2690));
    InMux I__7716 (
            .O(N__39223),
            .I(N__39220));
    LocalMux I__7715 (
            .O(N__39220),
            .I(N__39217));
    Span4Mux_h I__7714 (
            .O(N__39217),
            .I(N__39214));
    Odrv4 I__7713 (
            .O(N__39214),
            .I(n2698));
    CascadeMux I__7712 (
            .O(N__39211),
            .I(N__39208));
    InMux I__7711 (
            .O(N__39208),
            .I(N__39205));
    LocalMux I__7710 (
            .O(N__39205),
            .I(N__39202));
    Span4Mux_h I__7709 (
            .O(N__39202),
            .I(N__39199));
    Odrv4 I__7708 (
            .O(N__39199),
            .I(n2699));
    CascadeMux I__7707 (
            .O(N__39196),
            .I(N__39192));
    InMux I__7706 (
            .O(N__39195),
            .I(N__39189));
    InMux I__7705 (
            .O(N__39192),
            .I(N__39186));
    LocalMux I__7704 (
            .O(N__39189),
            .I(N__39183));
    LocalMux I__7703 (
            .O(N__39186),
            .I(N__39180));
    Span4Mux_h I__7702 (
            .O(N__39183),
            .I(N__39174));
    Span4Mux_v I__7701 (
            .O(N__39180),
            .I(N__39174));
    InMux I__7700 (
            .O(N__39179),
            .I(N__39171));
    Odrv4 I__7699 (
            .O(N__39174),
            .I(n2217));
    LocalMux I__7698 (
            .O(N__39171),
            .I(n2217));
    CascadeMux I__7697 (
            .O(N__39166),
            .I(N__39163));
    InMux I__7696 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__7695 (
            .O(N__39160),
            .I(N__39157));
    Span4Mux_h I__7694 (
            .O(N__39157),
            .I(N__39154));
    Odrv4 I__7693 (
            .O(N__39154),
            .I(n2284));
    InMux I__7692 (
            .O(N__39151),
            .I(N__39146));
    CascadeMux I__7691 (
            .O(N__39150),
            .I(N__39140));
    InMux I__7690 (
            .O(N__39149),
            .I(N__39135));
    LocalMux I__7689 (
            .O(N__39146),
            .I(N__39129));
    InMux I__7688 (
            .O(N__39145),
            .I(N__39126));
    CascadeMux I__7687 (
            .O(N__39144),
            .I(N__39123));
    CascadeMux I__7686 (
            .O(N__39143),
            .I(N__39120));
    InMux I__7685 (
            .O(N__39140),
            .I(N__39112));
    InMux I__7684 (
            .O(N__39139),
            .I(N__39112));
    InMux I__7683 (
            .O(N__39138),
            .I(N__39112));
    LocalMux I__7682 (
            .O(N__39135),
            .I(N__39109));
    InMux I__7681 (
            .O(N__39134),
            .I(N__39106));
    InMux I__7680 (
            .O(N__39133),
            .I(N__39099));
    InMux I__7679 (
            .O(N__39132),
            .I(N__39099));
    Span4Mux_h I__7678 (
            .O(N__39129),
            .I(N__39092));
    LocalMux I__7677 (
            .O(N__39126),
            .I(N__39089));
    InMux I__7676 (
            .O(N__39123),
            .I(N__39082));
    InMux I__7675 (
            .O(N__39120),
            .I(N__39082));
    InMux I__7674 (
            .O(N__39119),
            .I(N__39082));
    LocalMux I__7673 (
            .O(N__39112),
            .I(N__39079));
    Span4Mux_h I__7672 (
            .O(N__39109),
            .I(N__39076));
    LocalMux I__7671 (
            .O(N__39106),
            .I(N__39073));
    CascadeMux I__7670 (
            .O(N__39105),
            .I(N__39068));
    InMux I__7669 (
            .O(N__39104),
            .I(N__39064));
    LocalMux I__7668 (
            .O(N__39099),
            .I(N__39061));
    InMux I__7667 (
            .O(N__39098),
            .I(N__39056));
    InMux I__7666 (
            .O(N__39097),
            .I(N__39056));
    InMux I__7665 (
            .O(N__39096),
            .I(N__39051));
    InMux I__7664 (
            .O(N__39095),
            .I(N__39051));
    Span4Mux_v I__7663 (
            .O(N__39092),
            .I(N__39042));
    Span4Mux_h I__7662 (
            .O(N__39089),
            .I(N__39042));
    LocalMux I__7661 (
            .O(N__39082),
            .I(N__39042));
    Span4Mux_h I__7660 (
            .O(N__39079),
            .I(N__39042));
    Span4Mux_h I__7659 (
            .O(N__39076),
            .I(N__39037));
    Span4Mux_h I__7658 (
            .O(N__39073),
            .I(N__39037));
    InMux I__7657 (
            .O(N__39072),
            .I(N__39028));
    InMux I__7656 (
            .O(N__39071),
            .I(N__39028));
    InMux I__7655 (
            .O(N__39068),
            .I(N__39028));
    InMux I__7654 (
            .O(N__39067),
            .I(N__39028));
    LocalMux I__7653 (
            .O(N__39064),
            .I(n2247));
    Odrv4 I__7652 (
            .O(N__39061),
            .I(n2247));
    LocalMux I__7651 (
            .O(N__39056),
            .I(n2247));
    LocalMux I__7650 (
            .O(N__39051),
            .I(n2247));
    Odrv4 I__7649 (
            .O(N__39042),
            .I(n2247));
    Odrv4 I__7648 (
            .O(N__39037),
            .I(n2247));
    LocalMux I__7647 (
            .O(N__39028),
            .I(n2247));
    InMux I__7646 (
            .O(N__39013),
            .I(N__39008));
    InMux I__7645 (
            .O(N__39012),
            .I(N__39005));
    InMux I__7644 (
            .O(N__39011),
            .I(N__39002));
    LocalMux I__7643 (
            .O(N__39008),
            .I(N__38995));
    LocalMux I__7642 (
            .O(N__39005),
            .I(N__38995));
    LocalMux I__7641 (
            .O(N__39002),
            .I(N__38995));
    Span12Mux_s6_h I__7640 (
            .O(N__38995),
            .I(N__38992));
    Odrv12 I__7639 (
            .O(N__38992),
            .I(n2316));
    InMux I__7638 (
            .O(N__38989),
            .I(N__38986));
    LocalMux I__7637 (
            .O(N__38986),
            .I(N__38982));
    InMux I__7636 (
            .O(N__38985),
            .I(N__38979));
    Span4Mux_h I__7635 (
            .O(N__38982),
            .I(N__38976));
    LocalMux I__7634 (
            .O(N__38979),
            .I(N__38973));
    Span4Mux_h I__7633 (
            .O(N__38976),
            .I(N__38970));
    Span4Mux_v I__7632 (
            .O(N__38973),
            .I(N__38967));
    Odrv4 I__7631 (
            .O(N__38970),
            .I(n2533));
    Odrv4 I__7630 (
            .O(N__38967),
            .I(n2533));
    CascadeMux I__7629 (
            .O(N__38962),
            .I(N__38959));
    InMux I__7628 (
            .O(N__38959),
            .I(N__38956));
    LocalMux I__7627 (
            .O(N__38956),
            .I(N__38953));
    Span4Mux_v I__7626 (
            .O(N__38953),
            .I(N__38950));
    Span4Mux_h I__7625 (
            .O(N__38950),
            .I(N__38947));
    Odrv4 I__7624 (
            .O(N__38947),
            .I(n2600));
    InMux I__7623 (
            .O(N__38944),
            .I(N__38940));
    CascadeMux I__7622 (
            .O(N__38943),
            .I(N__38937));
    LocalMux I__7621 (
            .O(N__38940),
            .I(N__38927));
    InMux I__7620 (
            .O(N__38937),
            .I(N__38924));
    InMux I__7619 (
            .O(N__38936),
            .I(N__38919));
    InMux I__7618 (
            .O(N__38935),
            .I(N__38919));
    InMux I__7617 (
            .O(N__38934),
            .I(N__38916));
    CascadeMux I__7616 (
            .O(N__38933),
            .I(N__38913));
    CascadeMux I__7615 (
            .O(N__38932),
            .I(N__38910));
    InMux I__7614 (
            .O(N__38931),
            .I(N__38904));
    CascadeMux I__7613 (
            .O(N__38930),
            .I(N__38901));
    Span4Mux_v I__7612 (
            .O(N__38927),
            .I(N__38894));
    LocalMux I__7611 (
            .O(N__38924),
            .I(N__38891));
    LocalMux I__7610 (
            .O(N__38919),
            .I(N__38888));
    LocalMux I__7609 (
            .O(N__38916),
            .I(N__38885));
    InMux I__7608 (
            .O(N__38913),
            .I(N__38874));
    InMux I__7607 (
            .O(N__38910),
            .I(N__38874));
    InMux I__7606 (
            .O(N__38909),
            .I(N__38874));
    InMux I__7605 (
            .O(N__38908),
            .I(N__38874));
    InMux I__7604 (
            .O(N__38907),
            .I(N__38874));
    LocalMux I__7603 (
            .O(N__38904),
            .I(N__38871));
    InMux I__7602 (
            .O(N__38901),
            .I(N__38863));
    InMux I__7601 (
            .O(N__38900),
            .I(N__38863));
    CascadeMux I__7600 (
            .O(N__38899),
            .I(N__38857));
    CascadeMux I__7599 (
            .O(N__38898),
            .I(N__38854));
    CascadeMux I__7598 (
            .O(N__38897),
            .I(N__38851));
    Span4Mux_v I__7597 (
            .O(N__38894),
            .I(N__38838));
    Span4Mux_v I__7596 (
            .O(N__38891),
            .I(N__38838));
    Span4Mux_v I__7595 (
            .O(N__38888),
            .I(N__38838));
    Span4Mux_h I__7594 (
            .O(N__38885),
            .I(N__38838));
    LocalMux I__7593 (
            .O(N__38874),
            .I(N__38838));
    Span4Mux_h I__7592 (
            .O(N__38871),
            .I(N__38835));
    InMux I__7591 (
            .O(N__38870),
            .I(N__38828));
    InMux I__7590 (
            .O(N__38869),
            .I(N__38828));
    InMux I__7589 (
            .O(N__38868),
            .I(N__38828));
    LocalMux I__7588 (
            .O(N__38863),
            .I(N__38825));
    InMux I__7587 (
            .O(N__38862),
            .I(N__38820));
    InMux I__7586 (
            .O(N__38861),
            .I(N__38820));
    InMux I__7585 (
            .O(N__38860),
            .I(N__38807));
    InMux I__7584 (
            .O(N__38857),
            .I(N__38807));
    InMux I__7583 (
            .O(N__38854),
            .I(N__38807));
    InMux I__7582 (
            .O(N__38851),
            .I(N__38807));
    InMux I__7581 (
            .O(N__38850),
            .I(N__38807));
    InMux I__7580 (
            .O(N__38849),
            .I(N__38807));
    Odrv4 I__7579 (
            .O(N__38838),
            .I(n2544));
    Odrv4 I__7578 (
            .O(N__38835),
            .I(n2544));
    LocalMux I__7577 (
            .O(N__38828),
            .I(n2544));
    Odrv4 I__7576 (
            .O(N__38825),
            .I(n2544));
    LocalMux I__7575 (
            .O(N__38820),
            .I(n2544));
    LocalMux I__7574 (
            .O(N__38807),
            .I(n2544));
    CascadeMux I__7573 (
            .O(N__38794),
            .I(N__38791));
    InMux I__7572 (
            .O(N__38791),
            .I(N__38787));
    InMux I__7571 (
            .O(N__38790),
            .I(N__38784));
    LocalMux I__7570 (
            .O(N__38787),
            .I(N__38781));
    LocalMux I__7569 (
            .O(N__38784),
            .I(n2632));
    Odrv4 I__7568 (
            .O(N__38781),
            .I(n2632));
    InMux I__7567 (
            .O(N__38776),
            .I(N__38771));
    InMux I__7566 (
            .O(N__38775),
            .I(N__38768));
    InMux I__7565 (
            .O(N__38774),
            .I(N__38765));
    LocalMux I__7564 (
            .O(N__38771),
            .I(N__38762));
    LocalMux I__7563 (
            .O(N__38768),
            .I(N__38759));
    LocalMux I__7562 (
            .O(N__38765),
            .I(N__38756));
    Span4Mux_v I__7561 (
            .O(N__38762),
            .I(N__38753));
    Span4Mux_h I__7560 (
            .O(N__38759),
            .I(N__38748));
    Span4Mux_h I__7559 (
            .O(N__38756),
            .I(N__38748));
    Span4Mux_v I__7558 (
            .O(N__38753),
            .I(N__38745));
    Span4Mux_v I__7557 (
            .O(N__38748),
            .I(N__38742));
    Odrv4 I__7556 (
            .O(N__38745),
            .I(n312));
    Odrv4 I__7555 (
            .O(N__38742),
            .I(n312));
    InMux I__7554 (
            .O(N__38737),
            .I(N__38733));
    CascadeMux I__7553 (
            .O(N__38736),
            .I(N__38730));
    LocalMux I__7552 (
            .O(N__38733),
            .I(N__38726));
    InMux I__7551 (
            .O(N__38730),
            .I(N__38723));
    InMux I__7550 (
            .O(N__38729),
            .I(N__38720));
    Span4Mux_h I__7549 (
            .O(N__38726),
            .I(N__38717));
    LocalMux I__7548 (
            .O(N__38723),
            .I(N__38712));
    LocalMux I__7547 (
            .O(N__38720),
            .I(N__38712));
    Odrv4 I__7546 (
            .O(N__38717),
            .I(n2633));
    Odrv12 I__7545 (
            .O(N__38712),
            .I(n2633));
    CascadeMux I__7544 (
            .O(N__38707),
            .I(n2632_cascade_));
    InMux I__7543 (
            .O(N__38704),
            .I(N__38700));
    CascadeMux I__7542 (
            .O(N__38703),
            .I(N__38697));
    LocalMux I__7541 (
            .O(N__38700),
            .I(N__38693));
    InMux I__7540 (
            .O(N__38697),
            .I(N__38690));
    InMux I__7539 (
            .O(N__38696),
            .I(N__38687));
    Span4Mux_h I__7538 (
            .O(N__38693),
            .I(N__38684));
    LocalMux I__7537 (
            .O(N__38690),
            .I(N__38679));
    LocalMux I__7536 (
            .O(N__38687),
            .I(N__38679));
    Odrv4 I__7535 (
            .O(N__38684),
            .I(n2631));
    Odrv12 I__7534 (
            .O(N__38679),
            .I(n2631));
    InMux I__7533 (
            .O(N__38674),
            .I(N__38671));
    LocalMux I__7532 (
            .O(N__38671),
            .I(N__38668));
    Span4Mux_v I__7531 (
            .O(N__38668),
            .I(N__38665));
    Odrv4 I__7530 (
            .O(N__38665),
            .I(n11760));
    CascadeMux I__7529 (
            .O(N__38662),
            .I(n2732_cascade_));
    CascadeMux I__7528 (
            .O(N__38659),
            .I(n11666_cascade_));
    InMux I__7527 (
            .O(N__38656),
            .I(N__38653));
    LocalMux I__7526 (
            .O(N__38653),
            .I(N__38650));
    Span4Mux_h I__7525 (
            .O(N__38650),
            .I(N__38647));
    Odrv4 I__7524 (
            .O(N__38647),
            .I(n2691));
    CascadeMux I__7523 (
            .O(N__38644),
            .I(N__38640));
    CascadeMux I__7522 (
            .O(N__38643),
            .I(N__38637));
    InMux I__7521 (
            .O(N__38640),
            .I(N__38634));
    InMux I__7520 (
            .O(N__38637),
            .I(N__38631));
    LocalMux I__7519 (
            .O(N__38634),
            .I(N__38628));
    LocalMux I__7518 (
            .O(N__38631),
            .I(N__38625));
    Span4Mux_h I__7517 (
            .O(N__38628),
            .I(N__38619));
    Span4Mux_v I__7516 (
            .O(N__38625),
            .I(N__38619));
    InMux I__7515 (
            .O(N__38624),
            .I(N__38616));
    Odrv4 I__7514 (
            .O(N__38619),
            .I(n2624));
    LocalMux I__7513 (
            .O(N__38616),
            .I(n2624));
    InMux I__7512 (
            .O(N__38611),
            .I(N__38607));
    InMux I__7511 (
            .O(N__38610),
            .I(N__38604));
    LocalMux I__7510 (
            .O(N__38607),
            .I(N__38600));
    LocalMux I__7509 (
            .O(N__38604),
            .I(N__38597));
    InMux I__7508 (
            .O(N__38603),
            .I(N__38594));
    Span4Mux_h I__7507 (
            .O(N__38600),
            .I(N__38591));
    Span4Mux_v I__7506 (
            .O(N__38597),
            .I(N__38586));
    LocalMux I__7505 (
            .O(N__38594),
            .I(N__38586));
    Odrv4 I__7504 (
            .O(N__38591),
            .I(n2617));
    Odrv4 I__7503 (
            .O(N__38586),
            .I(n2617));
    InMux I__7502 (
            .O(N__38581),
            .I(N__38578));
    LocalMux I__7501 (
            .O(N__38578),
            .I(N__38575));
    Span4Mux_h I__7500 (
            .O(N__38575),
            .I(N__38572));
    Odrv4 I__7499 (
            .O(N__38572),
            .I(n2684));
    InMux I__7498 (
            .O(N__38569),
            .I(N__38566));
    LocalMux I__7497 (
            .O(N__38566),
            .I(N__38563));
    Span4Mux_v I__7496 (
            .O(N__38563),
            .I(N__38560));
    Odrv4 I__7495 (
            .O(N__38560),
            .I(n2701));
    CascadeMux I__7494 (
            .O(N__38557),
            .I(N__38554));
    InMux I__7493 (
            .O(N__38554),
            .I(N__38551));
    LocalMux I__7492 (
            .O(N__38551),
            .I(N__38546));
    InMux I__7491 (
            .O(N__38550),
            .I(N__38543));
    InMux I__7490 (
            .O(N__38549),
            .I(N__38540));
    Span4Mux_v I__7489 (
            .O(N__38546),
            .I(N__38537));
    LocalMux I__7488 (
            .O(N__38543),
            .I(N__38532));
    LocalMux I__7487 (
            .O(N__38540),
            .I(N__38532));
    Odrv4 I__7486 (
            .O(N__38537),
            .I(n2613));
    Odrv12 I__7485 (
            .O(N__38532),
            .I(n2613));
    CascadeMux I__7484 (
            .O(N__38527),
            .I(N__38524));
    InMux I__7483 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__7482 (
            .O(N__38521),
            .I(N__38518));
    Span4Mux_h I__7481 (
            .O(N__38518),
            .I(N__38515));
    Odrv4 I__7480 (
            .O(N__38515),
            .I(n2680));
    InMux I__7479 (
            .O(N__38512),
            .I(N__38508));
    InMux I__7478 (
            .O(N__38511),
            .I(N__38505));
    LocalMux I__7477 (
            .O(N__38508),
            .I(N__38501));
    LocalMux I__7476 (
            .O(N__38505),
            .I(N__38498));
    InMux I__7475 (
            .O(N__38504),
            .I(N__38495));
    Span4Mux_h I__7474 (
            .O(N__38501),
            .I(N__38492));
    Span4Mux_h I__7473 (
            .O(N__38498),
            .I(N__38487));
    LocalMux I__7472 (
            .O(N__38495),
            .I(N__38487));
    Odrv4 I__7471 (
            .O(N__38492),
            .I(n2611));
    Odrv4 I__7470 (
            .O(N__38487),
            .I(n2611));
    InMux I__7469 (
            .O(N__38482),
            .I(N__38479));
    LocalMux I__7468 (
            .O(N__38479),
            .I(N__38476));
    Span4Mux_h I__7467 (
            .O(N__38476),
            .I(N__38473));
    Odrv4 I__7466 (
            .O(N__38473),
            .I(n2678));
    InMux I__7465 (
            .O(N__38470),
            .I(N__38465));
    InMux I__7464 (
            .O(N__38469),
            .I(N__38462));
    CascadeMux I__7463 (
            .O(N__38468),
            .I(N__38459));
    LocalMux I__7462 (
            .O(N__38465),
            .I(N__38456));
    LocalMux I__7461 (
            .O(N__38462),
            .I(N__38453));
    InMux I__7460 (
            .O(N__38459),
            .I(N__38450));
    Span4Mux_v I__7459 (
            .O(N__38456),
            .I(N__38447));
    Span4Mux_v I__7458 (
            .O(N__38453),
            .I(N__38442));
    LocalMux I__7457 (
            .O(N__38450),
            .I(N__38442));
    Odrv4 I__7456 (
            .O(N__38447),
            .I(n2615));
    Odrv4 I__7455 (
            .O(N__38442),
            .I(n2615));
    CascadeMux I__7454 (
            .O(N__38437),
            .I(N__38434));
    InMux I__7453 (
            .O(N__38434),
            .I(N__38431));
    LocalMux I__7452 (
            .O(N__38431),
            .I(N__38428));
    Span4Mux_h I__7451 (
            .O(N__38428),
            .I(N__38425));
    Odrv4 I__7450 (
            .O(N__38425),
            .I(n2682));
    CascadeMux I__7449 (
            .O(N__38422),
            .I(n45_cascade_));
    InMux I__7448 (
            .O(N__38419),
            .I(N__38416));
    LocalMux I__7447 (
            .O(N__38416),
            .I(n16_adj_614));
    CascadeMux I__7446 (
            .O(N__38413),
            .I(n14843_cascade_));
    InMux I__7445 (
            .O(N__38410),
            .I(N__38407));
    LocalMux I__7444 (
            .O(N__38407),
            .I(n24_adj_619));
    CascadeMux I__7443 (
            .O(N__38404),
            .I(n14711_cascade_));
    InMux I__7442 (
            .O(N__38401),
            .I(N__38398));
    LocalMux I__7441 (
            .O(N__38398),
            .I(n8_adj_607));
    InMux I__7440 (
            .O(N__38395),
            .I(N__38390));
    InMux I__7439 (
            .O(N__38394),
            .I(N__38385));
    InMux I__7438 (
            .O(N__38393),
            .I(N__38385));
    LocalMux I__7437 (
            .O(N__38390),
            .I(n45));
    LocalMux I__7436 (
            .O(N__38385),
            .I(n45));
    CascadeMux I__7435 (
            .O(N__38380),
            .I(n14826_cascade_));
    InMux I__7434 (
            .O(N__38377),
            .I(N__38374));
    LocalMux I__7433 (
            .O(N__38374),
            .I(n14779));
    InMux I__7432 (
            .O(N__38371),
            .I(N__38368));
    LocalMux I__7431 (
            .O(N__38368),
            .I(N__38365));
    Odrv4 I__7430 (
            .O(N__38365),
            .I(n14864));
    CascadeMux I__7429 (
            .O(N__38362),
            .I(N__38359));
    InMux I__7428 (
            .O(N__38359),
            .I(N__38355));
    InMux I__7427 (
            .O(N__38358),
            .I(N__38352));
    LocalMux I__7426 (
            .O(N__38355),
            .I(n43));
    LocalMux I__7425 (
            .O(N__38352),
            .I(n43));
    InMux I__7424 (
            .O(N__38347),
            .I(N__38344));
    LocalMux I__7423 (
            .O(N__38344),
            .I(n14713));
    InMux I__7422 (
            .O(N__38341),
            .I(N__38338));
    LocalMux I__7421 (
            .O(N__38338),
            .I(N__38335));
    Span4Mux_h I__7420 (
            .O(N__38335),
            .I(N__38332));
    Odrv4 I__7419 (
            .O(N__38332),
            .I(n2700));
    CascadeMux I__7418 (
            .O(N__38329),
            .I(n41_cascade_));
    InMux I__7417 (
            .O(N__38326),
            .I(N__38323));
    LocalMux I__7416 (
            .O(N__38323),
            .I(n41));
    CascadeMux I__7415 (
            .O(N__38320),
            .I(n14715_cascade_));
    InMux I__7414 (
            .O(N__38317),
            .I(N__38314));
    LocalMux I__7413 (
            .O(N__38314),
            .I(n40));
    CascadeMux I__7412 (
            .O(N__38311),
            .I(n14866_cascade_));
    CascadeMux I__7411 (
            .O(N__38308),
            .I(n12_adj_598_cascade_));
    InMux I__7410 (
            .O(N__38305),
            .I(N__38301));
    InMux I__7409 (
            .O(N__38304),
            .I(N__38298));
    LocalMux I__7408 (
            .O(N__38301),
            .I(N__38294));
    LocalMux I__7407 (
            .O(N__38298),
            .I(N__38291));
    InMux I__7406 (
            .O(N__38297),
            .I(N__38288));
    Span4Mux_v I__7405 (
            .O(N__38294),
            .I(N__38283));
    Span4Mux_v I__7404 (
            .O(N__38291),
            .I(N__38283));
    LocalMux I__7403 (
            .O(N__38288),
            .I(encoder0_position_13));
    Odrv4 I__7402 (
            .O(N__38283),
            .I(encoder0_position_13));
    CascadeMux I__7401 (
            .O(N__38278),
            .I(N__38275));
    InMux I__7400 (
            .O(N__38275),
            .I(N__38272));
    LocalMux I__7399 (
            .O(N__38272),
            .I(N__38269));
    Span4Mux_h I__7398 (
            .O(N__38269),
            .I(N__38266));
    Odrv4 I__7397 (
            .O(N__38266),
            .I(n20_adj_644));
    InMux I__7396 (
            .O(N__38263),
            .I(N__38258));
    InMux I__7395 (
            .O(N__38262),
            .I(N__38252));
    InMux I__7394 (
            .O(N__38261),
            .I(N__38252));
    LocalMux I__7393 (
            .O(N__38258),
            .I(N__38249));
    InMux I__7392 (
            .O(N__38257),
            .I(N__38246));
    LocalMux I__7391 (
            .O(N__38252),
            .I(N__38243));
    Span4Mux_h I__7390 (
            .O(N__38249),
            .I(N__38240));
    LocalMux I__7389 (
            .O(N__38246),
            .I(encoder0_position_28));
    Odrv4 I__7388 (
            .O(N__38243),
            .I(encoder0_position_28));
    Odrv4 I__7387 (
            .O(N__38240),
            .I(encoder0_position_28));
    CascadeMux I__7386 (
            .O(N__38233),
            .I(N__38230));
    InMux I__7385 (
            .O(N__38230),
            .I(N__38227));
    LocalMux I__7384 (
            .O(N__38227),
            .I(N__38224));
    Odrv4 I__7383 (
            .O(N__38224),
            .I(n5_adj_629));
    InMux I__7382 (
            .O(N__38221),
            .I(N__38218));
    LocalMux I__7381 (
            .O(N__38218),
            .I(N__38215));
    Odrv4 I__7380 (
            .O(N__38215),
            .I(encoder0_position_scaled_9));
    InMux I__7379 (
            .O(N__38212),
            .I(N__38209));
    LocalMux I__7378 (
            .O(N__38209),
            .I(N__38206));
    Odrv4 I__7377 (
            .O(N__38206),
            .I(encoder0_position_scaled_10));
    CascadeMux I__7376 (
            .O(N__38203),
            .I(N__38200));
    InMux I__7375 (
            .O(N__38200),
            .I(N__38193));
    InMux I__7374 (
            .O(N__38199),
            .I(N__38193));
    InMux I__7373 (
            .O(N__38198),
            .I(N__38188));
    LocalMux I__7372 (
            .O(N__38193),
            .I(N__38185));
    InMux I__7371 (
            .O(N__38192),
            .I(N__38182));
    InMux I__7370 (
            .O(N__38191),
            .I(N__38179));
    LocalMux I__7369 (
            .O(N__38188),
            .I(N__38172));
    Span4Mux_h I__7368 (
            .O(N__38185),
            .I(N__38172));
    LocalMux I__7367 (
            .O(N__38182),
            .I(N__38172));
    LocalMux I__7366 (
            .O(N__38179),
            .I(N__38166));
    Span4Mux_v I__7365 (
            .O(N__38172),
            .I(N__38166));
    InMux I__7364 (
            .O(N__38171),
            .I(N__38163));
    Span4Mux_h I__7363 (
            .O(N__38166),
            .I(N__38160));
    LocalMux I__7362 (
            .O(N__38163),
            .I(h2));
    Odrv4 I__7361 (
            .O(N__38160),
            .I(h2));
    InMux I__7360 (
            .O(N__38155),
            .I(N__38151));
    InMux I__7359 (
            .O(N__38154),
            .I(N__38145));
    LocalMux I__7358 (
            .O(N__38151),
            .I(N__38142));
    InMux I__7357 (
            .O(N__38150),
            .I(N__38139));
    InMux I__7356 (
            .O(N__38149),
            .I(N__38136));
    InMux I__7355 (
            .O(N__38148),
            .I(N__38133));
    LocalMux I__7354 (
            .O(N__38145),
            .I(N__38129));
    Span4Mux_s2_v I__7353 (
            .O(N__38142),
            .I(N__38126));
    LocalMux I__7352 (
            .O(N__38139),
            .I(N__38119));
    LocalMux I__7351 (
            .O(N__38136),
            .I(N__38119));
    LocalMux I__7350 (
            .O(N__38133),
            .I(N__38119));
    InMux I__7349 (
            .O(N__38132),
            .I(N__38116));
    Span12Mux_s6_v I__7348 (
            .O(N__38129),
            .I(N__38113));
    Span4Mux_v I__7347 (
            .O(N__38126),
            .I(N__38110));
    Span4Mux_v I__7346 (
            .O(N__38119),
            .I(N__38107));
    LocalMux I__7345 (
            .O(N__38116),
            .I(h3));
    Odrv12 I__7344 (
            .O(N__38113),
            .I(h3));
    Odrv4 I__7343 (
            .O(N__38110),
            .I(h3));
    Odrv4 I__7342 (
            .O(N__38107),
            .I(h3));
    InMux I__7341 (
            .O(N__38098),
            .I(N__38092));
    InMux I__7340 (
            .O(N__38097),
            .I(N__38089));
    InMux I__7339 (
            .O(N__38096),
            .I(N__38083));
    InMux I__7338 (
            .O(N__38095),
            .I(N__38083));
    LocalMux I__7337 (
            .O(N__38092),
            .I(N__38080));
    LocalMux I__7336 (
            .O(N__38089),
            .I(N__38077));
    InMux I__7335 (
            .O(N__38088),
            .I(N__38074));
    LocalMux I__7334 (
            .O(N__38083),
            .I(N__38071));
    Span4Mux_h I__7333 (
            .O(N__38080),
            .I(N__38065));
    Span4Mux_h I__7332 (
            .O(N__38077),
            .I(N__38065));
    LocalMux I__7331 (
            .O(N__38074),
            .I(N__38062));
    Span4Mux_h I__7330 (
            .O(N__38071),
            .I(N__38059));
    InMux I__7329 (
            .O(N__38070),
            .I(N__38056));
    Span4Mux_h I__7328 (
            .O(N__38065),
            .I(N__38053));
    Span4Mux_h I__7327 (
            .O(N__38062),
            .I(N__38048));
    Span4Mux_h I__7326 (
            .O(N__38059),
            .I(N__38048));
    LocalMux I__7325 (
            .O(N__38056),
            .I(h1));
    Odrv4 I__7324 (
            .O(N__38053),
            .I(h1));
    Odrv4 I__7323 (
            .O(N__38048),
            .I(h1));
    CEMux I__7322 (
            .O(N__38041),
            .I(N__38038));
    LocalMux I__7321 (
            .O(N__38038),
            .I(N__38035));
    Span4Mux_v I__7320 (
            .O(N__38035),
            .I(N__38032));
    Odrv4 I__7319 (
            .O(N__38032),
            .I(n6_adj_592));
    SRMux I__7318 (
            .O(N__38029),
            .I(N__38026));
    LocalMux I__7317 (
            .O(N__38026),
            .I(N__38023));
    Span4Mux_h I__7316 (
            .O(N__38023),
            .I(N__38020));
    Odrv4 I__7315 (
            .O(N__38020),
            .I(commutation_state_7__N_261));
    InMux I__7314 (
            .O(N__38017),
            .I(N__38014));
    LocalMux I__7313 (
            .O(N__38014),
            .I(encoder0_position_scaled_4));
    CascadeMux I__7312 (
            .O(N__38011),
            .I(dti_N_333_cascade_));
    InMux I__7311 (
            .O(N__38008),
            .I(N__38005));
    LocalMux I__7310 (
            .O(N__38005),
            .I(encoder0_position_scaled_22));
    InMux I__7309 (
            .O(N__38002),
            .I(N__37999));
    LocalMux I__7308 (
            .O(N__37999),
            .I(N__37996));
    Span4Mux_h I__7307 (
            .O(N__37996),
            .I(N__37993));
    Odrv4 I__7306 (
            .O(N__37993),
            .I(n26));
    InMux I__7305 (
            .O(N__37990),
            .I(N__37987));
    LocalMux I__7304 (
            .O(N__37987),
            .I(N__37983));
    CascadeMux I__7303 (
            .O(N__37986),
            .I(N__37980));
    Span4Mux_h I__7302 (
            .O(N__37983),
            .I(N__37977));
    InMux I__7301 (
            .O(N__37980),
            .I(N__37973));
    Span4Mux_v I__7300 (
            .O(N__37977),
            .I(N__37970));
    InMux I__7299 (
            .O(N__37976),
            .I(N__37967));
    LocalMux I__7298 (
            .O(N__37973),
            .I(encoder0_position_7));
    Odrv4 I__7297 (
            .O(N__37970),
            .I(encoder0_position_7));
    LocalMux I__7296 (
            .O(N__37967),
            .I(encoder0_position_7));
    InMux I__7295 (
            .O(N__37960),
            .I(N__37957));
    LocalMux I__7294 (
            .O(N__37957),
            .I(encoder0_position_scaled_19));
    InMux I__7293 (
            .O(N__37954),
            .I(N__37951));
    LocalMux I__7292 (
            .O(N__37951),
            .I(encoder0_position_scaled_21));
    InMux I__7291 (
            .O(N__37948),
            .I(N__37945));
    LocalMux I__7290 (
            .O(N__37945),
            .I(encoder0_position_scaled_13));
    CEMux I__7289 (
            .O(N__37942),
            .I(N__37939));
    LocalMux I__7288 (
            .O(N__37939),
            .I(N__37936));
    Span4Mux_h I__7287 (
            .O(N__37936),
            .I(N__37933));
    Odrv4 I__7286 (
            .O(N__37933),
            .I(n4828));
    CascadeMux I__7285 (
            .O(N__37930),
            .I(n11593_cascade_));
    CascadeMux I__7284 (
            .O(N__37927),
            .I(n59_cascade_));
    CascadeMux I__7283 (
            .O(N__37924),
            .I(N__37920));
    InMux I__7282 (
            .O(N__37923),
            .I(N__37917));
    InMux I__7281 (
            .O(N__37920),
            .I(N__37914));
    LocalMux I__7280 (
            .O(N__37917),
            .I(n11838));
    LocalMux I__7279 (
            .O(N__37914),
            .I(n11838));
    InMux I__7278 (
            .O(N__37909),
            .I(N__37906));
    LocalMux I__7277 (
            .O(N__37906),
            .I(encoder0_position_scaled_0));
    InMux I__7276 (
            .O(N__37903),
            .I(N__37900));
    LocalMux I__7275 (
            .O(N__37900),
            .I(encoder0_position_scaled_15));
    InMux I__7274 (
            .O(N__37897),
            .I(N__37894));
    LocalMux I__7273 (
            .O(N__37894),
            .I(encoder0_position_scaled_12));
    InMux I__7272 (
            .O(N__37891),
            .I(N__37888));
    LocalMux I__7271 (
            .O(N__37888),
            .I(encoder0_position_scaled_2));
    InMux I__7270 (
            .O(N__37885),
            .I(n12461));
    InMux I__7269 (
            .O(N__37882),
            .I(n12462));
    InMux I__7268 (
            .O(N__37879),
            .I(n12463));
    InMux I__7267 (
            .O(N__37876),
            .I(N__37873));
    LocalMux I__7266 (
            .O(N__37873),
            .I(n15197));
    InMux I__7265 (
            .O(N__37870),
            .I(bfn_10_23_0_));
    InMux I__7264 (
            .O(N__37867),
            .I(n12453));
    InMux I__7263 (
            .O(N__37864),
            .I(n12454));
    InMux I__7262 (
            .O(N__37861),
            .I(n12455));
    InMux I__7261 (
            .O(N__37858),
            .I(n12456));
    InMux I__7260 (
            .O(N__37855),
            .I(n12457));
    InMux I__7259 (
            .O(N__37852),
            .I(n12458));
    InMux I__7258 (
            .O(N__37849),
            .I(n12459));
    InMux I__7257 (
            .O(N__37846),
            .I(bfn_10_24_0_));
    InMux I__7256 (
            .O(N__37843),
            .I(n12443));
    InMux I__7255 (
            .O(N__37840),
            .I(bfn_10_22_0_));
    InMux I__7254 (
            .O(N__37837),
            .I(n12445));
    InMux I__7253 (
            .O(N__37834),
            .I(n12446));
    InMux I__7252 (
            .O(N__37831),
            .I(n12447));
    InMux I__7251 (
            .O(N__37828),
            .I(n12448));
    InMux I__7250 (
            .O(N__37825),
            .I(n12449));
    InMux I__7249 (
            .O(N__37822),
            .I(n12450));
    InMux I__7248 (
            .O(N__37819),
            .I(n12451));
    CascadeMux I__7247 (
            .O(N__37816),
            .I(n3117_cascade_));
    InMux I__7246 (
            .O(N__37813),
            .I(N__37810));
    LocalMux I__7245 (
            .O(N__37810),
            .I(n13888));
    InMux I__7244 (
            .O(N__37807),
            .I(N__37804));
    LocalMux I__7243 (
            .O(N__37804),
            .I(n13886));
    InMux I__7242 (
            .O(N__37801),
            .I(bfn_10_21_0_));
    InMux I__7241 (
            .O(N__37798),
            .I(n12437));
    InMux I__7240 (
            .O(N__37795),
            .I(n12438));
    InMux I__7239 (
            .O(N__37792),
            .I(n12439));
    InMux I__7238 (
            .O(N__37789),
            .I(n12440));
    InMux I__7237 (
            .O(N__37786),
            .I(n12441));
    InMux I__7236 (
            .O(N__37783),
            .I(n12442));
    InMux I__7235 (
            .O(N__37780),
            .I(N__37777));
    LocalMux I__7234 (
            .O(N__37777),
            .I(N__37773));
    InMux I__7233 (
            .O(N__37776),
            .I(N__37769));
    Span4Mux_h I__7232 (
            .O(N__37773),
            .I(N__37766));
    InMux I__7231 (
            .O(N__37772),
            .I(N__37763));
    LocalMux I__7230 (
            .O(N__37769),
            .I(N__37758));
    Span4Mux_v I__7229 (
            .O(N__37766),
            .I(N__37758));
    LocalMux I__7228 (
            .O(N__37763),
            .I(encoder0_position_6));
    Odrv4 I__7227 (
            .O(N__37758),
            .I(encoder0_position_6));
    CascadeMux I__7226 (
            .O(N__37753),
            .I(N__37750));
    InMux I__7225 (
            .O(N__37750),
            .I(N__37747));
    LocalMux I__7224 (
            .O(N__37747),
            .I(N__37744));
    Span4Mux_v I__7223 (
            .O(N__37744),
            .I(N__37741));
    Span4Mux_h I__7222 (
            .O(N__37741),
            .I(N__37738));
    Odrv4 I__7221 (
            .O(N__37738),
            .I(n27_adj_651));
    InMux I__7220 (
            .O(N__37735),
            .I(N__37732));
    LocalMux I__7219 (
            .O(N__37732),
            .I(N__37729));
    Span4Mux_v I__7218 (
            .O(N__37729),
            .I(N__37726));
    Span4Mux_v I__7217 (
            .O(N__37726),
            .I(N__37723));
    Odrv4 I__7216 (
            .O(N__37723),
            .I(n24));
    InMux I__7215 (
            .O(N__37720),
            .I(N__37717));
    LocalMux I__7214 (
            .O(N__37717),
            .I(N__37714));
    Span4Mux_v I__7213 (
            .O(N__37714),
            .I(N__37709));
    InMux I__7212 (
            .O(N__37713),
            .I(N__37706));
    InMux I__7211 (
            .O(N__37712),
            .I(N__37703));
    Span4Mux_h I__7210 (
            .O(N__37709),
            .I(N__37700));
    LocalMux I__7209 (
            .O(N__37706),
            .I(N__37697));
    LocalMux I__7208 (
            .O(N__37703),
            .I(encoder0_position_9));
    Odrv4 I__7207 (
            .O(N__37700),
            .I(encoder0_position_9));
    Odrv12 I__7206 (
            .O(N__37697),
            .I(encoder0_position_9));
    InMux I__7205 (
            .O(N__37690),
            .I(N__37687));
    LocalMux I__7204 (
            .O(N__37687),
            .I(N__37683));
    InMux I__7203 (
            .O(N__37686),
            .I(N__37680));
    Span4Mux_v I__7202 (
            .O(N__37683),
            .I(N__37674));
    LocalMux I__7201 (
            .O(N__37680),
            .I(N__37674));
    InMux I__7200 (
            .O(N__37679),
            .I(N__37671));
    Span4Mux_h I__7199 (
            .O(N__37674),
            .I(N__37668));
    LocalMux I__7198 (
            .O(N__37671),
            .I(N__37665));
    Span4Mux_h I__7197 (
            .O(N__37668),
            .I(N__37662));
    Span12Mux_s9_h I__7196 (
            .O(N__37665),
            .I(N__37659));
    Odrv4 I__7195 (
            .O(N__37662),
            .I(n310));
    Odrv12 I__7194 (
            .O(N__37659),
            .I(n310));
    InMux I__7193 (
            .O(N__37654),
            .I(N__37651));
    LocalMux I__7192 (
            .O(N__37651),
            .I(N__37648));
    Span4Mux_v I__7191 (
            .O(N__37648),
            .I(N__37645));
    Span4Mux_v I__7190 (
            .O(N__37645),
            .I(N__37642));
    Span4Mux_h I__7189 (
            .O(N__37642),
            .I(N__37639));
    Odrv4 I__7188 (
            .O(N__37639),
            .I(n19));
    InMux I__7187 (
            .O(N__37636),
            .I(N__37633));
    LocalMux I__7186 (
            .O(N__37633),
            .I(N__37629));
    CascadeMux I__7185 (
            .O(N__37632),
            .I(N__37625));
    Span4Mux_h I__7184 (
            .O(N__37629),
            .I(N__37622));
    InMux I__7183 (
            .O(N__37628),
            .I(N__37619));
    InMux I__7182 (
            .O(N__37625),
            .I(N__37616));
    Span4Mux_v I__7181 (
            .O(N__37622),
            .I(N__37613));
    LocalMux I__7180 (
            .O(N__37619),
            .I(N__37610));
    LocalMux I__7179 (
            .O(N__37616),
            .I(encoder0_position_14));
    Odrv4 I__7178 (
            .O(N__37613),
            .I(encoder0_position_14));
    Odrv4 I__7177 (
            .O(N__37610),
            .I(encoder0_position_14));
    InMux I__7176 (
            .O(N__37603),
            .I(N__37600));
    LocalMux I__7175 (
            .O(N__37600),
            .I(N__37595));
    InMux I__7174 (
            .O(N__37599),
            .I(N__37592));
    InMux I__7173 (
            .O(N__37598),
            .I(N__37589));
    Span4Mux_v I__7172 (
            .O(N__37595),
            .I(N__37586));
    LocalMux I__7171 (
            .O(N__37592),
            .I(N__37581));
    LocalMux I__7170 (
            .O(N__37589),
            .I(N__37581));
    Span4Mux_h I__7169 (
            .O(N__37586),
            .I(N__37576));
    Span4Mux_v I__7168 (
            .O(N__37581),
            .I(N__37576));
    Span4Mux_h I__7167 (
            .O(N__37576),
            .I(N__37573));
    Odrv4 I__7166 (
            .O(N__37573),
            .I(n305));
    InMux I__7165 (
            .O(N__37570),
            .I(N__37567));
    LocalMux I__7164 (
            .O(N__37567),
            .I(N__37564));
    Span4Mux_v I__7163 (
            .O(N__37564),
            .I(N__37561));
    Span4Mux_v I__7162 (
            .O(N__37561),
            .I(N__37558));
    Odrv4 I__7161 (
            .O(N__37558),
            .I(n23));
    InMux I__7160 (
            .O(N__37555),
            .I(N__37551));
    InMux I__7159 (
            .O(N__37554),
            .I(N__37548));
    LocalMux I__7158 (
            .O(N__37551),
            .I(N__37544));
    LocalMux I__7157 (
            .O(N__37548),
            .I(N__37541));
    CascadeMux I__7156 (
            .O(N__37547),
            .I(N__37538));
    Span4Mux_h I__7155 (
            .O(N__37544),
            .I(N__37535));
    Span4Mux_v I__7154 (
            .O(N__37541),
            .I(N__37532));
    InMux I__7153 (
            .O(N__37538),
            .I(N__37529));
    Span4Mux_v I__7152 (
            .O(N__37535),
            .I(N__37526));
    Span4Mux_v I__7151 (
            .O(N__37532),
            .I(N__37523));
    LocalMux I__7150 (
            .O(N__37529),
            .I(encoder0_position_10));
    Odrv4 I__7149 (
            .O(N__37526),
            .I(encoder0_position_10));
    Odrv4 I__7148 (
            .O(N__37523),
            .I(encoder0_position_10));
    InMux I__7147 (
            .O(N__37516),
            .I(N__37513));
    LocalMux I__7146 (
            .O(N__37513),
            .I(N__37509));
    InMux I__7145 (
            .O(N__37512),
            .I(N__37506));
    Span4Mux_v I__7144 (
            .O(N__37509),
            .I(N__37500));
    LocalMux I__7143 (
            .O(N__37506),
            .I(N__37500));
    InMux I__7142 (
            .O(N__37505),
            .I(N__37497));
    Span4Mux_h I__7141 (
            .O(N__37500),
            .I(N__37494));
    LocalMux I__7140 (
            .O(N__37497),
            .I(N__37491));
    Span4Mux_h I__7139 (
            .O(N__37494),
            .I(N__37488));
    Odrv12 I__7138 (
            .O(N__37491),
            .I(n309));
    Odrv4 I__7137 (
            .O(N__37488),
            .I(n309));
    CascadeMux I__7136 (
            .O(N__37483),
            .I(N__37479));
    InMux I__7135 (
            .O(N__37482),
            .I(N__37476));
    InMux I__7134 (
            .O(N__37479),
            .I(N__37473));
    LocalMux I__7133 (
            .O(N__37476),
            .I(N__37467));
    LocalMux I__7132 (
            .O(N__37473),
            .I(N__37467));
    InMux I__7131 (
            .O(N__37472),
            .I(N__37464));
    Span4Mux_v I__7130 (
            .O(N__37467),
            .I(N__37459));
    LocalMux I__7129 (
            .O(N__37464),
            .I(N__37459));
    Odrv4 I__7128 (
            .O(N__37459),
            .I(n2616));
    CascadeMux I__7127 (
            .O(N__37456),
            .I(N__37453));
    InMux I__7126 (
            .O(N__37453),
            .I(N__37450));
    LocalMux I__7125 (
            .O(N__37450),
            .I(N__37447));
    Odrv4 I__7124 (
            .O(N__37447),
            .I(n2683));
    CascadeMux I__7123 (
            .O(N__37444),
            .I(n13884_cascade_));
    CascadeMux I__7122 (
            .O(N__37441),
            .I(N__37437));
    InMux I__7121 (
            .O(N__37440),
            .I(N__37434));
    InMux I__7120 (
            .O(N__37437),
            .I(N__37431));
    LocalMux I__7119 (
            .O(N__37434),
            .I(N__37426));
    LocalMux I__7118 (
            .O(N__37431),
            .I(N__37426));
    Span4Mux_v I__7117 (
            .O(N__37426),
            .I(N__37422));
    InMux I__7116 (
            .O(N__37425),
            .I(N__37419));
    Odrv4 I__7115 (
            .O(N__37422),
            .I(n2627));
    LocalMux I__7114 (
            .O(N__37419),
            .I(n2627));
    CascadeMux I__7113 (
            .O(N__37414),
            .I(N__37411));
    InMux I__7112 (
            .O(N__37411),
            .I(N__37408));
    LocalMux I__7111 (
            .O(N__37408),
            .I(n2694));
    InMux I__7110 (
            .O(N__37405),
            .I(N__37401));
    CascadeMux I__7109 (
            .O(N__37404),
            .I(N__37398));
    LocalMux I__7108 (
            .O(N__37401),
            .I(N__37395));
    InMux I__7107 (
            .O(N__37398),
            .I(N__37392));
    Span4Mux_h I__7106 (
            .O(N__37395),
            .I(N__37388));
    LocalMux I__7105 (
            .O(N__37392),
            .I(N__37385));
    InMux I__7104 (
            .O(N__37391),
            .I(N__37382));
    Odrv4 I__7103 (
            .O(N__37388),
            .I(n2521));
    Odrv4 I__7102 (
            .O(N__37385),
            .I(n2521));
    LocalMux I__7101 (
            .O(N__37382),
            .I(n2521));
    CascadeMux I__7100 (
            .O(N__37375),
            .I(N__37372));
    InMux I__7099 (
            .O(N__37372),
            .I(N__37369));
    LocalMux I__7098 (
            .O(N__37369),
            .I(N__37366));
    Span4Mux_v I__7097 (
            .O(N__37366),
            .I(N__37363));
    Odrv4 I__7096 (
            .O(N__37363),
            .I(n2588));
    CascadeMux I__7095 (
            .O(N__37360),
            .I(N__37357));
    InMux I__7094 (
            .O(N__37357),
            .I(N__37354));
    LocalMux I__7093 (
            .O(N__37354),
            .I(N__37350));
    InMux I__7092 (
            .O(N__37353),
            .I(N__37347));
    Odrv4 I__7091 (
            .O(N__37350),
            .I(n2620));
    LocalMux I__7090 (
            .O(N__37347),
            .I(n2620));
    InMux I__7089 (
            .O(N__37342),
            .I(N__37339));
    LocalMux I__7088 (
            .O(N__37339),
            .I(N__37336));
    Odrv4 I__7087 (
            .O(N__37336),
            .I(n2687));
    CascadeMux I__7086 (
            .O(N__37333),
            .I(n2620_cascade_));
    InMux I__7085 (
            .O(N__37330),
            .I(N__37327));
    LocalMux I__7084 (
            .O(N__37327),
            .I(N__37323));
    InMux I__7083 (
            .O(N__37326),
            .I(N__37320));
    Span4Mux_h I__7082 (
            .O(N__37323),
            .I(N__37317));
    LocalMux I__7081 (
            .O(N__37320),
            .I(N__37314));
    Span4Mux_v I__7080 (
            .O(N__37317),
            .I(N__37309));
    Span4Mux_h I__7079 (
            .O(N__37314),
            .I(N__37309));
    Odrv4 I__7078 (
            .O(N__37309),
            .I(n2610));
    CascadeMux I__7077 (
            .O(N__37306),
            .I(N__37303));
    InMux I__7076 (
            .O(N__37303),
            .I(N__37300));
    LocalMux I__7075 (
            .O(N__37300),
            .I(n14300));
    InMux I__7074 (
            .O(N__37297),
            .I(N__37293));
    InMux I__7073 (
            .O(N__37296),
            .I(N__37289));
    LocalMux I__7072 (
            .O(N__37293),
            .I(N__37286));
    InMux I__7071 (
            .O(N__37292),
            .I(N__37283));
    LocalMux I__7070 (
            .O(N__37289),
            .I(n2621));
    Odrv4 I__7069 (
            .O(N__37286),
            .I(n2621));
    LocalMux I__7068 (
            .O(N__37283),
            .I(n2621));
    CascadeMux I__7067 (
            .O(N__37276),
            .I(n2643_cascade_));
    InMux I__7066 (
            .O(N__37273),
            .I(N__37270));
    LocalMux I__7065 (
            .O(N__37270),
            .I(N__37267));
    Span4Mux_v I__7064 (
            .O(N__37267),
            .I(N__37264));
    Span4Mux_h I__7063 (
            .O(N__37264),
            .I(N__37261));
    Odrv4 I__7062 (
            .O(N__37261),
            .I(n2688));
    CascadeMux I__7061 (
            .O(N__37258),
            .I(n2720_cascade_));
    CascadeMux I__7060 (
            .O(N__37255),
            .I(n14038_cascade_));
    InMux I__7059 (
            .O(N__37252),
            .I(N__37249));
    LocalMux I__7058 (
            .O(N__37249),
            .I(n14042));
    InMux I__7057 (
            .O(N__37246),
            .I(N__37241));
    InMux I__7056 (
            .O(N__37245),
            .I(N__37238));
    InMux I__7055 (
            .O(N__37244),
            .I(N__37235));
    LocalMux I__7054 (
            .O(N__37241),
            .I(N__37232));
    LocalMux I__7053 (
            .O(N__37238),
            .I(N__37229));
    LocalMux I__7052 (
            .O(N__37235),
            .I(N__37226));
    Span4Mux_h I__7051 (
            .O(N__37232),
            .I(N__37223));
    Span4Mux_h I__7050 (
            .O(N__37229),
            .I(N__37218));
    Span4Mux_h I__7049 (
            .O(N__37226),
            .I(N__37218));
    Odrv4 I__7048 (
            .O(N__37223),
            .I(n2614));
    Odrv4 I__7047 (
            .O(N__37218),
            .I(n2614));
    InMux I__7046 (
            .O(N__37213),
            .I(N__37210));
    LocalMux I__7045 (
            .O(N__37210),
            .I(N__37207));
    Span4Mux_h I__7044 (
            .O(N__37207),
            .I(N__37204));
    Odrv4 I__7043 (
            .O(N__37204),
            .I(n2681));
    InMux I__7042 (
            .O(N__37201),
            .I(N__37198));
    LocalMux I__7041 (
            .O(N__37198),
            .I(N__37195));
    Odrv4 I__7040 (
            .O(N__37195),
            .I(n2685));
    CascadeMux I__7039 (
            .O(N__37192),
            .I(N__37187));
    InMux I__7038 (
            .O(N__37191),
            .I(N__37184));
    InMux I__7037 (
            .O(N__37190),
            .I(N__37181));
    InMux I__7036 (
            .O(N__37187),
            .I(N__37178));
    LocalMux I__7035 (
            .O(N__37184),
            .I(N__37175));
    LocalMux I__7034 (
            .O(N__37181),
            .I(N__37172));
    LocalMux I__7033 (
            .O(N__37178),
            .I(N__37169));
    Span4Mux_h I__7032 (
            .O(N__37175),
            .I(N__37164));
    Span4Mux_h I__7031 (
            .O(N__37172),
            .I(N__37164));
    Odrv4 I__7030 (
            .O(N__37169),
            .I(n2618));
    Odrv4 I__7029 (
            .O(N__37164),
            .I(n2618));
    InMux I__7028 (
            .O(N__37159),
            .I(N__37156));
    LocalMux I__7027 (
            .O(N__37156),
            .I(n14294));
    InMux I__7026 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__7025 (
            .O(N__37150),
            .I(N__37147));
    Odrv4 I__7024 (
            .O(N__37147),
            .I(n2693));
    InMux I__7023 (
            .O(N__37144),
            .I(N__37140));
    InMux I__7022 (
            .O(N__37143),
            .I(N__37137));
    LocalMux I__7021 (
            .O(N__37140),
            .I(N__37134));
    LocalMux I__7020 (
            .O(N__37137),
            .I(n2626));
    Odrv4 I__7019 (
            .O(N__37134),
            .I(n2626));
    CascadeMux I__7018 (
            .O(N__37129),
            .I(n2725_cascade_));
    CascadeMux I__7017 (
            .O(N__37126),
            .I(n14040_cascade_));
    CascadeMux I__7016 (
            .O(N__37123),
            .I(N__37119));
    InMux I__7015 (
            .O(N__37122),
            .I(N__37115));
    InMux I__7014 (
            .O(N__37119),
            .I(N__37112));
    InMux I__7013 (
            .O(N__37118),
            .I(N__37109));
    LocalMux I__7012 (
            .O(N__37115),
            .I(n2629));
    LocalMux I__7011 (
            .O(N__37112),
            .I(n2629));
    LocalMux I__7010 (
            .O(N__37109),
            .I(n2629));
    CascadeMux I__7009 (
            .O(N__37102),
            .I(N__37099));
    InMux I__7008 (
            .O(N__37099),
            .I(N__37096));
    LocalMux I__7007 (
            .O(N__37096),
            .I(N__37093));
    Odrv4 I__7006 (
            .O(N__37093),
            .I(n2696));
    CascadeMux I__7005 (
            .O(N__37090),
            .I(N__37087));
    InMux I__7004 (
            .O(N__37087),
            .I(N__37083));
    InMux I__7003 (
            .O(N__37086),
            .I(N__37080));
    LocalMux I__7002 (
            .O(N__37083),
            .I(N__37077));
    LocalMux I__7001 (
            .O(N__37080),
            .I(n2630));
    Odrv4 I__7000 (
            .O(N__37077),
            .I(n2630));
    InMux I__6999 (
            .O(N__37072),
            .I(N__37069));
    LocalMux I__6998 (
            .O(N__37069),
            .I(N__37066));
    Odrv4 I__6997 (
            .O(N__37066),
            .I(n2697));
    InMux I__6996 (
            .O(N__37063),
            .I(N__37060));
    LocalMux I__6995 (
            .O(N__37060),
            .I(N__37057));
    Odrv4 I__6994 (
            .O(N__37057),
            .I(n2695));
    CascadeMux I__6993 (
            .O(N__37054),
            .I(N__37050));
    CascadeMux I__6992 (
            .O(N__37053),
            .I(N__37047));
    InMux I__6991 (
            .O(N__37050),
            .I(N__37044));
    InMux I__6990 (
            .O(N__37047),
            .I(N__37041));
    LocalMux I__6989 (
            .O(N__37044),
            .I(N__37038));
    LocalMux I__6988 (
            .O(N__37041),
            .I(N__37035));
    Span4Mux_h I__6987 (
            .O(N__37038),
            .I(N__37032));
    Odrv12 I__6986 (
            .O(N__37035),
            .I(n2628));
    Odrv4 I__6985 (
            .O(N__37032),
            .I(n2628));
    CascadeMux I__6984 (
            .O(N__37027),
            .I(N__37023));
    InMux I__6983 (
            .O(N__37026),
            .I(N__37020));
    InMux I__6982 (
            .O(N__37023),
            .I(N__37016));
    LocalMux I__6981 (
            .O(N__37020),
            .I(N__37013));
    InMux I__6980 (
            .O(N__37019),
            .I(N__37010));
    LocalMux I__6979 (
            .O(N__37016),
            .I(n2619));
    Odrv4 I__6978 (
            .O(N__37013),
            .I(n2619));
    LocalMux I__6977 (
            .O(N__37010),
            .I(n2619));
    InMux I__6976 (
            .O(N__37003),
            .I(N__37000));
    LocalMux I__6975 (
            .O(N__37000),
            .I(N__36997));
    Span4Mux_h I__6974 (
            .O(N__36997),
            .I(N__36994));
    Odrv4 I__6973 (
            .O(N__36994),
            .I(n2686));
    InMux I__6972 (
            .O(N__36991),
            .I(N__36988));
    LocalMux I__6971 (
            .O(N__36988),
            .I(encoder0_position_scaled_23));
    InMux I__6970 (
            .O(N__36985),
            .I(N__36982));
    LocalMux I__6969 (
            .O(N__36982),
            .I(N__36979));
    Span4Mux_h I__6968 (
            .O(N__36979),
            .I(N__36976));
    Span4Mux_h I__6967 (
            .O(N__36976),
            .I(N__36973));
    Odrv4 I__6966 (
            .O(N__36973),
            .I(ENCODER0_A_N));
    InMux I__6965 (
            .O(N__36970),
            .I(N__36967));
    LocalMux I__6964 (
            .O(N__36967),
            .I(N__36963));
    InMux I__6963 (
            .O(N__36966),
            .I(N__36960));
    Span4Mux_v I__6962 (
            .O(N__36963),
            .I(N__36952));
    LocalMux I__6961 (
            .O(N__36960),
            .I(N__36952));
    CascadeMux I__6960 (
            .O(N__36959),
            .I(N__36945));
    CascadeMux I__6959 (
            .O(N__36958),
            .I(N__36942));
    InMux I__6958 (
            .O(N__36957),
            .I(N__36938));
    Span4Mux_h I__6957 (
            .O(N__36952),
            .I(N__36935));
    InMux I__6956 (
            .O(N__36951),
            .I(N__36932));
    InMux I__6955 (
            .O(N__36950),
            .I(N__36925));
    InMux I__6954 (
            .O(N__36949),
            .I(N__36925));
    InMux I__6953 (
            .O(N__36948),
            .I(N__36925));
    InMux I__6952 (
            .O(N__36945),
            .I(N__36918));
    InMux I__6951 (
            .O(N__36942),
            .I(N__36918));
    InMux I__6950 (
            .O(N__36941),
            .I(N__36918));
    LocalMux I__6949 (
            .O(N__36938),
            .I(N__36915));
    Odrv4 I__6948 (
            .O(N__36935),
            .I(n1059));
    LocalMux I__6947 (
            .O(N__36932),
            .I(n1059));
    LocalMux I__6946 (
            .O(N__36925),
            .I(n1059));
    LocalMux I__6945 (
            .O(N__36918),
            .I(n1059));
    Odrv4 I__6944 (
            .O(N__36915),
            .I(n1059));
    InMux I__6943 (
            .O(N__36904),
            .I(N__36901));
    LocalMux I__6942 (
            .O(N__36901),
            .I(N__36898));
    Span4Mux_h I__6941 (
            .O(N__36898),
            .I(N__36895));
    Odrv4 I__6940 (
            .O(N__36895),
            .I(n15210));
    CascadeMux I__6939 (
            .O(N__36892),
            .I(n14536_cascade_));
    InMux I__6938 (
            .O(N__36889),
            .I(N__36886));
    LocalMux I__6937 (
            .O(N__36886),
            .I(N__36883));
    Span12Mux_v I__6936 (
            .O(N__36883),
            .I(N__36879));
    InMux I__6935 (
            .O(N__36882),
            .I(N__36876));
    Odrv12 I__6934 (
            .O(N__36879),
            .I(blink_counter_25));
    LocalMux I__6933 (
            .O(N__36876),
            .I(blink_counter_25));
    IoInMux I__6932 (
            .O(N__36871),
            .I(N__36868));
    LocalMux I__6931 (
            .O(N__36868),
            .I(N__36865));
    Span4Mux_s2_v I__6930 (
            .O(N__36865),
            .I(N__36862));
    Span4Mux_h I__6929 (
            .O(N__36862),
            .I(N__36859));
    Odrv4 I__6928 (
            .O(N__36859),
            .I(LED_c));
    InMux I__6927 (
            .O(N__36856),
            .I(N__36850));
    InMux I__6926 (
            .O(N__36855),
            .I(N__36850));
    LocalMux I__6925 (
            .O(N__36850),
            .I(N__36847));
    Span4Mux_v I__6924 (
            .O(N__36847),
            .I(N__36844));
    Span4Mux_h I__6923 (
            .O(N__36844),
            .I(N__36840));
    InMux I__6922 (
            .O(N__36843),
            .I(N__36837));
    Odrv4 I__6921 (
            .O(N__36840),
            .I(blink_counter_24));
    LocalMux I__6920 (
            .O(N__36837),
            .I(blink_counter_24));
    InMux I__6919 (
            .O(N__36832),
            .I(N__36826));
    InMux I__6918 (
            .O(N__36831),
            .I(N__36826));
    LocalMux I__6917 (
            .O(N__36826),
            .I(N__36822));
    InMux I__6916 (
            .O(N__36825),
            .I(N__36819));
    Odrv12 I__6915 (
            .O(N__36822),
            .I(blink_counter_21));
    LocalMux I__6914 (
            .O(N__36819),
            .I(blink_counter_21));
    CascadeMux I__6913 (
            .O(N__36814),
            .I(N__36810));
    InMux I__6912 (
            .O(N__36813),
            .I(N__36805));
    InMux I__6911 (
            .O(N__36810),
            .I(N__36805));
    LocalMux I__6910 (
            .O(N__36805),
            .I(N__36801));
    InMux I__6909 (
            .O(N__36804),
            .I(N__36798));
    Odrv12 I__6908 (
            .O(N__36801),
            .I(blink_counter_22));
    LocalMux I__6907 (
            .O(N__36798),
            .I(blink_counter_22));
    CascadeMux I__6906 (
            .O(N__36793),
            .I(N__36790));
    InMux I__6905 (
            .O(N__36790),
            .I(N__36784));
    InMux I__6904 (
            .O(N__36789),
            .I(N__36784));
    LocalMux I__6903 (
            .O(N__36784),
            .I(N__36780));
    InMux I__6902 (
            .O(N__36783),
            .I(N__36777));
    Odrv12 I__6901 (
            .O(N__36780),
            .I(blink_counter_23));
    LocalMux I__6900 (
            .O(N__36777),
            .I(blink_counter_23));
    InMux I__6899 (
            .O(N__36772),
            .I(N__36769));
    LocalMux I__6898 (
            .O(N__36769),
            .I(n14535));
    InMux I__6897 (
            .O(N__36766),
            .I(N__36763));
    LocalMux I__6896 (
            .O(N__36763),
            .I(N__36760));
    Span4Mux_v I__6895 (
            .O(N__36760),
            .I(N__36757));
    Span4Mux_h I__6894 (
            .O(N__36757),
            .I(N__36753));
    InMux I__6893 (
            .O(N__36756),
            .I(N__36750));
    Odrv4 I__6892 (
            .O(N__36753),
            .I(n15259));
    LocalMux I__6891 (
            .O(N__36750),
            .I(n15259));
    InMux I__6890 (
            .O(N__36745),
            .I(N__36740));
    InMux I__6889 (
            .O(N__36744),
            .I(N__36734));
    InMux I__6888 (
            .O(N__36743),
            .I(N__36734));
    LocalMux I__6887 (
            .O(N__36740),
            .I(N__36729));
    CascadeMux I__6886 (
            .O(N__36739),
            .I(N__36726));
    LocalMux I__6885 (
            .O(N__36734),
            .I(N__36722));
    CascadeMux I__6884 (
            .O(N__36733),
            .I(N__36716));
    CascadeMux I__6883 (
            .O(N__36732),
            .I(N__36712));
    Span12Mux_v I__6882 (
            .O(N__36729),
            .I(N__36708));
    InMux I__6881 (
            .O(N__36726),
            .I(N__36703));
    InMux I__6880 (
            .O(N__36725),
            .I(N__36703));
    Span4Mux_s3_h I__6879 (
            .O(N__36722),
            .I(N__36700));
    InMux I__6878 (
            .O(N__36721),
            .I(N__36695));
    InMux I__6877 (
            .O(N__36720),
            .I(N__36695));
    InMux I__6876 (
            .O(N__36719),
            .I(N__36684));
    InMux I__6875 (
            .O(N__36716),
            .I(N__36684));
    InMux I__6874 (
            .O(N__36715),
            .I(N__36684));
    InMux I__6873 (
            .O(N__36712),
            .I(N__36684));
    InMux I__6872 (
            .O(N__36711),
            .I(N__36684));
    Odrv12 I__6871 (
            .O(N__36708),
            .I(n1356));
    LocalMux I__6870 (
            .O(N__36703),
            .I(n1356));
    Odrv4 I__6869 (
            .O(N__36700),
            .I(n1356));
    LocalMux I__6868 (
            .O(N__36695),
            .I(n1356));
    LocalMux I__6867 (
            .O(N__36684),
            .I(n1356));
    InMux I__6866 (
            .O(N__36673),
            .I(n12571));
    InMux I__6865 (
            .O(N__36670),
            .I(N__36667));
    LocalMux I__6864 (
            .O(N__36667),
            .I(N__36664));
    Span4Mux_v I__6863 (
            .O(N__36664),
            .I(N__36660));
    InMux I__6862 (
            .O(N__36663),
            .I(N__36657));
    Span4Mux_h I__6861 (
            .O(N__36660),
            .I(N__36654));
    LocalMux I__6860 (
            .O(N__36657),
            .I(N__36651));
    Odrv4 I__6859 (
            .O(N__36654),
            .I(n15243));
    Odrv4 I__6858 (
            .O(N__36651),
            .I(n15243));
    CascadeMux I__6857 (
            .O(N__36646),
            .I(N__36643));
    InMux I__6856 (
            .O(N__36643),
            .I(N__36640));
    LocalMux I__6855 (
            .O(N__36640),
            .I(N__36637));
    Span4Mux_v I__6854 (
            .O(N__36637),
            .I(N__36632));
    CascadeMux I__6853 (
            .O(N__36636),
            .I(N__36622));
    CascadeMux I__6852 (
            .O(N__36635),
            .I(N__36619));
    Span4Mux_h I__6851 (
            .O(N__36632),
            .I(N__36615));
    InMux I__6850 (
            .O(N__36631),
            .I(N__36612));
    InMux I__6849 (
            .O(N__36630),
            .I(N__36609));
    InMux I__6848 (
            .O(N__36629),
            .I(N__36604));
    InMux I__6847 (
            .O(N__36628),
            .I(N__36604));
    InMux I__6846 (
            .O(N__36627),
            .I(N__36601));
    InMux I__6845 (
            .O(N__36626),
            .I(N__36590));
    InMux I__6844 (
            .O(N__36625),
            .I(N__36590));
    InMux I__6843 (
            .O(N__36622),
            .I(N__36590));
    InMux I__6842 (
            .O(N__36619),
            .I(N__36590));
    InMux I__6841 (
            .O(N__36618),
            .I(N__36590));
    Odrv4 I__6840 (
            .O(N__36615),
            .I(n1257));
    LocalMux I__6839 (
            .O(N__36612),
            .I(n1257));
    LocalMux I__6838 (
            .O(N__36609),
            .I(n1257));
    LocalMux I__6837 (
            .O(N__36604),
            .I(n1257));
    LocalMux I__6836 (
            .O(N__36601),
            .I(n1257));
    LocalMux I__6835 (
            .O(N__36590),
            .I(n1257));
    InMux I__6834 (
            .O(N__36577),
            .I(n12572));
    InMux I__6833 (
            .O(N__36574),
            .I(N__36571));
    LocalMux I__6832 (
            .O(N__36571),
            .I(N__36567));
    InMux I__6831 (
            .O(N__36570),
            .I(N__36564));
    Span4Mux_h I__6830 (
            .O(N__36567),
            .I(N__36561));
    LocalMux I__6829 (
            .O(N__36564),
            .I(N__36558));
    Span4Mux_v I__6828 (
            .O(N__36561),
            .I(N__36553));
    Span4Mux_s1_v I__6827 (
            .O(N__36558),
            .I(N__36553));
    Odrv4 I__6826 (
            .O(N__36553),
            .I(n15224));
    InMux I__6825 (
            .O(N__36550),
            .I(N__36547));
    LocalMux I__6824 (
            .O(N__36547),
            .I(N__36542));
    CascadeMux I__6823 (
            .O(N__36546),
            .I(N__36533));
    CascadeMux I__6822 (
            .O(N__36545),
            .I(N__36530));
    Span12Mux_v I__6821 (
            .O(N__36542),
            .I(N__36526));
    InMux I__6820 (
            .O(N__36541),
            .I(N__36523));
    InMux I__6819 (
            .O(N__36540),
            .I(N__36520));
    InMux I__6818 (
            .O(N__36539),
            .I(N__36515));
    InMux I__6817 (
            .O(N__36538),
            .I(N__36515));
    InMux I__6816 (
            .O(N__36537),
            .I(N__36512));
    InMux I__6815 (
            .O(N__36536),
            .I(N__36503));
    InMux I__6814 (
            .O(N__36533),
            .I(N__36503));
    InMux I__6813 (
            .O(N__36530),
            .I(N__36503));
    InMux I__6812 (
            .O(N__36529),
            .I(N__36503));
    Odrv12 I__6811 (
            .O(N__36526),
            .I(n1158));
    LocalMux I__6810 (
            .O(N__36523),
            .I(n1158));
    LocalMux I__6809 (
            .O(N__36520),
            .I(n1158));
    LocalMux I__6808 (
            .O(N__36515),
            .I(n1158));
    LocalMux I__6807 (
            .O(N__36512),
            .I(n1158));
    LocalMux I__6806 (
            .O(N__36503),
            .I(n1158));
    InMux I__6805 (
            .O(N__36490),
            .I(n12573));
    CascadeMux I__6804 (
            .O(N__36487),
            .I(N__36466));
    CascadeMux I__6803 (
            .O(N__36486),
            .I(N__36463));
    CascadeMux I__6802 (
            .O(N__36485),
            .I(N__36459));
    CascadeMux I__6801 (
            .O(N__36484),
            .I(N__36455));
    CascadeMux I__6800 (
            .O(N__36483),
            .I(N__36451));
    CascadeMux I__6799 (
            .O(N__36482),
            .I(N__36448));
    CascadeMux I__6798 (
            .O(N__36481),
            .I(N__36445));
    CascadeMux I__6797 (
            .O(N__36480),
            .I(N__36442));
    CascadeMux I__6796 (
            .O(N__36479),
            .I(N__36439));
    CascadeMux I__6795 (
            .O(N__36478),
            .I(N__36435));
    CascadeMux I__6794 (
            .O(N__36477),
            .I(N__36432));
    CascadeMux I__6793 (
            .O(N__36476),
            .I(N__36429));
    CascadeMux I__6792 (
            .O(N__36475),
            .I(N__36426));
    CascadeMux I__6791 (
            .O(N__36474),
            .I(N__36423));
    CascadeMux I__6790 (
            .O(N__36473),
            .I(N__36420));
    CascadeMux I__6789 (
            .O(N__36472),
            .I(N__36417));
    CascadeMux I__6788 (
            .O(N__36471),
            .I(N__36413));
    CascadeMux I__6787 (
            .O(N__36470),
            .I(N__36410));
    CascadeMux I__6786 (
            .O(N__36469),
            .I(N__36407));
    InMux I__6785 (
            .O(N__36466),
            .I(N__36403));
    InMux I__6784 (
            .O(N__36463),
            .I(N__36388));
    InMux I__6783 (
            .O(N__36462),
            .I(N__36388));
    InMux I__6782 (
            .O(N__36459),
            .I(N__36388));
    InMux I__6781 (
            .O(N__36458),
            .I(N__36388));
    InMux I__6780 (
            .O(N__36455),
            .I(N__36388));
    InMux I__6779 (
            .O(N__36454),
            .I(N__36388));
    InMux I__6778 (
            .O(N__36451),
            .I(N__36388));
    InMux I__6777 (
            .O(N__36448),
            .I(N__36379));
    InMux I__6776 (
            .O(N__36445),
            .I(N__36379));
    InMux I__6775 (
            .O(N__36442),
            .I(N__36379));
    InMux I__6774 (
            .O(N__36439),
            .I(N__36379));
    CascadeMux I__6773 (
            .O(N__36438),
            .I(N__36376));
    InMux I__6772 (
            .O(N__36435),
            .I(N__36367));
    InMux I__6771 (
            .O(N__36432),
            .I(N__36367));
    InMux I__6770 (
            .O(N__36429),
            .I(N__36367));
    InMux I__6769 (
            .O(N__36426),
            .I(N__36367));
    InMux I__6768 (
            .O(N__36423),
            .I(N__36362));
    InMux I__6767 (
            .O(N__36420),
            .I(N__36362));
    InMux I__6766 (
            .O(N__36417),
            .I(N__36349));
    InMux I__6765 (
            .O(N__36416),
            .I(N__36349));
    InMux I__6764 (
            .O(N__36413),
            .I(N__36349));
    InMux I__6763 (
            .O(N__36410),
            .I(N__36349));
    InMux I__6762 (
            .O(N__36407),
            .I(N__36349));
    InMux I__6761 (
            .O(N__36406),
            .I(N__36349));
    LocalMux I__6760 (
            .O(N__36403),
            .I(N__36342));
    LocalMux I__6759 (
            .O(N__36388),
            .I(N__36342));
    LocalMux I__6758 (
            .O(N__36379),
            .I(N__36342));
    InMux I__6757 (
            .O(N__36376),
            .I(N__36339));
    LocalMux I__6756 (
            .O(N__36367),
            .I(N__36332));
    LocalMux I__6755 (
            .O(N__36362),
            .I(N__36332));
    LocalMux I__6754 (
            .O(N__36349),
            .I(N__36332));
    Span4Mux_v I__6753 (
            .O(N__36342),
            .I(N__36327));
    LocalMux I__6752 (
            .O(N__36339),
            .I(N__36327));
    Span4Mux_v I__6751 (
            .O(N__36332),
            .I(N__36324));
    Span4Mux_h I__6750 (
            .O(N__36327),
            .I(N__36321));
    Odrv4 I__6749 (
            .O(N__36324),
            .I(n2_adj_626));
    Odrv4 I__6748 (
            .O(N__36321),
            .I(n2_adj_626));
    InMux I__6747 (
            .O(N__36316),
            .I(n12574));
    InMux I__6746 (
            .O(N__36313),
            .I(N__36310));
    LocalMux I__6745 (
            .O(N__36310),
            .I(encoder0_position_scaled_17));
    InMux I__6744 (
            .O(N__36307),
            .I(N__36304));
    LocalMux I__6743 (
            .O(N__36304),
            .I(encoder0_position_scaled_20));
    CascadeMux I__6742 (
            .O(N__36301),
            .I(N__36298));
    InMux I__6741 (
            .O(N__36298),
            .I(N__36294));
    CascadeMux I__6740 (
            .O(N__36297),
            .I(N__36291));
    LocalMux I__6739 (
            .O(N__36294),
            .I(N__36288));
    InMux I__6738 (
            .O(N__36291),
            .I(N__36284));
    Span4Mux_h I__6737 (
            .O(N__36288),
            .I(N__36281));
    InMux I__6736 (
            .O(N__36287),
            .I(N__36278));
    LocalMux I__6735 (
            .O(N__36284),
            .I(encoder0_position_25));
    Odrv4 I__6734 (
            .O(N__36281),
            .I(encoder0_position_25));
    LocalMux I__6733 (
            .O(N__36278),
            .I(encoder0_position_25));
    InMux I__6732 (
            .O(N__36271),
            .I(N__36268));
    LocalMux I__6731 (
            .O(N__36268),
            .I(N__36265));
    Odrv4 I__6730 (
            .O(N__36265),
            .I(n8));
    InMux I__6729 (
            .O(N__36262),
            .I(N__36255));
    InMux I__6728 (
            .O(N__36261),
            .I(N__36255));
    InMux I__6727 (
            .O(N__36260),
            .I(N__36252));
    LocalMux I__6726 (
            .O(N__36255),
            .I(N__36249));
    LocalMux I__6725 (
            .O(N__36252),
            .I(N__36246));
    Span4Mux_v I__6724 (
            .O(N__36249),
            .I(N__36243));
    Span4Mux_h I__6723 (
            .O(N__36246),
            .I(N__36240));
    Odrv4 I__6722 (
            .O(N__36243),
            .I(n294));
    Odrv4 I__6721 (
            .O(N__36240),
            .I(n294));
    InMux I__6720 (
            .O(N__36235),
            .I(N__36232));
    LocalMux I__6719 (
            .O(N__36232),
            .I(N__36229));
    Span4Mux_v I__6718 (
            .O(N__36229),
            .I(N__36226));
    Span4Mux_v I__6717 (
            .O(N__36226),
            .I(N__36223));
    Span4Mux_h I__6716 (
            .O(N__36223),
            .I(N__36219));
    InMux I__6715 (
            .O(N__36222),
            .I(N__36216));
    Odrv4 I__6714 (
            .O(N__36219),
            .I(n15059));
    LocalMux I__6713 (
            .O(N__36216),
            .I(n15059));
    InMux I__6712 (
            .O(N__36211),
            .I(N__36208));
    LocalMux I__6711 (
            .O(N__36208),
            .I(N__36202));
    CascadeMux I__6710 (
            .O(N__36207),
            .I(N__36195));
    CascadeMux I__6709 (
            .O(N__36206),
            .I(N__36188));
    InMux I__6708 (
            .O(N__36205),
            .I(N__36185));
    Span4Mux_v I__6707 (
            .O(N__36202),
            .I(N__36182));
    InMux I__6706 (
            .O(N__36201),
            .I(N__36177));
    InMux I__6705 (
            .O(N__36200),
            .I(N__36177));
    InMux I__6704 (
            .O(N__36199),
            .I(N__36174));
    CascadeMux I__6703 (
            .O(N__36198),
            .I(N__36170));
    InMux I__6702 (
            .O(N__36195),
            .I(N__36163));
    InMux I__6701 (
            .O(N__36194),
            .I(N__36163));
    CascadeMux I__6700 (
            .O(N__36193),
            .I(N__36160));
    CascadeMux I__6699 (
            .O(N__36192),
            .I(N__36154));
    CascadeMux I__6698 (
            .O(N__36191),
            .I(N__36151));
    InMux I__6697 (
            .O(N__36188),
            .I(N__36146));
    LocalMux I__6696 (
            .O(N__36185),
            .I(N__36143));
    Span4Mux_h I__6695 (
            .O(N__36182),
            .I(N__36136));
    LocalMux I__6694 (
            .O(N__36177),
            .I(N__36136));
    LocalMux I__6693 (
            .O(N__36174),
            .I(N__36136));
    InMux I__6692 (
            .O(N__36173),
            .I(N__36129));
    InMux I__6691 (
            .O(N__36170),
            .I(N__36129));
    InMux I__6690 (
            .O(N__36169),
            .I(N__36129));
    InMux I__6689 (
            .O(N__36168),
            .I(N__36126));
    LocalMux I__6688 (
            .O(N__36163),
            .I(N__36123));
    InMux I__6687 (
            .O(N__36160),
            .I(N__36118));
    InMux I__6686 (
            .O(N__36159),
            .I(N__36118));
    InMux I__6685 (
            .O(N__36158),
            .I(N__36113));
    InMux I__6684 (
            .O(N__36157),
            .I(N__36113));
    InMux I__6683 (
            .O(N__36154),
            .I(N__36104));
    InMux I__6682 (
            .O(N__36151),
            .I(N__36104));
    InMux I__6681 (
            .O(N__36150),
            .I(N__36104));
    InMux I__6680 (
            .O(N__36149),
            .I(N__36104));
    LocalMux I__6679 (
            .O(N__36146),
            .I(N__36097));
    Span4Mux_v I__6678 (
            .O(N__36143),
            .I(N__36097));
    Span4Mux_v I__6677 (
            .O(N__36136),
            .I(N__36097));
    LocalMux I__6676 (
            .O(N__36129),
            .I(N__36094));
    LocalMux I__6675 (
            .O(N__36126),
            .I(N__36089));
    Span4Mux_h I__6674 (
            .O(N__36123),
            .I(N__36089));
    LocalMux I__6673 (
            .O(N__36118),
            .I(n2148));
    LocalMux I__6672 (
            .O(N__36113),
            .I(n2148));
    LocalMux I__6671 (
            .O(N__36104),
            .I(n2148));
    Odrv4 I__6670 (
            .O(N__36097),
            .I(n2148));
    Odrv12 I__6669 (
            .O(N__36094),
            .I(n2148));
    Odrv4 I__6668 (
            .O(N__36089),
            .I(n2148));
    InMux I__6667 (
            .O(N__36076),
            .I(n12563));
    InMux I__6666 (
            .O(N__36073),
            .I(N__36069));
    CascadeMux I__6665 (
            .O(N__36072),
            .I(N__36066));
    LocalMux I__6664 (
            .O(N__36069),
            .I(N__36063));
    InMux I__6663 (
            .O(N__36066),
            .I(N__36060));
    Span12Mux_h I__6662 (
            .O(N__36063),
            .I(N__36057));
    LocalMux I__6661 (
            .O(N__36060),
            .I(N__36054));
    Odrv12 I__6660 (
            .O(N__36057),
            .I(n15035));
    Odrv4 I__6659 (
            .O(N__36054),
            .I(n15035));
    InMux I__6658 (
            .O(N__36049),
            .I(N__36046));
    LocalMux I__6657 (
            .O(N__36046),
            .I(N__36041));
    CascadeMux I__6656 (
            .O(N__36045),
            .I(N__36038));
    InMux I__6655 (
            .O(N__36044),
            .I(N__36033));
    Span4Mux_v I__6654 (
            .O(N__36041),
            .I(N__36028));
    InMux I__6653 (
            .O(N__36038),
            .I(N__36025));
    InMux I__6652 (
            .O(N__36037),
            .I(N__36022));
    InMux I__6651 (
            .O(N__36036),
            .I(N__36019));
    LocalMux I__6650 (
            .O(N__36033),
            .I(N__36012));
    InMux I__6649 (
            .O(N__36032),
            .I(N__36007));
    InMux I__6648 (
            .O(N__36031),
            .I(N__36007));
    Span4Mux_h I__6647 (
            .O(N__36028),
            .I(N__35998));
    LocalMux I__6646 (
            .O(N__36025),
            .I(N__35998));
    LocalMux I__6645 (
            .O(N__36022),
            .I(N__35998));
    LocalMux I__6644 (
            .O(N__36019),
            .I(N__35998));
    InMux I__6643 (
            .O(N__36018),
            .I(N__35995));
    CascadeMux I__6642 (
            .O(N__36017),
            .I(N__35988));
    CascadeMux I__6641 (
            .O(N__36016),
            .I(N__35982));
    CascadeMux I__6640 (
            .O(N__36015),
            .I(N__35979));
    Span4Mux_h I__6639 (
            .O(N__36012),
            .I(N__35969));
    LocalMux I__6638 (
            .O(N__36007),
            .I(N__35969));
    Span4Mux_v I__6637 (
            .O(N__35998),
            .I(N__35969));
    LocalMux I__6636 (
            .O(N__35995),
            .I(N__35969));
    InMux I__6635 (
            .O(N__35994),
            .I(N__35966));
    InMux I__6634 (
            .O(N__35993),
            .I(N__35963));
    InMux I__6633 (
            .O(N__35992),
            .I(N__35960));
    InMux I__6632 (
            .O(N__35991),
            .I(N__35957));
    InMux I__6631 (
            .O(N__35988),
            .I(N__35950));
    InMux I__6630 (
            .O(N__35987),
            .I(N__35950));
    InMux I__6629 (
            .O(N__35986),
            .I(N__35950));
    InMux I__6628 (
            .O(N__35985),
            .I(N__35941));
    InMux I__6627 (
            .O(N__35982),
            .I(N__35941));
    InMux I__6626 (
            .O(N__35979),
            .I(N__35941));
    InMux I__6625 (
            .O(N__35978),
            .I(N__35941));
    Span4Mux_h I__6624 (
            .O(N__35969),
            .I(N__35938));
    LocalMux I__6623 (
            .O(N__35966),
            .I(n2049));
    LocalMux I__6622 (
            .O(N__35963),
            .I(n2049));
    LocalMux I__6621 (
            .O(N__35960),
            .I(n2049));
    LocalMux I__6620 (
            .O(N__35957),
            .I(n2049));
    LocalMux I__6619 (
            .O(N__35950),
            .I(n2049));
    LocalMux I__6618 (
            .O(N__35941),
            .I(n2049));
    Odrv4 I__6617 (
            .O(N__35938),
            .I(n2049));
    InMux I__6616 (
            .O(N__35923),
            .I(n12564));
    InMux I__6615 (
            .O(N__35920),
            .I(N__35917));
    LocalMux I__6614 (
            .O(N__35917),
            .I(N__35914));
    Span4Mux_h I__6613 (
            .O(N__35914),
            .I(N__35911));
    Span4Mux_h I__6612 (
            .O(N__35911),
            .I(N__35907));
    InMux I__6611 (
            .O(N__35910),
            .I(N__35904));
    Odrv4 I__6610 (
            .O(N__35907),
            .I(n15012));
    LocalMux I__6609 (
            .O(N__35904),
            .I(n15012));
    InMux I__6608 (
            .O(N__35899),
            .I(N__35896));
    LocalMux I__6607 (
            .O(N__35896),
            .I(N__35891));
    InMux I__6606 (
            .O(N__35895),
            .I(N__35885));
    CascadeMux I__6605 (
            .O(N__35894),
            .I(N__35882));
    Span4Mux_h I__6604 (
            .O(N__35891),
            .I(N__35879));
    CascadeMux I__6603 (
            .O(N__35890),
            .I(N__35876));
    CascadeMux I__6602 (
            .O(N__35889),
            .I(N__35864));
    CascadeMux I__6601 (
            .O(N__35888),
            .I(N__35859));
    LocalMux I__6600 (
            .O(N__35885),
            .I(N__35855));
    InMux I__6599 (
            .O(N__35882),
            .I(N__35852));
    Span4Mux_v I__6598 (
            .O(N__35879),
            .I(N__35849));
    InMux I__6597 (
            .O(N__35876),
            .I(N__35846));
    InMux I__6596 (
            .O(N__35875),
            .I(N__35843));
    InMux I__6595 (
            .O(N__35874),
            .I(N__35838));
    InMux I__6594 (
            .O(N__35873),
            .I(N__35838));
    InMux I__6593 (
            .O(N__35872),
            .I(N__35835));
    InMux I__6592 (
            .O(N__35871),
            .I(N__35832));
    InMux I__6591 (
            .O(N__35870),
            .I(N__35825));
    InMux I__6590 (
            .O(N__35869),
            .I(N__35825));
    InMux I__6589 (
            .O(N__35868),
            .I(N__35825));
    InMux I__6588 (
            .O(N__35867),
            .I(N__35812));
    InMux I__6587 (
            .O(N__35864),
            .I(N__35812));
    InMux I__6586 (
            .O(N__35863),
            .I(N__35812));
    InMux I__6585 (
            .O(N__35862),
            .I(N__35812));
    InMux I__6584 (
            .O(N__35859),
            .I(N__35812));
    InMux I__6583 (
            .O(N__35858),
            .I(N__35812));
    Span4Mux_s3_h I__6582 (
            .O(N__35855),
            .I(N__35807));
    LocalMux I__6581 (
            .O(N__35852),
            .I(N__35807));
    Odrv4 I__6580 (
            .O(N__35849),
            .I(n1950));
    LocalMux I__6579 (
            .O(N__35846),
            .I(n1950));
    LocalMux I__6578 (
            .O(N__35843),
            .I(n1950));
    LocalMux I__6577 (
            .O(N__35838),
            .I(n1950));
    LocalMux I__6576 (
            .O(N__35835),
            .I(n1950));
    LocalMux I__6575 (
            .O(N__35832),
            .I(n1950));
    LocalMux I__6574 (
            .O(N__35825),
            .I(n1950));
    LocalMux I__6573 (
            .O(N__35812),
            .I(n1950));
    Odrv4 I__6572 (
            .O(N__35807),
            .I(n1950));
    InMux I__6571 (
            .O(N__35788),
            .I(n12565));
    InMux I__6570 (
            .O(N__35785),
            .I(N__35782));
    LocalMux I__6569 (
            .O(N__35782),
            .I(N__35779));
    Span4Mux_v I__6568 (
            .O(N__35779),
            .I(N__35776));
    Span4Mux_h I__6567 (
            .O(N__35776),
            .I(N__35773));
    Odrv4 I__6566 (
            .O(N__35773),
            .I(n14990));
    InMux I__6565 (
            .O(N__35770),
            .I(N__35767));
    LocalMux I__6564 (
            .O(N__35767),
            .I(N__35762));
    InMux I__6563 (
            .O(N__35766),
            .I(N__35758));
    InMux I__6562 (
            .O(N__35765),
            .I(N__35755));
    Span4Mux_h I__6561 (
            .O(N__35762),
            .I(N__35748));
    CascadeMux I__6560 (
            .O(N__35761),
            .I(N__35744));
    LocalMux I__6559 (
            .O(N__35758),
            .I(N__35741));
    LocalMux I__6558 (
            .O(N__35755),
            .I(N__35738));
    CascadeMux I__6557 (
            .O(N__35754),
            .I(N__35734));
    CascadeMux I__6556 (
            .O(N__35753),
            .I(N__35730));
    CascadeMux I__6555 (
            .O(N__35752),
            .I(N__35722));
    InMux I__6554 (
            .O(N__35751),
            .I(N__35717));
    Span4Mux_v I__6553 (
            .O(N__35748),
            .I(N__35714));
    InMux I__6552 (
            .O(N__35747),
            .I(N__35711));
    InMux I__6551 (
            .O(N__35744),
            .I(N__35708));
    Span4Mux_s3_h I__6550 (
            .O(N__35741),
            .I(N__35705));
    Span4Mux_s3_h I__6549 (
            .O(N__35738),
            .I(N__35702));
    InMux I__6548 (
            .O(N__35737),
            .I(N__35689));
    InMux I__6547 (
            .O(N__35734),
            .I(N__35689));
    InMux I__6546 (
            .O(N__35733),
            .I(N__35689));
    InMux I__6545 (
            .O(N__35730),
            .I(N__35689));
    InMux I__6544 (
            .O(N__35729),
            .I(N__35689));
    InMux I__6543 (
            .O(N__35728),
            .I(N__35689));
    InMux I__6542 (
            .O(N__35727),
            .I(N__35680));
    InMux I__6541 (
            .O(N__35726),
            .I(N__35680));
    InMux I__6540 (
            .O(N__35725),
            .I(N__35680));
    InMux I__6539 (
            .O(N__35722),
            .I(N__35680));
    InMux I__6538 (
            .O(N__35721),
            .I(N__35675));
    InMux I__6537 (
            .O(N__35720),
            .I(N__35675));
    LocalMux I__6536 (
            .O(N__35717),
            .I(n1851));
    Odrv4 I__6535 (
            .O(N__35714),
            .I(n1851));
    LocalMux I__6534 (
            .O(N__35711),
            .I(n1851));
    LocalMux I__6533 (
            .O(N__35708),
            .I(n1851));
    Odrv4 I__6532 (
            .O(N__35705),
            .I(n1851));
    Odrv4 I__6531 (
            .O(N__35702),
            .I(n1851));
    LocalMux I__6530 (
            .O(N__35689),
            .I(n1851));
    LocalMux I__6529 (
            .O(N__35680),
            .I(n1851));
    LocalMux I__6528 (
            .O(N__35675),
            .I(n1851));
    InMux I__6527 (
            .O(N__35656),
            .I(n12566));
    InMux I__6526 (
            .O(N__35653),
            .I(N__35650));
    LocalMux I__6525 (
            .O(N__35650),
            .I(N__35647));
    Span4Mux_v I__6524 (
            .O(N__35647),
            .I(N__35643));
    CascadeMux I__6523 (
            .O(N__35646),
            .I(N__35640));
    Span4Mux_h I__6522 (
            .O(N__35643),
            .I(N__35637));
    InMux I__6521 (
            .O(N__35640),
            .I(N__35634));
    Odrv4 I__6520 (
            .O(N__35637),
            .I(n14969));
    LocalMux I__6519 (
            .O(N__35634),
            .I(n14969));
    InMux I__6518 (
            .O(N__35629),
            .I(N__35625));
    CascadeMux I__6517 (
            .O(N__35628),
            .I(N__35616));
    LocalMux I__6516 (
            .O(N__35625),
            .I(N__35612));
    CascadeMux I__6515 (
            .O(N__35624),
            .I(N__35608));
    InMux I__6514 (
            .O(N__35623),
            .I(N__35604));
    CascadeMux I__6513 (
            .O(N__35622),
            .I(N__35601));
    CascadeMux I__6512 (
            .O(N__35621),
            .I(N__35596));
    InMux I__6511 (
            .O(N__35620),
            .I(N__35585));
    InMux I__6510 (
            .O(N__35619),
            .I(N__35585));
    InMux I__6509 (
            .O(N__35616),
            .I(N__35585));
    InMux I__6508 (
            .O(N__35615),
            .I(N__35585));
    Span4Mux_v I__6507 (
            .O(N__35612),
            .I(N__35581));
    InMux I__6506 (
            .O(N__35611),
            .I(N__35574));
    InMux I__6505 (
            .O(N__35608),
            .I(N__35574));
    InMux I__6504 (
            .O(N__35607),
            .I(N__35574));
    LocalMux I__6503 (
            .O(N__35604),
            .I(N__35571));
    InMux I__6502 (
            .O(N__35601),
            .I(N__35566));
    InMux I__6501 (
            .O(N__35600),
            .I(N__35566));
    InMux I__6500 (
            .O(N__35599),
            .I(N__35559));
    InMux I__6499 (
            .O(N__35596),
            .I(N__35559));
    InMux I__6498 (
            .O(N__35595),
            .I(N__35559));
    InMux I__6497 (
            .O(N__35594),
            .I(N__35556));
    LocalMux I__6496 (
            .O(N__35585),
            .I(N__35553));
    InMux I__6495 (
            .O(N__35584),
            .I(N__35550));
    Span4Mux_h I__6494 (
            .O(N__35581),
            .I(N__35543));
    LocalMux I__6493 (
            .O(N__35574),
            .I(N__35543));
    Span4Mux_v I__6492 (
            .O(N__35571),
            .I(N__35543));
    LocalMux I__6491 (
            .O(N__35566),
            .I(n1752));
    LocalMux I__6490 (
            .O(N__35559),
            .I(n1752));
    LocalMux I__6489 (
            .O(N__35556),
            .I(n1752));
    Odrv4 I__6488 (
            .O(N__35553),
            .I(n1752));
    LocalMux I__6487 (
            .O(N__35550),
            .I(n1752));
    Odrv4 I__6486 (
            .O(N__35543),
            .I(n1752));
    InMux I__6485 (
            .O(N__35530),
            .I(bfn_9_27_0_));
    InMux I__6484 (
            .O(N__35527),
            .I(N__35524));
    LocalMux I__6483 (
            .O(N__35524),
            .I(N__35521));
    Span4Mux_v I__6482 (
            .O(N__35521),
            .I(N__35517));
    InMux I__6481 (
            .O(N__35520),
            .I(N__35514));
    Span4Mux_h I__6480 (
            .O(N__35517),
            .I(N__35511));
    LocalMux I__6479 (
            .O(N__35514),
            .I(N__35508));
    Odrv4 I__6478 (
            .O(N__35511),
            .I(n14949));
    Odrv4 I__6477 (
            .O(N__35508),
            .I(n14949));
    CascadeMux I__6476 (
            .O(N__35503),
            .I(N__35500));
    InMux I__6475 (
            .O(N__35500),
            .I(N__35497));
    LocalMux I__6474 (
            .O(N__35497),
            .I(N__35494));
    Span4Mux_h I__6473 (
            .O(N__35494),
            .I(N__35488));
    CascadeMux I__6472 (
            .O(N__35493),
            .I(N__35477));
    CascadeMux I__6471 (
            .O(N__35492),
            .I(N__35473));
    CascadeMux I__6470 (
            .O(N__35491),
            .I(N__35470));
    Span4Mux_h I__6469 (
            .O(N__35488),
            .I(N__35465));
    InMux I__6468 (
            .O(N__35487),
            .I(N__35462));
    InMux I__6467 (
            .O(N__35486),
            .I(N__35455));
    InMux I__6466 (
            .O(N__35485),
            .I(N__35455));
    InMux I__6465 (
            .O(N__35484),
            .I(N__35455));
    InMux I__6464 (
            .O(N__35483),
            .I(N__35446));
    InMux I__6463 (
            .O(N__35482),
            .I(N__35446));
    InMux I__6462 (
            .O(N__35481),
            .I(N__35446));
    InMux I__6461 (
            .O(N__35480),
            .I(N__35446));
    InMux I__6460 (
            .O(N__35477),
            .I(N__35433));
    InMux I__6459 (
            .O(N__35476),
            .I(N__35433));
    InMux I__6458 (
            .O(N__35473),
            .I(N__35433));
    InMux I__6457 (
            .O(N__35470),
            .I(N__35433));
    InMux I__6456 (
            .O(N__35469),
            .I(N__35433));
    InMux I__6455 (
            .O(N__35468),
            .I(N__35433));
    Odrv4 I__6454 (
            .O(N__35465),
            .I(n1653));
    LocalMux I__6453 (
            .O(N__35462),
            .I(n1653));
    LocalMux I__6452 (
            .O(N__35455),
            .I(n1653));
    LocalMux I__6451 (
            .O(N__35446),
            .I(n1653));
    LocalMux I__6450 (
            .O(N__35433),
            .I(n1653));
    InMux I__6449 (
            .O(N__35422),
            .I(n12568));
    InMux I__6448 (
            .O(N__35419),
            .I(N__35416));
    LocalMux I__6447 (
            .O(N__35416),
            .I(N__35413));
    Span4Mux_v I__6446 (
            .O(N__35413),
            .I(N__35410));
    Span4Mux_h I__6445 (
            .O(N__35410),
            .I(N__35406));
    InMux I__6444 (
            .O(N__35409),
            .I(N__35403));
    Odrv4 I__6443 (
            .O(N__35406),
            .I(n15292));
    LocalMux I__6442 (
            .O(N__35403),
            .I(n15292));
    InMux I__6441 (
            .O(N__35398),
            .I(N__35395));
    LocalMux I__6440 (
            .O(N__35395),
            .I(N__35392));
    Span4Mux_h I__6439 (
            .O(N__35392),
            .I(N__35385));
    CascadeMux I__6438 (
            .O(N__35391),
            .I(N__35379));
    CascadeMux I__6437 (
            .O(N__35390),
            .I(N__35375));
    CascadeMux I__6436 (
            .O(N__35389),
            .I(N__35369));
    CascadeMux I__6435 (
            .O(N__35388),
            .I(N__35366));
    Span4Mux_h I__6434 (
            .O(N__35385),
            .I(N__35361));
    InMux I__6433 (
            .O(N__35384),
            .I(N__35356));
    InMux I__6432 (
            .O(N__35383),
            .I(N__35356));
    InMux I__6431 (
            .O(N__35382),
            .I(N__35353));
    InMux I__6430 (
            .O(N__35379),
            .I(N__35342));
    InMux I__6429 (
            .O(N__35378),
            .I(N__35342));
    InMux I__6428 (
            .O(N__35375),
            .I(N__35342));
    InMux I__6427 (
            .O(N__35374),
            .I(N__35342));
    InMux I__6426 (
            .O(N__35373),
            .I(N__35342));
    InMux I__6425 (
            .O(N__35372),
            .I(N__35331));
    InMux I__6424 (
            .O(N__35369),
            .I(N__35331));
    InMux I__6423 (
            .O(N__35366),
            .I(N__35331));
    InMux I__6422 (
            .O(N__35365),
            .I(N__35331));
    InMux I__6421 (
            .O(N__35364),
            .I(N__35331));
    Odrv4 I__6420 (
            .O(N__35361),
            .I(n1554));
    LocalMux I__6419 (
            .O(N__35356),
            .I(n1554));
    LocalMux I__6418 (
            .O(N__35353),
            .I(n1554));
    LocalMux I__6417 (
            .O(N__35342),
            .I(n1554));
    LocalMux I__6416 (
            .O(N__35331),
            .I(n1554));
    InMux I__6415 (
            .O(N__35320),
            .I(n12569));
    InMux I__6414 (
            .O(N__35317),
            .I(N__35314));
    LocalMux I__6413 (
            .O(N__35314),
            .I(N__35311));
    Span4Mux_h I__6412 (
            .O(N__35311),
            .I(N__35307));
    CascadeMux I__6411 (
            .O(N__35310),
            .I(N__35304));
    Span4Mux_h I__6410 (
            .O(N__35307),
            .I(N__35301));
    InMux I__6409 (
            .O(N__35304),
            .I(N__35298));
    Odrv4 I__6408 (
            .O(N__35301),
            .I(n15276));
    LocalMux I__6407 (
            .O(N__35298),
            .I(n15276));
    CascadeMux I__6406 (
            .O(N__35293),
            .I(N__35290));
    InMux I__6405 (
            .O(N__35290),
            .I(N__35287));
    LocalMux I__6404 (
            .O(N__35287),
            .I(N__35283));
    CascadeMux I__6403 (
            .O(N__35286),
            .I(N__35276));
    Span4Mux_h I__6402 (
            .O(N__35283),
            .I(N__35271));
    InMux I__6401 (
            .O(N__35282),
            .I(N__35268));
    CascadeMux I__6400 (
            .O(N__35281),
            .I(N__35265));
    CascadeMux I__6399 (
            .O(N__35280),
            .I(N__35262));
    CascadeMux I__6398 (
            .O(N__35279),
            .I(N__35259));
    InMux I__6397 (
            .O(N__35276),
            .I(N__35251));
    InMux I__6396 (
            .O(N__35275),
            .I(N__35251));
    CascadeMux I__6395 (
            .O(N__35274),
            .I(N__35248));
    Span4Mux_h I__6394 (
            .O(N__35271),
            .I(N__35243));
    LocalMux I__6393 (
            .O(N__35268),
            .I(N__35240));
    InMux I__6392 (
            .O(N__35265),
            .I(N__35231));
    InMux I__6391 (
            .O(N__35262),
            .I(N__35231));
    InMux I__6390 (
            .O(N__35259),
            .I(N__35231));
    InMux I__6389 (
            .O(N__35258),
            .I(N__35231));
    InMux I__6388 (
            .O(N__35257),
            .I(N__35228));
    InMux I__6387 (
            .O(N__35256),
            .I(N__35225));
    LocalMux I__6386 (
            .O(N__35251),
            .I(N__35222));
    InMux I__6385 (
            .O(N__35248),
            .I(N__35215));
    InMux I__6384 (
            .O(N__35247),
            .I(N__35215));
    InMux I__6383 (
            .O(N__35246),
            .I(N__35215));
    Odrv4 I__6382 (
            .O(N__35243),
            .I(n1455));
    Odrv4 I__6381 (
            .O(N__35240),
            .I(n1455));
    LocalMux I__6380 (
            .O(N__35231),
            .I(n1455));
    LocalMux I__6379 (
            .O(N__35228),
            .I(n1455));
    LocalMux I__6378 (
            .O(N__35225),
            .I(n1455));
    Odrv4 I__6377 (
            .O(N__35222),
            .I(n1455));
    LocalMux I__6376 (
            .O(N__35215),
            .I(n1455));
    InMux I__6375 (
            .O(N__35200),
            .I(n12570));
    InMux I__6374 (
            .O(N__35197),
            .I(n12555));
    InMux I__6373 (
            .O(N__35194),
            .I(n12556));
    InMux I__6372 (
            .O(N__35191),
            .I(n12557));
    InMux I__6371 (
            .O(N__35188),
            .I(N__35185));
    LocalMux I__6370 (
            .O(N__35185),
            .I(N__35181));
    CascadeMux I__6369 (
            .O(N__35184),
            .I(N__35178));
    Span4Mux_v I__6368 (
            .O(N__35181),
            .I(N__35175));
    InMux I__6367 (
            .O(N__35178),
            .I(N__35172));
    Odrv4 I__6366 (
            .O(N__35175),
            .I(n15437));
    LocalMux I__6365 (
            .O(N__35172),
            .I(n15437));
    InMux I__6364 (
            .O(N__35167),
            .I(n12558));
    InMux I__6363 (
            .O(N__35164),
            .I(N__35161));
    LocalMux I__6362 (
            .O(N__35161),
            .I(N__35158));
    Sp12to4 I__6361 (
            .O(N__35158),
            .I(N__35154));
    CascadeMux I__6360 (
            .O(N__35157),
            .I(N__35151));
    Span12Mux_v I__6359 (
            .O(N__35154),
            .I(N__35148));
    InMux I__6358 (
            .O(N__35151),
            .I(N__35145));
    Odrv12 I__6357 (
            .O(N__35148),
            .I(n15401));
    LocalMux I__6356 (
            .O(N__35145),
            .I(n15401));
    InMux I__6355 (
            .O(N__35140),
            .I(bfn_9_26_0_));
    InMux I__6354 (
            .O(N__35137),
            .I(N__35134));
    LocalMux I__6353 (
            .O(N__35134),
            .I(N__35130));
    CascadeMux I__6352 (
            .O(N__35133),
            .I(N__35127));
    Span4Mux_h I__6351 (
            .O(N__35130),
            .I(N__35124));
    InMux I__6350 (
            .O(N__35127),
            .I(N__35121));
    Sp12to4 I__6349 (
            .O(N__35124),
            .I(N__35116));
    LocalMux I__6348 (
            .O(N__35121),
            .I(N__35116));
    Odrv12 I__6347 (
            .O(N__35116),
            .I(n15375));
    InMux I__6346 (
            .O(N__35113),
            .I(N__35110));
    LocalMux I__6345 (
            .O(N__35110),
            .I(N__35098));
    CascadeMux I__6344 (
            .O(N__35109),
            .I(N__35094));
    CascadeMux I__6343 (
            .O(N__35108),
            .I(N__35089));
    CascadeMux I__6342 (
            .O(N__35107),
            .I(N__35086));
    CascadeMux I__6341 (
            .O(N__35106),
            .I(N__35081));
    InMux I__6340 (
            .O(N__35105),
            .I(N__35076));
    InMux I__6339 (
            .O(N__35104),
            .I(N__35076));
    CascadeMux I__6338 (
            .O(N__35103),
            .I(N__35071));
    CascadeMux I__6337 (
            .O(N__35102),
            .I(N__35068));
    InMux I__6336 (
            .O(N__35101),
            .I(N__35064));
    Span4Mux_v I__6335 (
            .O(N__35098),
            .I(N__35061));
    InMux I__6334 (
            .O(N__35097),
            .I(N__35054));
    InMux I__6333 (
            .O(N__35094),
            .I(N__35054));
    InMux I__6332 (
            .O(N__35093),
            .I(N__35054));
    CascadeMux I__6331 (
            .O(N__35092),
            .I(N__35049));
    InMux I__6330 (
            .O(N__35089),
            .I(N__35039));
    InMux I__6329 (
            .O(N__35086),
            .I(N__35039));
    InMux I__6328 (
            .O(N__35085),
            .I(N__35039));
    InMux I__6327 (
            .O(N__35084),
            .I(N__35034));
    InMux I__6326 (
            .O(N__35081),
            .I(N__35034));
    LocalMux I__6325 (
            .O(N__35076),
            .I(N__35031));
    InMux I__6324 (
            .O(N__35075),
            .I(N__35026));
    InMux I__6323 (
            .O(N__35074),
            .I(N__35026));
    InMux I__6322 (
            .O(N__35071),
            .I(N__35023));
    InMux I__6321 (
            .O(N__35068),
            .I(N__35018));
    InMux I__6320 (
            .O(N__35067),
            .I(N__35018));
    LocalMux I__6319 (
            .O(N__35064),
            .I(N__35015));
    Span4Mux_v I__6318 (
            .O(N__35061),
            .I(N__35010));
    LocalMux I__6317 (
            .O(N__35054),
            .I(N__35010));
    InMux I__6316 (
            .O(N__35053),
            .I(N__35007));
    InMux I__6315 (
            .O(N__35052),
            .I(N__35004));
    InMux I__6314 (
            .O(N__35049),
            .I(N__34997));
    InMux I__6313 (
            .O(N__35048),
            .I(N__34997));
    InMux I__6312 (
            .O(N__35047),
            .I(N__34997));
    InMux I__6311 (
            .O(N__35046),
            .I(N__34994));
    LocalMux I__6310 (
            .O(N__35039),
            .I(N__34989));
    LocalMux I__6309 (
            .O(N__35034),
            .I(N__34989));
    Span4Mux_v I__6308 (
            .O(N__35031),
            .I(N__34978));
    LocalMux I__6307 (
            .O(N__35026),
            .I(N__34978));
    LocalMux I__6306 (
            .O(N__35023),
            .I(N__34978));
    LocalMux I__6305 (
            .O(N__35018),
            .I(N__34978));
    Span4Mux_h I__6304 (
            .O(N__35015),
            .I(N__34978));
    Span4Mux_h I__6303 (
            .O(N__35010),
            .I(N__34975));
    LocalMux I__6302 (
            .O(N__35007),
            .I(n2445));
    LocalMux I__6301 (
            .O(N__35004),
            .I(n2445));
    LocalMux I__6300 (
            .O(N__34997),
            .I(n2445));
    LocalMux I__6299 (
            .O(N__34994),
            .I(n2445));
    Odrv4 I__6298 (
            .O(N__34989),
            .I(n2445));
    Odrv4 I__6297 (
            .O(N__34978),
            .I(n2445));
    Odrv4 I__6296 (
            .O(N__34975),
            .I(n2445));
    InMux I__6295 (
            .O(N__34960),
            .I(n12560));
    InMux I__6294 (
            .O(N__34957),
            .I(N__34954));
    LocalMux I__6293 (
            .O(N__34954),
            .I(N__34951));
    Span12Mux_h I__6292 (
            .O(N__34951),
            .I(N__34947));
    InMux I__6291 (
            .O(N__34950),
            .I(N__34944));
    Odrv12 I__6290 (
            .O(N__34947),
            .I(n15348));
    LocalMux I__6289 (
            .O(N__34944),
            .I(n15348));
    InMux I__6288 (
            .O(N__34939),
            .I(N__34936));
    LocalMux I__6287 (
            .O(N__34936),
            .I(N__34932));
    InMux I__6286 (
            .O(N__34935),
            .I(N__34921));
    Span4Mux_h I__6285 (
            .O(N__34932),
            .I(N__34916));
    InMux I__6284 (
            .O(N__34931),
            .I(N__34913));
    InMux I__6283 (
            .O(N__34930),
            .I(N__34910));
    InMux I__6282 (
            .O(N__34929),
            .I(N__34907));
    CascadeMux I__6281 (
            .O(N__34928),
            .I(N__34901));
    CascadeMux I__6280 (
            .O(N__34927),
            .I(N__34897));
    CascadeMux I__6279 (
            .O(N__34926),
            .I(N__34891));
    InMux I__6278 (
            .O(N__34925),
            .I(N__34885));
    InMux I__6277 (
            .O(N__34924),
            .I(N__34885));
    LocalMux I__6276 (
            .O(N__34921),
            .I(N__34882));
    InMux I__6275 (
            .O(N__34920),
            .I(N__34877));
    InMux I__6274 (
            .O(N__34919),
            .I(N__34877));
    Span4Mux_v I__6273 (
            .O(N__34916),
            .I(N__34872));
    LocalMux I__6272 (
            .O(N__34913),
            .I(N__34872));
    LocalMux I__6271 (
            .O(N__34910),
            .I(N__34869));
    LocalMux I__6270 (
            .O(N__34907),
            .I(N__34866));
    InMux I__6269 (
            .O(N__34906),
            .I(N__34861));
    InMux I__6268 (
            .O(N__34905),
            .I(N__34852));
    InMux I__6267 (
            .O(N__34904),
            .I(N__34852));
    InMux I__6266 (
            .O(N__34901),
            .I(N__34852));
    InMux I__6265 (
            .O(N__34900),
            .I(N__34852));
    InMux I__6264 (
            .O(N__34897),
            .I(N__34847));
    InMux I__6263 (
            .O(N__34896),
            .I(N__34847));
    InMux I__6262 (
            .O(N__34895),
            .I(N__34838));
    InMux I__6261 (
            .O(N__34894),
            .I(N__34838));
    InMux I__6260 (
            .O(N__34891),
            .I(N__34838));
    InMux I__6259 (
            .O(N__34890),
            .I(N__34838));
    LocalMux I__6258 (
            .O(N__34885),
            .I(N__34835));
    Span4Mux_s3_h I__6257 (
            .O(N__34882),
            .I(N__34830));
    LocalMux I__6256 (
            .O(N__34877),
            .I(N__34830));
    Span4Mux_h I__6255 (
            .O(N__34872),
            .I(N__34823));
    Span4Mux_h I__6254 (
            .O(N__34869),
            .I(N__34823));
    Span4Mux_s3_h I__6253 (
            .O(N__34866),
            .I(N__34823));
    InMux I__6252 (
            .O(N__34865),
            .I(N__34818));
    InMux I__6251 (
            .O(N__34864),
            .I(N__34818));
    LocalMux I__6250 (
            .O(N__34861),
            .I(n2346));
    LocalMux I__6249 (
            .O(N__34852),
            .I(n2346));
    LocalMux I__6248 (
            .O(N__34847),
            .I(n2346));
    LocalMux I__6247 (
            .O(N__34838),
            .I(n2346));
    Odrv4 I__6246 (
            .O(N__34835),
            .I(n2346));
    Odrv4 I__6245 (
            .O(N__34830),
            .I(n2346));
    Odrv4 I__6244 (
            .O(N__34823),
            .I(n2346));
    LocalMux I__6243 (
            .O(N__34818),
            .I(n2346));
    InMux I__6242 (
            .O(N__34801),
            .I(n12561));
    InMux I__6241 (
            .O(N__34798),
            .I(N__34795));
    LocalMux I__6240 (
            .O(N__34795),
            .I(N__34791));
    CascadeMux I__6239 (
            .O(N__34794),
            .I(N__34788));
    Span4Mux_v I__6238 (
            .O(N__34791),
            .I(N__34785));
    InMux I__6237 (
            .O(N__34788),
            .I(N__34782));
    Odrv4 I__6236 (
            .O(N__34785),
            .I(n15322));
    LocalMux I__6235 (
            .O(N__34782),
            .I(n15322));
    InMux I__6234 (
            .O(N__34777),
            .I(n12562));
    CascadeMux I__6233 (
            .O(N__34774),
            .I(n3138_cascade_));
    CascadeMux I__6232 (
            .O(N__34771),
            .I(n3229_cascade_));
    InMux I__6231 (
            .O(N__34768),
            .I(N__34765));
    LocalMux I__6230 (
            .O(N__34765),
            .I(n11658));
    InMux I__6229 (
            .O(N__34762),
            .I(bfn_9_25_0_));
    InMux I__6228 (
            .O(N__34759),
            .I(n12552));
    InMux I__6227 (
            .O(N__34756),
            .I(n12553));
    InMux I__6226 (
            .O(N__34753),
            .I(n12554));
    CascadeMux I__6225 (
            .O(N__34750),
            .I(n11750_cascade_));
    CascadeMux I__6224 (
            .O(N__34747),
            .I(n13900_cascade_));
    CascadeMux I__6223 (
            .O(N__34744),
            .I(n3232_cascade_));
    InMux I__6222 (
            .O(N__34741),
            .I(N__34738));
    LocalMux I__6221 (
            .O(N__34738),
            .I(n13906));
    CascadeMux I__6220 (
            .O(N__34735),
            .I(n13912_cascade_));
    InMux I__6219 (
            .O(N__34732),
            .I(n12381));
    InMux I__6218 (
            .O(N__34729),
            .I(n12382));
    InMux I__6217 (
            .O(N__34726),
            .I(n12383));
    InMux I__6216 (
            .O(N__34723),
            .I(n12384));
    InMux I__6215 (
            .O(N__34720),
            .I(bfn_9_22_0_));
    InMux I__6214 (
            .O(N__34717),
            .I(N__34712));
    InMux I__6213 (
            .O(N__34716),
            .I(N__34709));
    InMux I__6212 (
            .O(N__34715),
            .I(N__34706));
    LocalMux I__6211 (
            .O(N__34712),
            .I(N__34699));
    LocalMux I__6210 (
            .O(N__34709),
            .I(N__34699));
    LocalMux I__6209 (
            .O(N__34706),
            .I(N__34699));
    Span4Mux_v I__6208 (
            .O(N__34699),
            .I(N__34696));
    Odrv4 I__6207 (
            .O(N__34696),
            .I(n2622));
    InMux I__6206 (
            .O(N__34693),
            .I(N__34690));
    LocalMux I__6205 (
            .O(N__34690),
            .I(N__34687));
    Odrv4 I__6204 (
            .O(N__34687),
            .I(n2689));
    InMux I__6203 (
            .O(N__34684),
            .I(n12373));
    InMux I__6202 (
            .O(N__34681),
            .I(n12374));
    InMux I__6201 (
            .O(N__34678),
            .I(n12375));
    InMux I__6200 (
            .O(N__34675),
            .I(n12376));
    InMux I__6199 (
            .O(N__34672),
            .I(bfn_9_21_0_));
    InMux I__6198 (
            .O(N__34669),
            .I(n12378));
    InMux I__6197 (
            .O(N__34666),
            .I(n12379));
    InMux I__6196 (
            .O(N__34663),
            .I(n12380));
    InMux I__6195 (
            .O(N__34660),
            .I(n12364));
    InMux I__6194 (
            .O(N__34657),
            .I(n12365));
    InMux I__6193 (
            .O(N__34654),
            .I(n12366));
    InMux I__6192 (
            .O(N__34651),
            .I(n12367));
    InMux I__6191 (
            .O(N__34648),
            .I(n12368));
    InMux I__6190 (
            .O(N__34645),
            .I(bfn_9_20_0_));
    InMux I__6189 (
            .O(N__34642),
            .I(N__34639));
    LocalMux I__6188 (
            .O(N__34639),
            .I(N__34635));
    InMux I__6187 (
            .O(N__34638),
            .I(N__34632));
    Odrv4 I__6186 (
            .O(N__34635),
            .I(n2625));
    LocalMux I__6185 (
            .O(N__34632),
            .I(n2625));
    InMux I__6184 (
            .O(N__34627),
            .I(N__34624));
    LocalMux I__6183 (
            .O(N__34624),
            .I(N__34621));
    Odrv4 I__6182 (
            .O(N__34621),
            .I(n2692));
    InMux I__6181 (
            .O(N__34618),
            .I(n12370));
    InMux I__6180 (
            .O(N__34615),
            .I(n12371));
    InMux I__6179 (
            .O(N__34612),
            .I(n12372));
    CascadeMux I__6178 (
            .O(N__34609),
            .I(N__34605));
    InMux I__6177 (
            .O(N__34608),
            .I(N__34602));
    InMux I__6176 (
            .O(N__34605),
            .I(N__34599));
    LocalMux I__6175 (
            .O(N__34602),
            .I(N__34595));
    LocalMux I__6174 (
            .O(N__34599),
            .I(N__34592));
    InMux I__6173 (
            .O(N__34598),
            .I(N__34589));
    Span4Mux_v I__6172 (
            .O(N__34595),
            .I(N__34586));
    Span4Mux_v I__6171 (
            .O(N__34592),
            .I(N__34581));
    LocalMux I__6170 (
            .O(N__34589),
            .I(N__34581));
    Odrv4 I__6169 (
            .O(N__34586),
            .I(n2520));
    Odrv4 I__6168 (
            .O(N__34581),
            .I(n2520));
    CascadeMux I__6167 (
            .O(N__34576),
            .I(N__34573));
    InMux I__6166 (
            .O(N__34573),
            .I(N__34570));
    LocalMux I__6165 (
            .O(N__34570),
            .I(N__34567));
    Span4Mux_h I__6164 (
            .O(N__34567),
            .I(N__34564));
    Odrv4 I__6163 (
            .O(N__34564),
            .I(n2587));
    InMux I__6162 (
            .O(N__34561),
            .I(N__34558));
    LocalMux I__6161 (
            .O(N__34558),
            .I(N__34555));
    Span4Mux_h I__6160 (
            .O(N__34555),
            .I(N__34552));
    Odrv4 I__6159 (
            .O(N__34552),
            .I(n2580));
    InMux I__6158 (
            .O(N__34549),
            .I(N__34544));
    InMux I__6157 (
            .O(N__34548),
            .I(N__34541));
    InMux I__6156 (
            .O(N__34547),
            .I(N__34538));
    LocalMux I__6155 (
            .O(N__34544),
            .I(N__34533));
    LocalMux I__6154 (
            .O(N__34541),
            .I(N__34533));
    LocalMux I__6153 (
            .O(N__34538),
            .I(N__34530));
    Span4Mux_h I__6152 (
            .O(N__34533),
            .I(N__34527));
    Odrv12 I__6151 (
            .O(N__34530),
            .I(n2513));
    Odrv4 I__6150 (
            .O(N__34527),
            .I(n2513));
    CascadeMux I__6149 (
            .O(N__34522),
            .I(n2721_cascade_));
    InMux I__6148 (
            .O(N__34519),
            .I(N__34515));
    CascadeMux I__6147 (
            .O(N__34518),
            .I(N__34512));
    LocalMux I__6146 (
            .O(N__34515),
            .I(N__34508));
    InMux I__6145 (
            .O(N__34512),
            .I(N__34505));
    CascadeMux I__6144 (
            .O(N__34511),
            .I(N__34502));
    Span4Mux_h I__6143 (
            .O(N__34508),
            .I(N__34497));
    LocalMux I__6142 (
            .O(N__34505),
            .I(N__34497));
    InMux I__6141 (
            .O(N__34502),
            .I(N__34494));
    Odrv4 I__6140 (
            .O(N__34497),
            .I(n2526));
    LocalMux I__6139 (
            .O(N__34494),
            .I(n2526));
    CascadeMux I__6138 (
            .O(N__34489),
            .I(N__34486));
    InMux I__6137 (
            .O(N__34486),
            .I(N__34483));
    LocalMux I__6136 (
            .O(N__34483),
            .I(N__34480));
    Span4Mux_v I__6135 (
            .O(N__34480),
            .I(N__34477));
    Odrv4 I__6134 (
            .O(N__34477),
            .I(n2593));
    CascadeMux I__6133 (
            .O(N__34474),
            .I(n2625_cascade_));
    InMux I__6132 (
            .O(N__34471),
            .I(bfn_9_19_0_));
    InMux I__6131 (
            .O(N__34468),
            .I(n12362));
    InMux I__6130 (
            .O(N__34465),
            .I(n12363));
    InMux I__6129 (
            .O(N__34462),
            .I(N__34458));
    CascadeMux I__6128 (
            .O(N__34461),
            .I(N__34455));
    LocalMux I__6127 (
            .O(N__34458),
            .I(N__34452));
    InMux I__6126 (
            .O(N__34455),
            .I(N__34449));
    Span4Mux_h I__6125 (
            .O(N__34452),
            .I(N__34444));
    LocalMux I__6124 (
            .O(N__34449),
            .I(N__34444));
    Sp12to4 I__6123 (
            .O(N__34444),
            .I(N__34440));
    InMux I__6122 (
            .O(N__34443),
            .I(N__34437));
    Odrv12 I__6121 (
            .O(N__34440),
            .I(n2531));
    LocalMux I__6120 (
            .O(N__34437),
            .I(n2531));
    InMux I__6119 (
            .O(N__34432),
            .I(N__34429));
    LocalMux I__6118 (
            .O(N__34429),
            .I(N__34426));
    Span4Mux_h I__6117 (
            .O(N__34426),
            .I(N__34423));
    Odrv4 I__6116 (
            .O(N__34423),
            .I(n2598));
    CascadeMux I__6115 (
            .O(N__34420),
            .I(n2630_cascade_));
    CascadeMux I__6114 (
            .O(N__34417),
            .I(n14288_cascade_));
    CascadeMux I__6113 (
            .O(N__34414),
            .I(N__34410));
    InMux I__6112 (
            .O(N__34413),
            .I(N__34407));
    InMux I__6111 (
            .O(N__34410),
            .I(N__34404));
    LocalMux I__6110 (
            .O(N__34407),
            .I(N__34401));
    LocalMux I__6109 (
            .O(N__34404),
            .I(N__34398));
    Odrv12 I__6108 (
            .O(N__34401),
            .I(n2527));
    Odrv4 I__6107 (
            .O(N__34398),
            .I(n2527));
    CascadeMux I__6106 (
            .O(N__34393),
            .I(N__34390));
    InMux I__6105 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__6104 (
            .O(N__34387),
            .I(N__34384));
    Span4Mux_v I__6103 (
            .O(N__34384),
            .I(N__34381));
    Odrv4 I__6102 (
            .O(N__34381),
            .I(n2594));
    CascadeMux I__6101 (
            .O(N__34378),
            .I(n2626_cascade_));
    InMux I__6100 (
            .O(N__34375),
            .I(N__34372));
    LocalMux I__6099 (
            .O(N__34372),
            .I(N__34369));
    Odrv4 I__6098 (
            .O(N__34369),
            .I(n14278));
    CascadeMux I__6097 (
            .O(N__34366),
            .I(n14280_cascade_));
    InMux I__6096 (
            .O(N__34363),
            .I(N__34360));
    LocalMux I__6095 (
            .O(N__34360),
            .I(n14286));
    CascadeMux I__6094 (
            .O(N__34357),
            .I(N__34354));
    InMux I__6093 (
            .O(N__34354),
            .I(N__34350));
    CascadeMux I__6092 (
            .O(N__34353),
            .I(N__34347));
    LocalMux I__6091 (
            .O(N__34350),
            .I(N__34343));
    InMux I__6090 (
            .O(N__34347),
            .I(N__34340));
    InMux I__6089 (
            .O(N__34346),
            .I(N__34337));
    Span4Mux_h I__6088 (
            .O(N__34343),
            .I(N__34334));
    LocalMux I__6087 (
            .O(N__34340),
            .I(N__34331));
    LocalMux I__6086 (
            .O(N__34337),
            .I(N__34328));
    Odrv4 I__6085 (
            .O(N__34334),
            .I(n2522));
    Odrv4 I__6084 (
            .O(N__34331),
            .I(n2522));
    Odrv4 I__6083 (
            .O(N__34328),
            .I(n2522));
    InMux I__6082 (
            .O(N__34321),
            .I(N__34318));
    LocalMux I__6081 (
            .O(N__34318),
            .I(N__34315));
    Span4Mux_h I__6080 (
            .O(N__34315),
            .I(N__34312));
    Odrv4 I__6079 (
            .O(N__34312),
            .I(n2589));
    InMux I__6078 (
            .O(N__34309),
            .I(N__34306));
    LocalMux I__6077 (
            .O(N__34306),
            .I(N__34303));
    Span4Mux_v I__6076 (
            .O(N__34303),
            .I(N__34300));
    Odrv4 I__6075 (
            .O(N__34300),
            .I(n2597));
    CascadeMux I__6074 (
            .O(N__34297),
            .I(N__34293));
    InMux I__6073 (
            .O(N__34296),
            .I(N__34290));
    InMux I__6072 (
            .O(N__34293),
            .I(N__34287));
    LocalMux I__6071 (
            .O(N__34290),
            .I(N__34284));
    LocalMux I__6070 (
            .O(N__34287),
            .I(N__34281));
    Span4Mux_h I__6069 (
            .O(N__34284),
            .I(N__34277));
    Span4Mux_v I__6068 (
            .O(N__34281),
            .I(N__34274));
    InMux I__6067 (
            .O(N__34280),
            .I(N__34271));
    Odrv4 I__6066 (
            .O(N__34277),
            .I(n2530));
    Odrv4 I__6065 (
            .O(N__34274),
            .I(n2530));
    LocalMux I__6064 (
            .O(N__34271),
            .I(n2530));
    InMux I__6063 (
            .O(N__34264),
            .I(N__34261));
    LocalMux I__6062 (
            .O(N__34261),
            .I(N__34258));
    Odrv4 I__6061 (
            .O(N__34258),
            .I(n898));
    CascadeMux I__6060 (
            .O(N__34255),
            .I(N__34252));
    InMux I__6059 (
            .O(N__34252),
            .I(N__34247));
    CascadeMux I__6058 (
            .O(N__34251),
            .I(N__34244));
    CascadeMux I__6057 (
            .O(N__34250),
            .I(N__34241));
    LocalMux I__6056 (
            .O(N__34247),
            .I(N__34238));
    InMux I__6055 (
            .O(N__34244),
            .I(N__34235));
    InMux I__6054 (
            .O(N__34241),
            .I(N__34232));
    Odrv4 I__6053 (
            .O(N__34238),
            .I(n831));
    LocalMux I__6052 (
            .O(N__34235),
            .I(n831));
    LocalMux I__6051 (
            .O(N__34232),
            .I(n831));
    CascadeMux I__6050 (
            .O(N__34225),
            .I(N__34220));
    CascadeMux I__6049 (
            .O(N__34224),
            .I(N__34216));
    InMux I__6048 (
            .O(N__34223),
            .I(N__34211));
    InMux I__6047 (
            .O(N__34220),
            .I(N__34206));
    InMux I__6046 (
            .O(N__34219),
            .I(N__34206));
    InMux I__6045 (
            .O(N__34216),
            .I(N__34199));
    InMux I__6044 (
            .O(N__34215),
            .I(N__34199));
    InMux I__6043 (
            .O(N__34214),
            .I(N__34199));
    LocalMux I__6042 (
            .O(N__34211),
            .I(n861));
    LocalMux I__6041 (
            .O(N__34206),
            .I(n861));
    LocalMux I__6040 (
            .O(N__34199),
            .I(n861));
    CascadeMux I__6039 (
            .O(N__34192),
            .I(N__34188));
    CascadeMux I__6038 (
            .O(N__34191),
            .I(N__34185));
    InMux I__6037 (
            .O(N__34188),
            .I(N__34182));
    InMux I__6036 (
            .O(N__34185),
            .I(N__34179));
    LocalMux I__6035 (
            .O(N__34182),
            .I(n930));
    LocalMux I__6034 (
            .O(N__34179),
            .I(n930));
    CascadeMux I__6033 (
            .O(N__34174),
            .I(n930_cascade_));
    InMux I__6032 (
            .O(N__34171),
            .I(N__34167));
    CascadeMux I__6031 (
            .O(N__34170),
            .I(N__34164));
    LocalMux I__6030 (
            .O(N__34167),
            .I(N__34160));
    InMux I__6029 (
            .O(N__34164),
            .I(N__34157));
    InMux I__6028 (
            .O(N__34163),
            .I(N__34154));
    Odrv4 I__6027 (
            .O(N__34160),
            .I(n929));
    LocalMux I__6026 (
            .O(N__34157),
            .I(n929));
    LocalMux I__6025 (
            .O(N__34154),
            .I(n929));
    CascadeMux I__6024 (
            .O(N__34147),
            .I(N__34143));
    InMux I__6023 (
            .O(N__34146),
            .I(N__34140));
    InMux I__6022 (
            .O(N__34143),
            .I(N__34137));
    LocalMux I__6021 (
            .O(N__34140),
            .I(N__34134));
    LocalMux I__6020 (
            .O(N__34137),
            .I(n927));
    Odrv4 I__6019 (
            .O(N__34134),
            .I(n927));
    InMux I__6018 (
            .O(N__34129),
            .I(N__34125));
    CascadeMux I__6017 (
            .O(N__34128),
            .I(N__34122));
    LocalMux I__6016 (
            .O(N__34125),
            .I(N__34118));
    InMux I__6015 (
            .O(N__34122),
            .I(N__34115));
    InMux I__6014 (
            .O(N__34121),
            .I(N__34112));
    Odrv4 I__6013 (
            .O(N__34118),
            .I(n928));
    LocalMux I__6012 (
            .O(N__34115),
            .I(n928));
    LocalMux I__6011 (
            .O(N__34112),
            .I(n928));
    CascadeMux I__6010 (
            .O(N__34105),
            .I(n13726_cascade_));
    InMux I__6009 (
            .O(N__34102),
            .I(N__34099));
    LocalMux I__6008 (
            .O(N__34099),
            .I(n11710));
    InMux I__6007 (
            .O(N__34096),
            .I(N__34093));
    LocalMux I__6006 (
            .O(N__34093),
            .I(n1000));
    CascadeMux I__6005 (
            .O(N__34090),
            .I(n960_cascade_));
    CascadeMux I__6004 (
            .O(N__34087),
            .I(N__34083));
    InMux I__6003 (
            .O(N__34086),
            .I(N__34079));
    InMux I__6002 (
            .O(N__34083),
            .I(N__34076));
    InMux I__6001 (
            .O(N__34082),
            .I(N__34073));
    LocalMux I__6000 (
            .O(N__34079),
            .I(n933));
    LocalMux I__5999 (
            .O(N__34076),
            .I(n933));
    LocalMux I__5998 (
            .O(N__34073),
            .I(n933));
    InMux I__5997 (
            .O(N__34066),
            .I(N__34061));
    InMux I__5996 (
            .O(N__34065),
            .I(N__34058));
    InMux I__5995 (
            .O(N__34064),
            .I(N__34055));
    LocalMux I__5994 (
            .O(N__34061),
            .I(n295));
    LocalMux I__5993 (
            .O(N__34058),
            .I(n295));
    LocalMux I__5992 (
            .O(N__34055),
            .I(n295));
    CascadeMux I__5991 (
            .O(N__34048),
            .I(N__34045));
    InMux I__5990 (
            .O(N__34045),
            .I(N__34042));
    LocalMux I__5989 (
            .O(N__34042),
            .I(n1001));
    CascadeMux I__5988 (
            .O(N__34039),
            .I(N__34035));
    InMux I__5987 (
            .O(N__34038),
            .I(N__34031));
    InMux I__5986 (
            .O(N__34035),
            .I(N__34028));
    InMux I__5985 (
            .O(N__34034),
            .I(N__34025));
    LocalMux I__5984 (
            .O(N__34031),
            .I(n931));
    LocalMux I__5983 (
            .O(N__34028),
            .I(n931));
    LocalMux I__5982 (
            .O(N__34025),
            .I(n931));
    InMux I__5981 (
            .O(N__34018),
            .I(N__34011));
    CascadeMux I__5980 (
            .O(N__34017),
            .I(N__34008));
    CascadeMux I__5979 (
            .O(N__34016),
            .I(N__34005));
    InMux I__5978 (
            .O(N__34015),
            .I(N__34000));
    InMux I__5977 (
            .O(N__34014),
            .I(N__33997));
    LocalMux I__5976 (
            .O(N__34011),
            .I(N__33994));
    InMux I__5975 (
            .O(N__34008),
            .I(N__33985));
    InMux I__5974 (
            .O(N__34005),
            .I(N__33985));
    InMux I__5973 (
            .O(N__34004),
            .I(N__33985));
    InMux I__5972 (
            .O(N__34003),
            .I(N__33985));
    LocalMux I__5971 (
            .O(N__34000),
            .I(n960));
    LocalMux I__5970 (
            .O(N__33997),
            .I(n960));
    Odrv4 I__5969 (
            .O(N__33994),
            .I(n960));
    LocalMux I__5968 (
            .O(N__33985),
            .I(n960));
    InMux I__5967 (
            .O(N__33976),
            .I(N__33973));
    LocalMux I__5966 (
            .O(N__33973),
            .I(n998));
    CascadeMux I__5965 (
            .O(N__33970),
            .I(N__33966));
    InMux I__5964 (
            .O(N__33969),
            .I(N__33962));
    InMux I__5963 (
            .O(N__33966),
            .I(N__33959));
    InMux I__5962 (
            .O(N__33965),
            .I(N__33956));
    LocalMux I__5961 (
            .O(N__33962),
            .I(n1032));
    LocalMux I__5960 (
            .O(N__33959),
            .I(n1032));
    LocalMux I__5959 (
            .O(N__33956),
            .I(n1032));
    CascadeMux I__5958 (
            .O(N__33949),
            .I(N__33944));
    InMux I__5957 (
            .O(N__33948),
            .I(N__33941));
    InMux I__5956 (
            .O(N__33947),
            .I(N__33938));
    InMux I__5955 (
            .O(N__33944),
            .I(N__33935));
    LocalMux I__5954 (
            .O(N__33941),
            .I(n296));
    LocalMux I__5953 (
            .O(N__33938),
            .I(n296));
    LocalMux I__5952 (
            .O(N__33935),
            .I(n296));
    InMux I__5951 (
            .O(N__33928),
            .I(N__33924));
    CascadeMux I__5950 (
            .O(N__33927),
            .I(N__33921));
    LocalMux I__5949 (
            .O(N__33924),
            .I(N__33917));
    InMux I__5948 (
            .O(N__33921),
            .I(N__33914));
    InMux I__5947 (
            .O(N__33920),
            .I(N__33911));
    Odrv4 I__5946 (
            .O(N__33917),
            .I(n1033));
    LocalMux I__5945 (
            .O(N__33914),
            .I(n1033));
    LocalMux I__5944 (
            .O(N__33911),
            .I(n1033));
    CascadeMux I__5943 (
            .O(N__33904),
            .I(N__33901));
    InMux I__5942 (
            .O(N__33901),
            .I(N__33898));
    LocalMux I__5941 (
            .O(N__33898),
            .I(N__33894));
    CascadeMux I__5940 (
            .O(N__33897),
            .I(N__33891));
    Span4Mux_s1_v I__5939 (
            .O(N__33894),
            .I(N__33887));
    InMux I__5938 (
            .O(N__33891),
            .I(N__33884));
    InMux I__5937 (
            .O(N__33890),
            .I(N__33881));
    Odrv4 I__5936 (
            .O(N__33887),
            .I(n1031));
    LocalMux I__5935 (
            .O(N__33884),
            .I(n1031));
    LocalMux I__5934 (
            .O(N__33881),
            .I(n1031));
    CascadeMux I__5933 (
            .O(N__33874),
            .I(N__33870));
    InMux I__5932 (
            .O(N__33873),
            .I(N__33866));
    InMux I__5931 (
            .O(N__33870),
            .I(N__33863));
    InMux I__5930 (
            .O(N__33869),
            .I(N__33860));
    LocalMux I__5929 (
            .O(N__33866),
            .I(n1029));
    LocalMux I__5928 (
            .O(N__33863),
            .I(n1029));
    LocalMux I__5927 (
            .O(N__33860),
            .I(n1029));
    CascadeMux I__5926 (
            .O(N__33853),
            .I(n11646_cascade_));
    InMux I__5925 (
            .O(N__33850),
            .I(N__33846));
    CascadeMux I__5924 (
            .O(N__33849),
            .I(N__33843));
    LocalMux I__5923 (
            .O(N__33846),
            .I(N__33839));
    InMux I__5922 (
            .O(N__33843),
            .I(N__33836));
    InMux I__5921 (
            .O(N__33842),
            .I(N__33833));
    Odrv12 I__5920 (
            .O(N__33839),
            .I(n1030));
    LocalMux I__5919 (
            .O(N__33836),
            .I(n1030));
    LocalMux I__5918 (
            .O(N__33833),
            .I(n1030));
    InMux I__5917 (
            .O(N__33826),
            .I(N__33823));
    LocalMux I__5916 (
            .O(N__33823),
            .I(n13323));
    InMux I__5915 (
            .O(N__33820),
            .I(n12107));
    InMux I__5914 (
            .O(N__33817),
            .I(n12108));
    InMux I__5913 (
            .O(N__33814),
            .I(n12109));
    InMux I__5912 (
            .O(N__33811),
            .I(n12110));
    CascadeMux I__5911 (
            .O(N__33808),
            .I(N__33805));
    InMux I__5910 (
            .O(N__33805),
            .I(N__33802));
    LocalMux I__5909 (
            .O(N__33802),
            .I(N__33799));
    Odrv4 I__5908 (
            .O(N__33799),
            .I(n996));
    InMux I__5907 (
            .O(N__33796),
            .I(n12111));
    CascadeMux I__5906 (
            .O(N__33793),
            .I(N__33790));
    InMux I__5905 (
            .O(N__33790),
            .I(N__33787));
    LocalMux I__5904 (
            .O(N__33787),
            .I(n995));
    InMux I__5903 (
            .O(N__33784),
            .I(n12112));
    InMux I__5902 (
            .O(N__33781),
            .I(n12113));
    CascadeMux I__5901 (
            .O(N__33778),
            .I(N__33775));
    InMux I__5900 (
            .O(N__33775),
            .I(N__33772));
    LocalMux I__5899 (
            .O(N__33772),
            .I(N__33767));
    InMux I__5898 (
            .O(N__33771),
            .I(N__33762));
    InMux I__5897 (
            .O(N__33770),
            .I(N__33762));
    Span4Mux_s2_v I__5896 (
            .O(N__33767),
            .I(N__33759));
    LocalMux I__5895 (
            .O(N__33762),
            .I(N__33756));
    Odrv4 I__5894 (
            .O(N__33759),
            .I(n1026));
    Odrv4 I__5893 (
            .O(N__33756),
            .I(n1026));
    InMux I__5892 (
            .O(N__33751),
            .I(N__33748));
    LocalMux I__5891 (
            .O(N__33748),
            .I(n997));
    InMux I__5890 (
            .O(N__33745),
            .I(N__33742));
    LocalMux I__5889 (
            .O(N__33742),
            .I(n999));
    InMux I__5888 (
            .O(N__33739),
            .I(N__33734));
    CascadeMux I__5887 (
            .O(N__33738),
            .I(N__33731));
    CascadeMux I__5886 (
            .O(N__33737),
            .I(N__33728));
    LocalMux I__5885 (
            .O(N__33734),
            .I(N__33725));
    InMux I__5884 (
            .O(N__33731),
            .I(N__33722));
    InMux I__5883 (
            .O(N__33728),
            .I(N__33719));
    Odrv4 I__5882 (
            .O(N__33725),
            .I(n932));
    LocalMux I__5881 (
            .O(N__33722),
            .I(n932));
    LocalMux I__5880 (
            .O(N__33719),
            .I(n932));
    InMux I__5879 (
            .O(N__33712),
            .I(n12101));
    CascadeMux I__5878 (
            .O(N__33709),
            .I(N__33704));
    InMux I__5877 (
            .O(N__33708),
            .I(N__33699));
    InMux I__5876 (
            .O(N__33707),
            .I(N__33699));
    InMux I__5875 (
            .O(N__33704),
            .I(N__33696));
    LocalMux I__5874 (
            .O(N__33699),
            .I(N__33693));
    LocalMux I__5873 (
            .O(N__33696),
            .I(N__33690));
    Span4Mux_s3_v I__5872 (
            .O(N__33693),
            .I(N__33687));
    Span4Mux_h I__5871 (
            .O(N__33690),
            .I(N__33684));
    Odrv4 I__5870 (
            .O(N__33687),
            .I(n832));
    Odrv4 I__5869 (
            .O(N__33684),
            .I(n832));
    CascadeMux I__5868 (
            .O(N__33679),
            .I(N__33676));
    InMux I__5867 (
            .O(N__33676),
            .I(N__33673));
    LocalMux I__5866 (
            .O(N__33673),
            .I(n899));
    InMux I__5865 (
            .O(N__33670),
            .I(n12102));
    InMux I__5864 (
            .O(N__33667),
            .I(n12103));
    CascadeMux I__5863 (
            .O(N__33664),
            .I(N__33661));
    InMux I__5862 (
            .O(N__33661),
            .I(N__33658));
    LocalMux I__5861 (
            .O(N__33658),
            .I(N__33653));
    InMux I__5860 (
            .O(N__33657),
            .I(N__33648));
    InMux I__5859 (
            .O(N__33656),
            .I(N__33648));
    Span4Mux_v I__5858 (
            .O(N__33653),
            .I(N__33645));
    LocalMux I__5857 (
            .O(N__33648),
            .I(N__33642));
    Odrv4 I__5856 (
            .O(N__33645),
            .I(n830));
    Odrv4 I__5855 (
            .O(N__33642),
            .I(n830));
    CascadeMux I__5854 (
            .O(N__33637),
            .I(N__33634));
    InMux I__5853 (
            .O(N__33634),
            .I(N__33631));
    LocalMux I__5852 (
            .O(N__33631),
            .I(n897));
    InMux I__5851 (
            .O(N__33628),
            .I(n12104));
    CascadeMux I__5850 (
            .O(N__33625),
            .I(N__33622));
    InMux I__5849 (
            .O(N__33622),
            .I(N__33617));
    InMux I__5848 (
            .O(N__33621),
            .I(N__33612));
    InMux I__5847 (
            .O(N__33620),
            .I(N__33612));
    LocalMux I__5846 (
            .O(N__33617),
            .I(n829));
    LocalMux I__5845 (
            .O(N__33612),
            .I(n829));
    InMux I__5844 (
            .O(N__33607),
            .I(N__33604));
    LocalMux I__5843 (
            .O(N__33604),
            .I(n896));
    InMux I__5842 (
            .O(N__33601),
            .I(n12105));
    InMux I__5841 (
            .O(N__33598),
            .I(N__33594));
    InMux I__5840 (
            .O(N__33597),
            .I(N__33591));
    LocalMux I__5839 (
            .O(N__33594),
            .I(N__33588));
    LocalMux I__5838 (
            .O(N__33591),
            .I(n828));
    Odrv4 I__5837 (
            .O(N__33588),
            .I(n828));
    InMux I__5836 (
            .O(N__33583),
            .I(n12106));
    InMux I__5835 (
            .O(N__33580),
            .I(N__33577));
    LocalMux I__5834 (
            .O(N__33577),
            .I(n900));
    CascadeMux I__5833 (
            .O(N__33574),
            .I(N__33569));
    CascadeMux I__5832 (
            .O(N__33573),
            .I(N__33566));
    InMux I__5831 (
            .O(N__33572),
            .I(N__33563));
    InMux I__5830 (
            .O(N__33569),
            .I(N__33558));
    InMux I__5829 (
            .O(N__33566),
            .I(N__33558));
    LocalMux I__5828 (
            .O(N__33563),
            .I(n833));
    LocalMux I__5827 (
            .O(N__33558),
            .I(n833));
    InMux I__5826 (
            .O(N__33553),
            .I(bfn_7_30_0_));
    CascadeMux I__5825 (
            .O(N__33550),
            .I(N__33547));
    InMux I__5824 (
            .O(N__33547),
            .I(N__33544));
    LocalMux I__5823 (
            .O(N__33544),
            .I(N__33541));
    Span4Mux_h I__5822 (
            .O(N__33541),
            .I(N__33538));
    Odrv4 I__5821 (
            .O(N__33538),
            .I(n8_adj_632));
    InMux I__5820 (
            .O(N__33535),
            .I(n12599));
    CascadeMux I__5819 (
            .O(N__33532),
            .I(N__33529));
    InMux I__5818 (
            .O(N__33529),
            .I(N__33526));
    LocalMux I__5817 (
            .O(N__33526),
            .I(n7_adj_631));
    InMux I__5816 (
            .O(N__33523),
            .I(N__33517));
    InMux I__5815 (
            .O(N__33522),
            .I(N__33517));
    LocalMux I__5814 (
            .O(N__33517),
            .I(n7));
    InMux I__5813 (
            .O(N__33514),
            .I(n12600));
    CascadeMux I__5812 (
            .O(N__33511),
            .I(N__33508));
    InMux I__5811 (
            .O(N__33508),
            .I(N__33505));
    LocalMux I__5810 (
            .O(N__33505),
            .I(N__33502));
    Span4Mux_h I__5809 (
            .O(N__33502),
            .I(N__33499));
    Odrv4 I__5808 (
            .O(N__33499),
            .I(n6_adj_630));
    InMux I__5807 (
            .O(N__33496),
            .I(N__33493));
    LocalMux I__5806 (
            .O(N__33493),
            .I(N__33488));
    InMux I__5805 (
            .O(N__33492),
            .I(N__33485));
    InMux I__5804 (
            .O(N__33491),
            .I(N__33482));
    Odrv4 I__5803 (
            .O(N__33488),
            .I(n6));
    LocalMux I__5802 (
            .O(N__33485),
            .I(n6));
    LocalMux I__5801 (
            .O(N__33482),
            .I(n6));
    InMux I__5800 (
            .O(N__33475),
            .I(n12601));
    CascadeMux I__5799 (
            .O(N__33472),
            .I(N__33469));
    InMux I__5798 (
            .O(N__33469),
            .I(N__33466));
    LocalMux I__5797 (
            .O(N__33466),
            .I(N__33463));
    Span4Mux_v I__5796 (
            .O(N__33463),
            .I(N__33458));
    InMux I__5795 (
            .O(N__33462),
            .I(N__33455));
    InMux I__5794 (
            .O(N__33461),
            .I(N__33452));
    Odrv4 I__5793 (
            .O(N__33458),
            .I(n5));
    LocalMux I__5792 (
            .O(N__33455),
            .I(n5));
    LocalMux I__5791 (
            .O(N__33452),
            .I(n5));
    InMux I__5790 (
            .O(N__33445),
            .I(n12602));
    CascadeMux I__5789 (
            .O(N__33442),
            .I(N__33439));
    InMux I__5788 (
            .O(N__33439),
            .I(N__33436));
    LocalMux I__5787 (
            .O(N__33436),
            .I(N__33433));
    Span4Mux_h I__5786 (
            .O(N__33433),
            .I(N__33430));
    Odrv4 I__5785 (
            .O(N__33430),
            .I(n4_adj_628));
    InMux I__5784 (
            .O(N__33427),
            .I(N__33424));
    LocalMux I__5783 (
            .O(N__33424),
            .I(N__33421));
    Span4Mux_h I__5782 (
            .O(N__33421),
            .I(N__33416));
    InMux I__5781 (
            .O(N__33420),
            .I(N__33411));
    InMux I__5780 (
            .O(N__33419),
            .I(N__33411));
    Odrv4 I__5779 (
            .O(N__33416),
            .I(n4));
    LocalMux I__5778 (
            .O(N__33411),
            .I(n4));
    InMux I__5777 (
            .O(N__33406),
            .I(n12603));
    CascadeMux I__5776 (
            .O(N__33403),
            .I(N__33400));
    InMux I__5775 (
            .O(N__33400),
            .I(N__33397));
    LocalMux I__5774 (
            .O(N__33397),
            .I(n3_adj_627));
    CascadeMux I__5773 (
            .O(N__33394),
            .I(N__33389));
    InMux I__5772 (
            .O(N__33393),
            .I(N__33383));
    InMux I__5771 (
            .O(N__33392),
            .I(N__33383));
    InMux I__5770 (
            .O(N__33389),
            .I(N__33378));
    InMux I__5769 (
            .O(N__33388),
            .I(N__33378));
    LocalMux I__5768 (
            .O(N__33383),
            .I(n3_adj_567));
    LocalMux I__5767 (
            .O(N__33378),
            .I(n3_adj_567));
    InMux I__5766 (
            .O(N__33373),
            .I(n12604));
    InMux I__5765 (
            .O(N__33370),
            .I(n12605));
    InMux I__5764 (
            .O(N__33367),
            .I(N__33364));
    LocalMux I__5763 (
            .O(N__33364),
            .I(N__33359));
    InMux I__5762 (
            .O(N__33363),
            .I(N__33354));
    InMux I__5761 (
            .O(N__33362),
            .I(N__33354));
    Span4Mux_h I__5760 (
            .O(N__33359),
            .I(N__33351));
    LocalMux I__5759 (
            .O(N__33354),
            .I(n2_adj_568));
    Odrv4 I__5758 (
            .O(N__33351),
            .I(n2_adj_568));
    InMux I__5757 (
            .O(N__33346),
            .I(N__33343));
    LocalMux I__5756 (
            .O(N__33343),
            .I(n901));
    InMux I__5755 (
            .O(N__33340),
            .I(bfn_7_29_0_));
    CascadeMux I__5754 (
            .O(N__33337),
            .I(N__33334));
    InMux I__5753 (
            .O(N__33334),
            .I(N__33331));
    LocalMux I__5752 (
            .O(N__33331),
            .I(N__33328));
    Odrv4 I__5751 (
            .O(N__33328),
            .I(n16_adj_640));
    InMux I__5750 (
            .O(N__33325),
            .I(N__33322));
    LocalMux I__5749 (
            .O(N__33322),
            .I(N__33319));
    Odrv4 I__5748 (
            .O(N__33319),
            .I(n16));
    InMux I__5747 (
            .O(N__33316),
            .I(n12591));
    CascadeMux I__5746 (
            .O(N__33313),
            .I(N__33310));
    InMux I__5745 (
            .O(N__33310),
            .I(N__33307));
    LocalMux I__5744 (
            .O(N__33307),
            .I(N__33304));
    Odrv4 I__5743 (
            .O(N__33304),
            .I(n15_adj_639));
    InMux I__5742 (
            .O(N__33301),
            .I(N__33298));
    LocalMux I__5741 (
            .O(N__33298),
            .I(N__33295));
    Span4Mux_v I__5740 (
            .O(N__33295),
            .I(N__33292));
    Span4Mux_h I__5739 (
            .O(N__33292),
            .I(N__33289));
    Odrv4 I__5738 (
            .O(N__33289),
            .I(n15));
    InMux I__5737 (
            .O(N__33286),
            .I(n12592));
    CascadeMux I__5736 (
            .O(N__33283),
            .I(N__33280));
    InMux I__5735 (
            .O(N__33280),
            .I(N__33277));
    LocalMux I__5734 (
            .O(N__33277),
            .I(N__33274));
    Odrv12 I__5733 (
            .O(N__33274),
            .I(n14_adj_638));
    InMux I__5732 (
            .O(N__33271),
            .I(N__33268));
    LocalMux I__5731 (
            .O(N__33268),
            .I(N__33265));
    Odrv12 I__5730 (
            .O(N__33265),
            .I(n14));
    InMux I__5729 (
            .O(N__33262),
            .I(n12593));
    CascadeMux I__5728 (
            .O(N__33259),
            .I(N__33256));
    InMux I__5727 (
            .O(N__33256),
            .I(N__33253));
    LocalMux I__5726 (
            .O(N__33253),
            .I(N__33250));
    Span4Mux_h I__5725 (
            .O(N__33250),
            .I(N__33247));
    Odrv4 I__5724 (
            .O(N__33247),
            .I(n13_adj_637));
    InMux I__5723 (
            .O(N__33244),
            .I(N__33241));
    LocalMux I__5722 (
            .O(N__33241),
            .I(N__33238));
    Span4Mux_h I__5721 (
            .O(N__33238),
            .I(N__33235));
    Odrv4 I__5720 (
            .O(N__33235),
            .I(n13));
    InMux I__5719 (
            .O(N__33232),
            .I(n12594));
    CascadeMux I__5718 (
            .O(N__33229),
            .I(N__33226));
    InMux I__5717 (
            .O(N__33226),
            .I(N__33223));
    LocalMux I__5716 (
            .O(N__33223),
            .I(N__33220));
    Span4Mux_h I__5715 (
            .O(N__33220),
            .I(N__33217));
    Odrv4 I__5714 (
            .O(N__33217),
            .I(n12_adj_636));
    InMux I__5713 (
            .O(N__33214),
            .I(N__33211));
    LocalMux I__5712 (
            .O(N__33211),
            .I(N__33208));
    Span4Mux_h I__5711 (
            .O(N__33208),
            .I(N__33205));
    Odrv4 I__5710 (
            .O(N__33205),
            .I(n12));
    InMux I__5709 (
            .O(N__33202),
            .I(n12595));
    CascadeMux I__5708 (
            .O(N__33199),
            .I(N__33196));
    InMux I__5707 (
            .O(N__33196),
            .I(N__33193));
    LocalMux I__5706 (
            .O(N__33193),
            .I(N__33190));
    Span4Mux_h I__5705 (
            .O(N__33190),
            .I(N__33187));
    Odrv4 I__5704 (
            .O(N__33187),
            .I(n11_adj_635));
    InMux I__5703 (
            .O(N__33184),
            .I(N__33181));
    LocalMux I__5702 (
            .O(N__33181),
            .I(N__33178));
    Span4Mux_h I__5701 (
            .O(N__33178),
            .I(N__33175));
    Odrv4 I__5700 (
            .O(N__33175),
            .I(n11));
    InMux I__5699 (
            .O(N__33172),
            .I(n12596));
    CascadeMux I__5698 (
            .O(N__33169),
            .I(N__33166));
    InMux I__5697 (
            .O(N__33166),
            .I(N__33163));
    LocalMux I__5696 (
            .O(N__33163),
            .I(N__33160));
    Span4Mux_h I__5695 (
            .O(N__33160),
            .I(N__33157));
    Span4Mux_v I__5694 (
            .O(N__33157),
            .I(N__33154));
    Odrv4 I__5693 (
            .O(N__33154),
            .I(n10_adj_634));
    CascadeMux I__5692 (
            .O(N__33151),
            .I(N__33148));
    InMux I__5691 (
            .O(N__33148),
            .I(N__33145));
    LocalMux I__5690 (
            .O(N__33145),
            .I(N__33142));
    Span4Mux_s2_v I__5689 (
            .O(N__33142),
            .I(N__33139));
    Odrv4 I__5688 (
            .O(N__33139),
            .I(n10));
    InMux I__5687 (
            .O(N__33136),
            .I(n12597));
    CascadeMux I__5686 (
            .O(N__33133),
            .I(N__33130));
    InMux I__5685 (
            .O(N__33130),
            .I(N__33127));
    LocalMux I__5684 (
            .O(N__33127),
            .I(N__33124));
    Span4Mux_v I__5683 (
            .O(N__33124),
            .I(N__33121));
    Odrv4 I__5682 (
            .O(N__33121),
            .I(n9_adj_633));
    CascadeMux I__5681 (
            .O(N__33118),
            .I(N__33115));
    InMux I__5680 (
            .O(N__33115),
            .I(N__33112));
    LocalMux I__5679 (
            .O(N__33112),
            .I(N__33109));
    Odrv4 I__5678 (
            .O(N__33109),
            .I(n9));
    InMux I__5677 (
            .O(N__33106),
            .I(bfn_7_28_0_));
    CascadeMux I__5676 (
            .O(N__33103),
            .I(N__33100));
    InMux I__5675 (
            .O(N__33100),
            .I(N__33097));
    LocalMux I__5674 (
            .O(N__33097),
            .I(n24_adj_648));
    InMux I__5673 (
            .O(N__33094),
            .I(n12583));
    CascadeMux I__5672 (
            .O(N__33091),
            .I(N__33088));
    InMux I__5671 (
            .O(N__33088),
            .I(N__33085));
    LocalMux I__5670 (
            .O(N__33085),
            .I(N__33082));
    Span12Mux_v I__5669 (
            .O(N__33082),
            .I(N__33079));
    Odrv12 I__5668 (
            .O(N__33079),
            .I(n23_adj_647));
    InMux I__5667 (
            .O(N__33076),
            .I(n12584));
    CascadeMux I__5666 (
            .O(N__33073),
            .I(N__33070));
    InMux I__5665 (
            .O(N__33070),
            .I(N__33067));
    LocalMux I__5664 (
            .O(N__33067),
            .I(N__33064));
    Odrv4 I__5663 (
            .O(N__33064),
            .I(n22_adj_646));
    InMux I__5662 (
            .O(N__33061),
            .I(N__33058));
    LocalMux I__5661 (
            .O(N__33058),
            .I(N__33055));
    Odrv4 I__5660 (
            .O(N__33055),
            .I(n22));
    InMux I__5659 (
            .O(N__33052),
            .I(n12585));
    CascadeMux I__5658 (
            .O(N__33049),
            .I(N__33046));
    InMux I__5657 (
            .O(N__33046),
            .I(N__33043));
    LocalMux I__5656 (
            .O(N__33043),
            .I(N__33040));
    Span4Mux_h I__5655 (
            .O(N__33040),
            .I(N__33037));
    Odrv4 I__5654 (
            .O(N__33037),
            .I(n21_adj_645));
    InMux I__5653 (
            .O(N__33034),
            .I(N__33031));
    LocalMux I__5652 (
            .O(N__33031),
            .I(N__33028));
    Odrv4 I__5651 (
            .O(N__33028),
            .I(n21));
    InMux I__5650 (
            .O(N__33025),
            .I(n12586));
    InMux I__5649 (
            .O(N__33022),
            .I(N__33019));
    LocalMux I__5648 (
            .O(N__33019),
            .I(N__33016));
    Odrv4 I__5647 (
            .O(N__33016),
            .I(n20));
    InMux I__5646 (
            .O(N__33013),
            .I(n12587));
    InMux I__5645 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__5644 (
            .O(N__33007),
            .I(n19_adj_643));
    InMux I__5643 (
            .O(N__33004),
            .I(n12588));
    CascadeMux I__5642 (
            .O(N__33001),
            .I(N__32998));
    InMux I__5641 (
            .O(N__32998),
            .I(N__32995));
    LocalMux I__5640 (
            .O(N__32995),
            .I(n18_adj_642));
    InMux I__5639 (
            .O(N__32992),
            .I(N__32989));
    LocalMux I__5638 (
            .O(N__32989),
            .I(N__32986));
    Odrv4 I__5637 (
            .O(N__32986),
            .I(n18));
    InMux I__5636 (
            .O(N__32983),
            .I(n12589));
    CascadeMux I__5635 (
            .O(N__32980),
            .I(N__32977));
    InMux I__5634 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__5633 (
            .O(N__32974),
            .I(n17_adj_641));
    InMux I__5632 (
            .O(N__32971),
            .I(N__32968));
    LocalMux I__5631 (
            .O(N__32968),
            .I(N__32965));
    Span4Mux_h I__5630 (
            .O(N__32965),
            .I(N__32962));
    Odrv4 I__5629 (
            .O(N__32962),
            .I(n17));
    InMux I__5628 (
            .O(N__32959),
            .I(bfn_7_27_0_));
    CascadeMux I__5627 (
            .O(N__32956),
            .I(N__32953));
    InMux I__5626 (
            .O(N__32953),
            .I(N__32950));
    LocalMux I__5625 (
            .O(N__32950),
            .I(n32_adj_656));
    InMux I__5624 (
            .O(N__32947),
            .I(N__32944));
    LocalMux I__5623 (
            .O(N__32944),
            .I(n32));
    InMux I__5622 (
            .O(N__32941),
            .I(n12575));
    InMux I__5621 (
            .O(N__32938),
            .I(N__32935));
    LocalMux I__5620 (
            .O(N__32935),
            .I(N__32932));
    Odrv4 I__5619 (
            .O(N__32932),
            .I(n31_adj_655));
    InMux I__5618 (
            .O(N__32929),
            .I(N__32926));
    LocalMux I__5617 (
            .O(N__32926),
            .I(N__32923));
    Span4Mux_v I__5616 (
            .O(N__32923),
            .I(N__32920));
    Span4Mux_h I__5615 (
            .O(N__32920),
            .I(N__32917));
    Odrv4 I__5614 (
            .O(N__32917),
            .I(n31));
    InMux I__5613 (
            .O(N__32914),
            .I(n12576));
    CascadeMux I__5612 (
            .O(N__32911),
            .I(N__32908));
    InMux I__5611 (
            .O(N__32908),
            .I(N__32905));
    LocalMux I__5610 (
            .O(N__32905),
            .I(N__32902));
    Span4Mux_h I__5609 (
            .O(N__32902),
            .I(N__32899));
    Odrv4 I__5608 (
            .O(N__32899),
            .I(n30_adj_654));
    InMux I__5607 (
            .O(N__32896),
            .I(N__32893));
    LocalMux I__5606 (
            .O(N__32893),
            .I(N__32890));
    Odrv4 I__5605 (
            .O(N__32890),
            .I(n30));
    InMux I__5604 (
            .O(N__32887),
            .I(n12577));
    CascadeMux I__5603 (
            .O(N__32884),
            .I(N__32881));
    InMux I__5602 (
            .O(N__32881),
            .I(N__32878));
    LocalMux I__5601 (
            .O(N__32878),
            .I(N__32875));
    Odrv4 I__5600 (
            .O(N__32875),
            .I(n29_adj_653));
    InMux I__5599 (
            .O(N__32872),
            .I(n12578));
    CascadeMux I__5598 (
            .O(N__32869),
            .I(N__32866));
    InMux I__5597 (
            .O(N__32866),
            .I(N__32863));
    LocalMux I__5596 (
            .O(N__32863),
            .I(n28_adj_652));
    InMux I__5595 (
            .O(N__32860),
            .I(N__32857));
    LocalMux I__5594 (
            .O(N__32857),
            .I(N__32854));
    Span4Mux_h I__5593 (
            .O(N__32854),
            .I(N__32851));
    Odrv4 I__5592 (
            .O(N__32851),
            .I(n28));
    InMux I__5591 (
            .O(N__32848),
            .I(n12579));
    InMux I__5590 (
            .O(N__32845),
            .I(N__32842));
    LocalMux I__5589 (
            .O(N__32842),
            .I(N__32839));
    Odrv12 I__5588 (
            .O(N__32839),
            .I(n27));
    InMux I__5587 (
            .O(N__32836),
            .I(n12580));
    CascadeMux I__5586 (
            .O(N__32833),
            .I(N__32830));
    InMux I__5585 (
            .O(N__32830),
            .I(N__32827));
    LocalMux I__5584 (
            .O(N__32827),
            .I(n26_adj_650));
    InMux I__5583 (
            .O(N__32824),
            .I(n12581));
    CascadeMux I__5582 (
            .O(N__32821),
            .I(N__32818));
    InMux I__5581 (
            .O(N__32818),
            .I(N__32815));
    LocalMux I__5580 (
            .O(N__32815),
            .I(n25_adj_649));
    InMux I__5579 (
            .O(N__32812),
            .I(N__32809));
    LocalMux I__5578 (
            .O(N__32809),
            .I(N__32806));
    Odrv4 I__5577 (
            .O(N__32806),
            .I(n25));
    InMux I__5576 (
            .O(N__32803),
            .I(bfn_7_26_0_));
    CascadeMux I__5575 (
            .O(N__32800),
            .I(N__32796));
    InMux I__5574 (
            .O(N__32799),
            .I(N__32792));
    InMux I__5573 (
            .O(N__32796),
            .I(N__32789));
    InMux I__5572 (
            .O(N__32795),
            .I(N__32786));
    LocalMux I__5571 (
            .O(N__32792),
            .I(N__32783));
    LocalMux I__5570 (
            .O(N__32789),
            .I(encoder0_position_8));
    LocalMux I__5569 (
            .O(N__32786),
            .I(encoder0_position_8));
    Odrv12 I__5568 (
            .O(N__32783),
            .I(encoder0_position_8));
    InMux I__5567 (
            .O(N__32776),
            .I(N__32772));
    InMux I__5566 (
            .O(N__32775),
            .I(N__32768));
    LocalMux I__5565 (
            .O(N__32772),
            .I(N__32765));
    InMux I__5564 (
            .O(N__32771),
            .I(N__32762));
    LocalMux I__5563 (
            .O(N__32768),
            .I(N__32759));
    Sp12to4 I__5562 (
            .O(N__32765),
            .I(N__32756));
    LocalMux I__5561 (
            .O(N__32762),
            .I(N__32753));
    Span4Mux_v I__5560 (
            .O(N__32759),
            .I(N__32750));
    Span12Mux_v I__5559 (
            .O(N__32756),
            .I(N__32747));
    Span4Mux_h I__5558 (
            .O(N__32753),
            .I(N__32744));
    Odrv4 I__5557 (
            .O(N__32750),
            .I(n311));
    Odrv12 I__5556 (
            .O(N__32747),
            .I(n311));
    Odrv4 I__5555 (
            .O(N__32744),
            .I(n311));
    CascadeMux I__5554 (
            .O(N__32737),
            .I(N__32734));
    InMux I__5553 (
            .O(N__32734),
            .I(N__32729));
    InMux I__5552 (
            .O(N__32733),
            .I(N__32726));
    InMux I__5551 (
            .O(N__32732),
            .I(N__32723));
    LocalMux I__5550 (
            .O(N__32729),
            .I(encoder0_position_5));
    LocalMux I__5549 (
            .O(N__32726),
            .I(encoder0_position_5));
    LocalMux I__5548 (
            .O(N__32723),
            .I(encoder0_position_5));
    InMux I__5547 (
            .O(N__32716),
            .I(N__32711));
    InMux I__5546 (
            .O(N__32715),
            .I(N__32708));
    InMux I__5545 (
            .O(N__32714),
            .I(N__32705));
    LocalMux I__5544 (
            .O(N__32711),
            .I(N__32702));
    LocalMux I__5543 (
            .O(N__32708),
            .I(encoder0_position_15));
    LocalMux I__5542 (
            .O(N__32705),
            .I(encoder0_position_15));
    Odrv4 I__5541 (
            .O(N__32702),
            .I(encoder0_position_15));
    InMux I__5540 (
            .O(N__32695),
            .I(N__32691));
    InMux I__5539 (
            .O(N__32694),
            .I(N__32687));
    LocalMux I__5538 (
            .O(N__32691),
            .I(N__32684));
    InMux I__5537 (
            .O(N__32690),
            .I(N__32681));
    LocalMux I__5536 (
            .O(N__32687),
            .I(N__32678));
    Span4Mux_h I__5535 (
            .O(N__32684),
            .I(N__32675));
    LocalMux I__5534 (
            .O(N__32681),
            .I(N__32672));
    Span12Mux_s6_h I__5533 (
            .O(N__32678),
            .I(N__32669));
    Odrv4 I__5532 (
            .O(N__32675),
            .I(n304));
    Odrv12 I__5531 (
            .O(N__32672),
            .I(n304));
    Odrv12 I__5530 (
            .O(N__32669),
            .I(n304));
    InMux I__5529 (
            .O(N__32662),
            .I(N__32659));
    LocalMux I__5528 (
            .O(N__32659),
            .I(N__32656));
    Span4Mux_v I__5527 (
            .O(N__32656),
            .I(N__32652));
    InMux I__5526 (
            .O(N__32655),
            .I(N__32649));
    Span4Mux_h I__5525 (
            .O(N__32652),
            .I(N__32646));
    LocalMux I__5524 (
            .O(N__32649),
            .I(n2320));
    Odrv4 I__5523 (
            .O(N__32646),
            .I(n2320));
    InMux I__5522 (
            .O(N__32641),
            .I(N__32637));
    CascadeMux I__5521 (
            .O(N__32640),
            .I(N__32634));
    LocalMux I__5520 (
            .O(N__32637),
            .I(N__32631));
    InMux I__5519 (
            .O(N__32634),
            .I(N__32628));
    Span12Mux_v I__5518 (
            .O(N__32631),
            .I(N__32625));
    LocalMux I__5517 (
            .O(N__32628),
            .I(n2319));
    Odrv12 I__5516 (
            .O(N__32625),
            .I(n2319));
    CascadeMux I__5515 (
            .O(N__32620),
            .I(N__32617));
    InMux I__5514 (
            .O(N__32617),
            .I(N__32614));
    LocalMux I__5513 (
            .O(N__32614),
            .I(n14008));
    InMux I__5512 (
            .O(N__32611),
            .I(N__32608));
    LocalMux I__5511 (
            .O(N__32608),
            .I(n14006));
    InMux I__5510 (
            .O(N__32605),
            .I(N__32602));
    LocalMux I__5509 (
            .O(N__32602),
            .I(N__32599));
    Span4Mux_h I__5508 (
            .O(N__32599),
            .I(N__32596));
    Span4Mux_v I__5507 (
            .O(N__32596),
            .I(N__32593));
    Odrv4 I__5506 (
            .O(N__32593),
            .I(n14014));
    CascadeMux I__5505 (
            .O(N__32590),
            .I(N__32587));
    InMux I__5504 (
            .O(N__32587),
            .I(N__32582));
    InMux I__5503 (
            .O(N__32586),
            .I(N__32577));
    InMux I__5502 (
            .O(N__32585),
            .I(N__32577));
    LocalMux I__5501 (
            .O(N__32582),
            .I(encoder0_position_1));
    LocalMux I__5500 (
            .O(N__32577),
            .I(encoder0_position_1));
    InMux I__5499 (
            .O(N__32572),
            .I(N__32569));
    LocalMux I__5498 (
            .O(N__32569),
            .I(N__32565));
    InMux I__5497 (
            .O(N__32568),
            .I(N__32561));
    Span4Mux_v I__5496 (
            .O(N__32565),
            .I(N__32558));
    InMux I__5495 (
            .O(N__32564),
            .I(N__32555));
    LocalMux I__5494 (
            .O(N__32561),
            .I(encoder0_position_0));
    Odrv4 I__5493 (
            .O(N__32558),
            .I(encoder0_position_0));
    LocalMux I__5492 (
            .O(N__32555),
            .I(encoder0_position_0));
    CascadeMux I__5491 (
            .O(N__32548),
            .I(N__32545));
    InMux I__5490 (
            .O(N__32545),
            .I(N__32542));
    LocalMux I__5489 (
            .O(N__32542),
            .I(n33_adj_657));
    CascadeMux I__5488 (
            .O(N__32539),
            .I(N__32536));
    InMux I__5487 (
            .O(N__32536),
            .I(N__32533));
    LocalMux I__5486 (
            .O(N__32533),
            .I(N__32530));
    Span4Mux_v I__5485 (
            .O(N__32530),
            .I(N__32527));
    Odrv4 I__5484 (
            .O(N__32527),
            .I(n33));
    InMux I__5483 (
            .O(N__32524),
            .I(bfn_7_25_0_));
    InMux I__5482 (
            .O(N__32521),
            .I(N__32518));
    LocalMux I__5481 (
            .O(N__32518),
            .I(N__32515));
    Odrv4 I__5480 (
            .O(N__32515),
            .I(n2295));
    CascadeMux I__5479 (
            .O(N__32512),
            .I(N__32508));
    CascadeMux I__5478 (
            .O(N__32511),
            .I(N__32505));
    InMux I__5477 (
            .O(N__32508),
            .I(N__32502));
    InMux I__5476 (
            .O(N__32505),
            .I(N__32499));
    LocalMux I__5475 (
            .O(N__32502),
            .I(N__32495));
    LocalMux I__5474 (
            .O(N__32499),
            .I(N__32492));
    InMux I__5473 (
            .O(N__32498),
            .I(N__32489));
    Span4Mux_v I__5472 (
            .O(N__32495),
            .I(N__32482));
    Span4Mux_h I__5471 (
            .O(N__32492),
            .I(N__32482));
    LocalMux I__5470 (
            .O(N__32489),
            .I(N__32482));
    Odrv4 I__5469 (
            .O(N__32482),
            .I(n2228));
    InMux I__5468 (
            .O(N__32479),
            .I(N__32476));
    LocalMux I__5467 (
            .O(N__32476),
            .I(N__32472));
    InMux I__5466 (
            .O(N__32475),
            .I(N__32468));
    Span4Mux_v I__5465 (
            .O(N__32472),
            .I(N__32465));
    InMux I__5464 (
            .O(N__32471),
            .I(N__32462));
    LocalMux I__5463 (
            .O(N__32468),
            .I(encoder0_position_2));
    Odrv4 I__5462 (
            .O(N__32465),
            .I(encoder0_position_2));
    LocalMux I__5461 (
            .O(N__32462),
            .I(encoder0_position_2));
    CascadeMux I__5460 (
            .O(N__32455),
            .I(N__32452));
    InMux I__5459 (
            .O(N__32452),
            .I(N__32448));
    InMux I__5458 (
            .O(N__32451),
            .I(N__32444));
    LocalMux I__5457 (
            .O(N__32448),
            .I(N__32441));
    InMux I__5456 (
            .O(N__32447),
            .I(N__32438));
    LocalMux I__5455 (
            .O(N__32444),
            .I(N__32433));
    Span4Mux_h I__5454 (
            .O(N__32441),
            .I(N__32433));
    LocalMux I__5453 (
            .O(N__32438),
            .I(N__32430));
    Odrv4 I__5452 (
            .O(N__32433),
            .I(n2321));
    Odrv4 I__5451 (
            .O(N__32430),
            .I(n2321));
    CascadeMux I__5450 (
            .O(N__32425),
            .I(N__32422));
    InMux I__5449 (
            .O(N__32422),
            .I(N__32418));
    InMux I__5448 (
            .O(N__32421),
            .I(N__32415));
    LocalMux I__5447 (
            .O(N__32418),
            .I(N__32412));
    LocalMux I__5446 (
            .O(N__32415),
            .I(N__32408));
    Span4Mux_h I__5445 (
            .O(N__32412),
            .I(N__32405));
    InMux I__5444 (
            .O(N__32411),
            .I(N__32402));
    Odrv12 I__5443 (
            .O(N__32408),
            .I(n2324));
    Odrv4 I__5442 (
            .O(N__32405),
            .I(n2324));
    LocalMux I__5441 (
            .O(N__32402),
            .I(n2324));
    CascadeMux I__5440 (
            .O(N__32395),
            .I(N__32391));
    CascadeMux I__5439 (
            .O(N__32394),
            .I(N__32388));
    InMux I__5438 (
            .O(N__32391),
            .I(N__32385));
    InMux I__5437 (
            .O(N__32388),
            .I(N__32381));
    LocalMux I__5436 (
            .O(N__32385),
            .I(N__32378));
    InMux I__5435 (
            .O(N__32384),
            .I(N__32375));
    LocalMux I__5434 (
            .O(N__32381),
            .I(N__32372));
    Span4Mux_h I__5433 (
            .O(N__32378),
            .I(N__32369));
    LocalMux I__5432 (
            .O(N__32375),
            .I(n2328));
    Odrv4 I__5431 (
            .O(N__32372),
            .I(n2328));
    Odrv4 I__5430 (
            .O(N__32369),
            .I(n2328));
    CascadeMux I__5429 (
            .O(N__32362),
            .I(N__32359));
    InMux I__5428 (
            .O(N__32359),
            .I(N__32355));
    InMux I__5427 (
            .O(N__32358),
            .I(N__32352));
    LocalMux I__5426 (
            .O(N__32355),
            .I(N__32349));
    LocalMux I__5425 (
            .O(N__32352),
            .I(N__32343));
    Span12Mux_s6_h I__5424 (
            .O(N__32349),
            .I(N__32343));
    InMux I__5423 (
            .O(N__32348),
            .I(N__32340));
    Odrv12 I__5422 (
            .O(N__32343),
            .I(n2327));
    LocalMux I__5421 (
            .O(N__32340),
            .I(n2327));
    CascadeMux I__5420 (
            .O(N__32335),
            .I(N__32331));
    InMux I__5419 (
            .O(N__32334),
            .I(N__32328));
    InMux I__5418 (
            .O(N__32331),
            .I(N__32325));
    LocalMux I__5417 (
            .O(N__32328),
            .I(N__32322));
    LocalMux I__5416 (
            .O(N__32325),
            .I(N__32319));
    Span4Mux_h I__5415 (
            .O(N__32322),
            .I(N__32315));
    Span4Mux_h I__5414 (
            .O(N__32319),
            .I(N__32312));
    InMux I__5413 (
            .O(N__32318),
            .I(N__32309));
    Odrv4 I__5412 (
            .O(N__32315),
            .I(n2322));
    Odrv4 I__5411 (
            .O(N__32312),
            .I(n2322));
    LocalMux I__5410 (
            .O(N__32309),
            .I(n2322));
    CascadeMux I__5409 (
            .O(N__32302),
            .I(N__32299));
    InMux I__5408 (
            .O(N__32299),
            .I(N__32295));
    InMux I__5407 (
            .O(N__32298),
            .I(N__32292));
    LocalMux I__5406 (
            .O(N__32295),
            .I(N__32289));
    LocalMux I__5405 (
            .O(N__32292),
            .I(N__32286));
    Span4Mux_v I__5404 (
            .O(N__32289),
            .I(N__32281));
    Span4Mux_v I__5403 (
            .O(N__32286),
            .I(N__32281));
    Odrv4 I__5402 (
            .O(N__32281),
            .I(n2326));
    CascadeMux I__5401 (
            .O(N__32278),
            .I(N__32273));
    CascadeMux I__5400 (
            .O(N__32277),
            .I(N__32270));
    InMux I__5399 (
            .O(N__32276),
            .I(N__32267));
    InMux I__5398 (
            .O(N__32273),
            .I(N__32264));
    InMux I__5397 (
            .O(N__32270),
            .I(N__32261));
    LocalMux I__5396 (
            .O(N__32267),
            .I(N__32256));
    LocalMux I__5395 (
            .O(N__32264),
            .I(N__32256));
    LocalMux I__5394 (
            .O(N__32261),
            .I(N__32253));
    Span4Mux_v I__5393 (
            .O(N__32256),
            .I(N__32248));
    Span4Mux_v I__5392 (
            .O(N__32253),
            .I(N__32248));
    Odrv4 I__5391 (
            .O(N__32248),
            .I(n2325));
    CascadeMux I__5390 (
            .O(N__32245),
            .I(N__32242));
    InMux I__5389 (
            .O(N__32242),
            .I(N__32238));
    InMux I__5388 (
            .O(N__32241),
            .I(N__32235));
    LocalMux I__5387 (
            .O(N__32238),
            .I(N__32232));
    LocalMux I__5386 (
            .O(N__32235),
            .I(N__32229));
    Span4Mux_s3_h I__5385 (
            .O(N__32232),
            .I(N__32226));
    Span4Mux_h I__5384 (
            .O(N__32229),
            .I(N__32222));
    Span4Mux_v I__5383 (
            .O(N__32226),
            .I(N__32219));
    InMux I__5382 (
            .O(N__32225),
            .I(N__32216));
    Odrv4 I__5381 (
            .O(N__32222),
            .I(n2323));
    Odrv4 I__5380 (
            .O(N__32219),
            .I(n2323));
    LocalMux I__5379 (
            .O(N__32216),
            .I(n2323));
    InMux I__5378 (
            .O(N__32209),
            .I(N__32205));
    CascadeMux I__5377 (
            .O(N__32208),
            .I(N__32202));
    LocalMux I__5376 (
            .O(N__32205),
            .I(N__32198));
    InMux I__5375 (
            .O(N__32202),
            .I(N__32195));
    InMux I__5374 (
            .O(N__32201),
            .I(N__32192));
    Span4Mux_v I__5373 (
            .O(N__32198),
            .I(N__32189));
    LocalMux I__5372 (
            .O(N__32195),
            .I(encoder0_position_3));
    LocalMux I__5371 (
            .O(N__32192),
            .I(encoder0_position_3));
    Odrv4 I__5370 (
            .O(N__32189),
            .I(encoder0_position_3));
    InMux I__5369 (
            .O(N__32182),
            .I(N__32177));
    InMux I__5368 (
            .O(N__32181),
            .I(N__32174));
    InMux I__5367 (
            .O(N__32180),
            .I(N__32171));
    LocalMux I__5366 (
            .O(N__32177),
            .I(N__32168));
    LocalMux I__5365 (
            .O(N__32174),
            .I(encoder0_position_11));
    LocalMux I__5364 (
            .O(N__32171),
            .I(encoder0_position_11));
    Odrv4 I__5363 (
            .O(N__32168),
            .I(encoder0_position_11));
    InMux I__5362 (
            .O(N__32161),
            .I(N__32157));
    InMux I__5361 (
            .O(N__32160),
            .I(N__32154));
    LocalMux I__5360 (
            .O(N__32157),
            .I(N__32149));
    LocalMux I__5359 (
            .O(N__32154),
            .I(N__32149));
    Span4Mux_h I__5358 (
            .O(N__32149),
            .I(N__32145));
    InMux I__5357 (
            .O(N__32148),
            .I(N__32142));
    Span4Mux_s3_h I__5356 (
            .O(N__32145),
            .I(N__32137));
    LocalMux I__5355 (
            .O(N__32142),
            .I(N__32137));
    Span4Mux_h I__5354 (
            .O(N__32137),
            .I(N__32134));
    Odrv4 I__5353 (
            .O(N__32134),
            .I(n308));
    InMux I__5352 (
            .O(N__32131),
            .I(n12289));
    InMux I__5351 (
            .O(N__32128),
            .I(N__32125));
    LocalMux I__5350 (
            .O(N__32125),
            .I(N__32122));
    Span4Mux_v I__5349 (
            .O(N__32122),
            .I(N__32118));
    InMux I__5348 (
            .O(N__32121),
            .I(N__32115));
    Odrv4 I__5347 (
            .O(N__32118),
            .I(n2219));
    LocalMux I__5346 (
            .O(N__32115),
            .I(n2219));
    InMux I__5345 (
            .O(N__32110),
            .I(N__32107));
    LocalMux I__5344 (
            .O(N__32107),
            .I(N__32104));
    Span4Mux_h I__5343 (
            .O(N__32104),
            .I(N__32101));
    Odrv4 I__5342 (
            .O(N__32101),
            .I(n2286_adj_600));
    InMux I__5341 (
            .O(N__32098),
            .I(n12290));
    InMux I__5340 (
            .O(N__32095),
            .I(N__32092));
    LocalMux I__5339 (
            .O(N__32092),
            .I(N__32089));
    Span4Mux_h I__5338 (
            .O(N__32089),
            .I(N__32084));
    InMux I__5337 (
            .O(N__32088),
            .I(N__32079));
    InMux I__5336 (
            .O(N__32087),
            .I(N__32079));
    Odrv4 I__5335 (
            .O(N__32084),
            .I(n2218));
    LocalMux I__5334 (
            .O(N__32079),
            .I(n2218));
    CascadeMux I__5333 (
            .O(N__32074),
            .I(N__32071));
    InMux I__5332 (
            .O(N__32071),
            .I(N__32068));
    LocalMux I__5331 (
            .O(N__32068),
            .I(N__32065));
    Span4Mux_v I__5330 (
            .O(N__32065),
            .I(N__32062));
    Span4Mux_h I__5329 (
            .O(N__32062),
            .I(N__32059));
    Odrv4 I__5328 (
            .O(N__32059),
            .I(n2285_adj_599));
    InMux I__5327 (
            .O(N__32056),
            .I(bfn_7_22_0_));
    InMux I__5326 (
            .O(N__32053),
            .I(n12292));
    InMux I__5325 (
            .O(N__32050),
            .I(N__32047));
    LocalMux I__5324 (
            .O(N__32047),
            .I(N__32043));
    InMux I__5323 (
            .O(N__32046),
            .I(N__32040));
    Span4Mux_v I__5322 (
            .O(N__32043),
            .I(N__32036));
    LocalMux I__5321 (
            .O(N__32040),
            .I(N__32033));
    InMux I__5320 (
            .O(N__32039),
            .I(N__32030));
    Span4Mux_h I__5319 (
            .O(N__32036),
            .I(N__32027));
    Span4Mux_v I__5318 (
            .O(N__32033),
            .I(N__32022));
    LocalMux I__5317 (
            .O(N__32030),
            .I(N__32022));
    Odrv4 I__5316 (
            .O(N__32027),
            .I(n2216));
    Odrv4 I__5315 (
            .O(N__32022),
            .I(n2216));
    InMux I__5314 (
            .O(N__32017),
            .I(N__32014));
    LocalMux I__5313 (
            .O(N__32014),
            .I(n2283));
    InMux I__5312 (
            .O(N__32011),
            .I(n12293));
    CascadeMux I__5311 (
            .O(N__32008),
            .I(N__32004));
    InMux I__5310 (
            .O(N__32007),
            .I(N__32001));
    InMux I__5309 (
            .O(N__32004),
            .I(N__31998));
    LocalMux I__5308 (
            .O(N__32001),
            .I(N__31995));
    LocalMux I__5307 (
            .O(N__31998),
            .I(N__31992));
    Span4Mux_h I__5306 (
            .O(N__31995),
            .I(N__31988));
    Span4Mux_v I__5305 (
            .O(N__31992),
            .I(N__31985));
    InMux I__5304 (
            .O(N__31991),
            .I(N__31982));
    Span4Mux_h I__5303 (
            .O(N__31988),
            .I(N__31979));
    Span4Mux_h I__5302 (
            .O(N__31985),
            .I(N__31974));
    LocalMux I__5301 (
            .O(N__31982),
            .I(N__31974));
    Odrv4 I__5300 (
            .O(N__31979),
            .I(n2215));
    Odrv4 I__5299 (
            .O(N__31974),
            .I(n2215));
    InMux I__5298 (
            .O(N__31969),
            .I(N__31966));
    LocalMux I__5297 (
            .O(N__31966),
            .I(N__31963));
    Span4Mux_v I__5296 (
            .O(N__31963),
            .I(N__31960));
    Odrv4 I__5295 (
            .O(N__31960),
            .I(n2282));
    InMux I__5294 (
            .O(N__31957),
            .I(n12294));
    InMux I__5293 (
            .O(N__31954),
            .I(N__31950));
    CascadeMux I__5292 (
            .O(N__31953),
            .I(N__31947));
    LocalMux I__5291 (
            .O(N__31950),
            .I(N__31944));
    InMux I__5290 (
            .O(N__31947),
            .I(N__31941));
    Span4Mux_h I__5289 (
            .O(N__31944),
            .I(N__31938));
    LocalMux I__5288 (
            .O(N__31941),
            .I(N__31935));
    Span4Mux_h I__5287 (
            .O(N__31938),
            .I(N__31932));
    Span4Mux_v I__5286 (
            .O(N__31935),
            .I(N__31929));
    Odrv4 I__5285 (
            .O(N__31932),
            .I(n2214));
    Odrv4 I__5284 (
            .O(N__31929),
            .I(n2214));
    InMux I__5283 (
            .O(N__31924),
            .I(n12295));
    CascadeMux I__5282 (
            .O(N__31921),
            .I(N__31918));
    InMux I__5281 (
            .O(N__31918),
            .I(N__31914));
    InMux I__5280 (
            .O(N__31917),
            .I(N__31911));
    LocalMux I__5279 (
            .O(N__31914),
            .I(N__31906));
    LocalMux I__5278 (
            .O(N__31911),
            .I(N__31906));
    Span4Mux_v I__5277 (
            .O(N__31906),
            .I(N__31903));
    Odrv4 I__5276 (
            .O(N__31903),
            .I(n2313));
    InMux I__5275 (
            .O(N__31900),
            .I(N__31896));
    CascadeMux I__5274 (
            .O(N__31899),
            .I(N__31893));
    LocalMux I__5273 (
            .O(N__31896),
            .I(N__31889));
    InMux I__5272 (
            .O(N__31893),
            .I(N__31886));
    InMux I__5271 (
            .O(N__31892),
            .I(N__31883));
    Odrv4 I__5270 (
            .O(N__31889),
            .I(n2225));
    LocalMux I__5269 (
            .O(N__31886),
            .I(n2225));
    LocalMux I__5268 (
            .O(N__31883),
            .I(n2225));
    CascadeMux I__5267 (
            .O(N__31876),
            .I(N__31873));
    InMux I__5266 (
            .O(N__31873),
            .I(N__31870));
    LocalMux I__5265 (
            .O(N__31870),
            .I(n2292));
    InMux I__5264 (
            .O(N__31867),
            .I(N__31863));
    CascadeMux I__5263 (
            .O(N__31866),
            .I(N__31860));
    LocalMux I__5262 (
            .O(N__31863),
            .I(N__31857));
    InMux I__5261 (
            .O(N__31860),
            .I(N__31854));
    Odrv4 I__5260 (
            .O(N__31857),
            .I(n2224));
    LocalMux I__5259 (
            .O(N__31854),
            .I(n2224));
    InMux I__5258 (
            .O(N__31849),
            .I(N__31846));
    LocalMux I__5257 (
            .O(N__31846),
            .I(n2291));
    InMux I__5256 (
            .O(N__31843),
            .I(n12281));
    CascadeMux I__5255 (
            .O(N__31840),
            .I(N__31836));
    InMux I__5254 (
            .O(N__31839),
            .I(N__31832));
    InMux I__5253 (
            .O(N__31836),
            .I(N__31829));
    InMux I__5252 (
            .O(N__31835),
            .I(N__31826));
    LocalMux I__5251 (
            .O(N__31832),
            .I(N__31819));
    LocalMux I__5250 (
            .O(N__31829),
            .I(N__31819));
    LocalMux I__5249 (
            .O(N__31826),
            .I(N__31819));
    Odrv12 I__5248 (
            .O(N__31819),
            .I(n2227));
    CascadeMux I__5247 (
            .O(N__31816),
            .I(N__31813));
    InMux I__5246 (
            .O(N__31813),
            .I(N__31810));
    LocalMux I__5245 (
            .O(N__31810),
            .I(N__31807));
    Odrv4 I__5244 (
            .O(N__31807),
            .I(n2294));
    InMux I__5243 (
            .O(N__31804),
            .I(n12282));
    CascadeMux I__5242 (
            .O(N__31801),
            .I(N__31797));
    CascadeMux I__5241 (
            .O(N__31800),
            .I(N__31794));
    InMux I__5240 (
            .O(N__31797),
            .I(N__31790));
    InMux I__5239 (
            .O(N__31794),
            .I(N__31787));
    InMux I__5238 (
            .O(N__31793),
            .I(N__31784));
    LocalMux I__5237 (
            .O(N__31790),
            .I(n2226));
    LocalMux I__5236 (
            .O(N__31787),
            .I(n2226));
    LocalMux I__5235 (
            .O(N__31784),
            .I(n2226));
    InMux I__5234 (
            .O(N__31777),
            .I(N__31774));
    LocalMux I__5233 (
            .O(N__31774),
            .I(n2293));
    InMux I__5232 (
            .O(N__31771),
            .I(bfn_7_21_0_));
    InMux I__5231 (
            .O(N__31768),
            .I(n12284));
    InMux I__5230 (
            .O(N__31765),
            .I(n12285));
    CascadeMux I__5229 (
            .O(N__31762),
            .I(N__31758));
    InMux I__5228 (
            .O(N__31761),
            .I(N__31755));
    InMux I__5227 (
            .O(N__31758),
            .I(N__31752));
    LocalMux I__5226 (
            .O(N__31755),
            .I(N__31749));
    LocalMux I__5225 (
            .O(N__31752),
            .I(n2223));
    Odrv4 I__5224 (
            .O(N__31749),
            .I(n2223));
    InMux I__5223 (
            .O(N__31744),
            .I(N__31741));
    LocalMux I__5222 (
            .O(N__31741),
            .I(n2290_adj_604));
    InMux I__5221 (
            .O(N__31738),
            .I(n12286));
    InMux I__5220 (
            .O(N__31735),
            .I(N__31731));
    InMux I__5219 (
            .O(N__31734),
            .I(N__31727));
    LocalMux I__5218 (
            .O(N__31731),
            .I(N__31724));
    InMux I__5217 (
            .O(N__31730),
            .I(N__31721));
    LocalMux I__5216 (
            .O(N__31727),
            .I(n2222));
    Odrv12 I__5215 (
            .O(N__31724),
            .I(n2222));
    LocalMux I__5214 (
            .O(N__31721),
            .I(n2222));
    CascadeMux I__5213 (
            .O(N__31714),
            .I(N__31711));
    InMux I__5212 (
            .O(N__31711),
            .I(N__31708));
    LocalMux I__5211 (
            .O(N__31708),
            .I(n2289_adj_603));
    InMux I__5210 (
            .O(N__31705),
            .I(n12287));
    InMux I__5209 (
            .O(N__31702),
            .I(N__31698));
    InMux I__5208 (
            .O(N__31701),
            .I(N__31695));
    LocalMux I__5207 (
            .O(N__31698),
            .I(N__31692));
    LocalMux I__5206 (
            .O(N__31695),
            .I(N__31689));
    Span4Mux_v I__5205 (
            .O(N__31692),
            .I(N__31686));
    Span4Mux_h I__5204 (
            .O(N__31689),
            .I(N__31683));
    Odrv4 I__5203 (
            .O(N__31686),
            .I(n2221));
    Odrv4 I__5202 (
            .O(N__31683),
            .I(n2221));
    InMux I__5201 (
            .O(N__31678),
            .I(N__31675));
    LocalMux I__5200 (
            .O(N__31675),
            .I(N__31672));
    Span4Mux_h I__5199 (
            .O(N__31672),
            .I(N__31669));
    Odrv4 I__5198 (
            .O(N__31669),
            .I(n2288_adj_602));
    InMux I__5197 (
            .O(N__31666),
            .I(n12288));
    InMux I__5196 (
            .O(N__31663),
            .I(N__31660));
    LocalMux I__5195 (
            .O(N__31660),
            .I(N__31656));
    InMux I__5194 (
            .O(N__31659),
            .I(N__31653));
    Span4Mux_v I__5193 (
            .O(N__31656),
            .I(N__31648));
    LocalMux I__5192 (
            .O(N__31653),
            .I(N__31648));
    Span4Mux_h I__5191 (
            .O(N__31648),
            .I(N__31645));
    Odrv4 I__5190 (
            .O(N__31645),
            .I(n2220));
    InMux I__5189 (
            .O(N__31642),
            .I(N__31639));
    LocalMux I__5188 (
            .O(N__31639),
            .I(N__31636));
    Span4Mux_s2_h I__5187 (
            .O(N__31636),
            .I(N__31633));
    Span4Mux_h I__5186 (
            .O(N__31633),
            .I(N__31630));
    Odrv4 I__5185 (
            .O(N__31630),
            .I(n2287_adj_601));
    CascadeMux I__5184 (
            .O(N__31627),
            .I(N__31624));
    InMux I__5183 (
            .O(N__31624),
            .I(N__31620));
    InMux I__5182 (
            .O(N__31623),
            .I(N__31616));
    LocalMux I__5181 (
            .O(N__31620),
            .I(N__31613));
    InMux I__5180 (
            .O(N__31619),
            .I(N__31610));
    LocalMux I__5179 (
            .O(N__31616),
            .I(n2532));
    Odrv12 I__5178 (
            .O(N__31613),
            .I(n2532));
    LocalMux I__5177 (
            .O(N__31610),
            .I(n2532));
    CascadeMux I__5176 (
            .O(N__31603),
            .I(N__31600));
    InMux I__5175 (
            .O(N__31600),
            .I(N__31597));
    LocalMux I__5174 (
            .O(N__31597),
            .I(N__31594));
    Span4Mux_v I__5173 (
            .O(N__31594),
            .I(N__31591));
    Odrv4 I__5172 (
            .O(N__31591),
            .I(n2599));
    InMux I__5171 (
            .O(N__31588),
            .I(N__31585));
    LocalMux I__5170 (
            .O(N__31585),
            .I(n2483));
    InMux I__5169 (
            .O(N__31582),
            .I(N__31579));
    LocalMux I__5168 (
            .O(N__31579),
            .I(N__31575));
    InMux I__5167 (
            .O(N__31578),
            .I(N__31572));
    Span4Mux_h I__5166 (
            .O(N__31575),
            .I(N__31568));
    LocalMux I__5165 (
            .O(N__31572),
            .I(N__31565));
    InMux I__5164 (
            .O(N__31571),
            .I(N__31562));
    Odrv4 I__5163 (
            .O(N__31568),
            .I(n2416));
    Odrv4 I__5162 (
            .O(N__31565),
            .I(n2416));
    LocalMux I__5161 (
            .O(N__31562),
            .I(n2416));
    InMux I__5160 (
            .O(N__31555),
            .I(N__31552));
    LocalMux I__5159 (
            .O(N__31552),
            .I(N__31549));
    Span4Mux_h I__5158 (
            .O(N__31549),
            .I(N__31544));
    InMux I__5157 (
            .O(N__31548),
            .I(N__31539));
    InMux I__5156 (
            .O(N__31547),
            .I(N__31539));
    Odrv4 I__5155 (
            .O(N__31544),
            .I(n2515));
    LocalMux I__5154 (
            .O(N__31539),
            .I(n2515));
    InMux I__5153 (
            .O(N__31534),
            .I(N__31531));
    LocalMux I__5152 (
            .O(N__31531),
            .I(N__31528));
    Odrv12 I__5151 (
            .O(N__31528),
            .I(n2301));
    InMux I__5150 (
            .O(N__31525),
            .I(bfn_7_20_0_));
    CascadeMux I__5149 (
            .O(N__31522),
            .I(N__31518));
    InMux I__5148 (
            .O(N__31521),
            .I(N__31514));
    InMux I__5147 (
            .O(N__31518),
            .I(N__31511));
    InMux I__5146 (
            .O(N__31517),
            .I(N__31508));
    LocalMux I__5145 (
            .O(N__31514),
            .I(N__31503));
    LocalMux I__5144 (
            .O(N__31511),
            .I(N__31503));
    LocalMux I__5143 (
            .O(N__31508),
            .I(n2233));
    Odrv12 I__5142 (
            .O(N__31503),
            .I(n2233));
    CascadeMux I__5141 (
            .O(N__31498),
            .I(N__31495));
    InMux I__5140 (
            .O(N__31495),
            .I(N__31492));
    LocalMux I__5139 (
            .O(N__31492),
            .I(N__31489));
    Span4Mux_h I__5138 (
            .O(N__31489),
            .I(N__31486));
    Odrv4 I__5137 (
            .O(N__31486),
            .I(n2300));
    InMux I__5136 (
            .O(N__31483),
            .I(n12276));
    CascadeMux I__5135 (
            .O(N__31480),
            .I(N__31477));
    InMux I__5134 (
            .O(N__31477),
            .I(N__31473));
    InMux I__5133 (
            .O(N__31476),
            .I(N__31470));
    LocalMux I__5132 (
            .O(N__31473),
            .I(N__31467));
    LocalMux I__5131 (
            .O(N__31470),
            .I(N__31462));
    Span4Mux_h I__5130 (
            .O(N__31467),
            .I(N__31462));
    Span4Mux_h I__5129 (
            .O(N__31462),
            .I(N__31459));
    Odrv4 I__5128 (
            .O(N__31459),
            .I(n2232));
    InMux I__5127 (
            .O(N__31456),
            .I(N__31453));
    LocalMux I__5126 (
            .O(N__31453),
            .I(N__31450));
    Span12Mux_s6_h I__5125 (
            .O(N__31450),
            .I(N__31447));
    Odrv12 I__5124 (
            .O(N__31447),
            .I(n2299));
    InMux I__5123 (
            .O(N__31444),
            .I(n12277));
    CascadeMux I__5122 (
            .O(N__31441),
            .I(N__31438));
    InMux I__5121 (
            .O(N__31438),
            .I(N__31434));
    CascadeMux I__5120 (
            .O(N__31437),
            .I(N__31430));
    LocalMux I__5119 (
            .O(N__31434),
            .I(N__31427));
    InMux I__5118 (
            .O(N__31433),
            .I(N__31422));
    InMux I__5117 (
            .O(N__31430),
            .I(N__31422));
    Span4Mux_h I__5116 (
            .O(N__31427),
            .I(N__31419));
    LocalMux I__5115 (
            .O(N__31422),
            .I(n2231));
    Odrv4 I__5114 (
            .O(N__31419),
            .I(n2231));
    InMux I__5113 (
            .O(N__31414),
            .I(N__31411));
    LocalMux I__5112 (
            .O(N__31411),
            .I(N__31408));
    Odrv4 I__5111 (
            .O(N__31408),
            .I(n2298));
    InMux I__5110 (
            .O(N__31405),
            .I(n12278));
    CascadeMux I__5109 (
            .O(N__31402),
            .I(N__31399));
    InMux I__5108 (
            .O(N__31399),
            .I(N__31396));
    LocalMux I__5107 (
            .O(N__31396),
            .I(N__31392));
    CascadeMux I__5106 (
            .O(N__31395),
            .I(N__31389));
    Span4Mux_v I__5105 (
            .O(N__31392),
            .I(N__31386));
    InMux I__5104 (
            .O(N__31389),
            .I(N__31383));
    Odrv4 I__5103 (
            .O(N__31386),
            .I(n2230));
    LocalMux I__5102 (
            .O(N__31383),
            .I(n2230));
    InMux I__5101 (
            .O(N__31378),
            .I(N__31375));
    LocalMux I__5100 (
            .O(N__31375),
            .I(N__31372));
    Span4Mux_v I__5099 (
            .O(N__31372),
            .I(N__31369));
    Odrv4 I__5098 (
            .O(N__31369),
            .I(n2297));
    InMux I__5097 (
            .O(N__31366),
            .I(n12279));
    CascadeMux I__5096 (
            .O(N__31363),
            .I(N__31359));
    CascadeMux I__5095 (
            .O(N__31362),
            .I(N__31355));
    InMux I__5094 (
            .O(N__31359),
            .I(N__31352));
    InMux I__5093 (
            .O(N__31358),
            .I(N__31349));
    InMux I__5092 (
            .O(N__31355),
            .I(N__31346));
    LocalMux I__5091 (
            .O(N__31352),
            .I(N__31343));
    LocalMux I__5090 (
            .O(N__31349),
            .I(N__31340));
    LocalMux I__5089 (
            .O(N__31346),
            .I(n2229));
    Odrv12 I__5088 (
            .O(N__31343),
            .I(n2229));
    Odrv4 I__5087 (
            .O(N__31340),
            .I(n2229));
    InMux I__5086 (
            .O(N__31333),
            .I(N__31330));
    LocalMux I__5085 (
            .O(N__31330),
            .I(N__31327));
    Odrv12 I__5084 (
            .O(N__31327),
            .I(n2296));
    InMux I__5083 (
            .O(N__31324),
            .I(n12280));
    InMux I__5082 (
            .O(N__31321),
            .I(N__31318));
    LocalMux I__5081 (
            .O(N__31318),
            .I(N__31315));
    Odrv4 I__5080 (
            .O(N__31315),
            .I(n2591));
    CascadeMux I__5079 (
            .O(N__31312),
            .I(n2524_cascade_));
    CascadeMux I__5078 (
            .O(N__31309),
            .I(N__31306));
    InMux I__5077 (
            .O(N__31306),
            .I(N__31303));
    LocalMux I__5076 (
            .O(N__31303),
            .I(N__31300));
    Odrv12 I__5075 (
            .O(N__31300),
            .I(n2391));
    CascadeMux I__5074 (
            .O(N__31297),
            .I(N__31293));
    CascadeMux I__5073 (
            .O(N__31296),
            .I(N__31289));
    InMux I__5072 (
            .O(N__31293),
            .I(N__31286));
    InMux I__5071 (
            .O(N__31292),
            .I(N__31283));
    InMux I__5070 (
            .O(N__31289),
            .I(N__31280));
    LocalMux I__5069 (
            .O(N__31286),
            .I(N__31275));
    LocalMux I__5068 (
            .O(N__31283),
            .I(N__31275));
    LocalMux I__5067 (
            .O(N__31280),
            .I(n2423));
    Odrv4 I__5066 (
            .O(N__31275),
            .I(n2423));
    InMux I__5065 (
            .O(N__31270),
            .I(N__31267));
    LocalMux I__5064 (
            .O(N__31267),
            .I(N__31264));
    Span4Mux_v I__5063 (
            .O(N__31264),
            .I(N__31261));
    Odrv4 I__5062 (
            .O(N__31261),
            .I(n2601));
    CascadeMux I__5061 (
            .O(N__31258),
            .I(N__31255));
    InMux I__5060 (
            .O(N__31255),
            .I(N__31252));
    LocalMux I__5059 (
            .O(N__31252),
            .I(N__31249));
    Span4Mux_h I__5058 (
            .O(N__31249),
            .I(N__31246));
    Span4Mux_h I__5057 (
            .O(N__31246),
            .I(N__31243));
    Odrv4 I__5056 (
            .O(N__31243),
            .I(n2394));
    CascadeMux I__5055 (
            .O(N__31240),
            .I(N__31236));
    CascadeMux I__5054 (
            .O(N__31239),
            .I(N__31233));
    InMux I__5053 (
            .O(N__31236),
            .I(N__31229));
    InMux I__5052 (
            .O(N__31233),
            .I(N__31226));
    CascadeMux I__5051 (
            .O(N__31232),
            .I(N__31223));
    LocalMux I__5050 (
            .O(N__31229),
            .I(N__31218));
    LocalMux I__5049 (
            .O(N__31226),
            .I(N__31218));
    InMux I__5048 (
            .O(N__31223),
            .I(N__31215));
    Span4Mux_v I__5047 (
            .O(N__31218),
            .I(N__31212));
    LocalMux I__5046 (
            .O(N__31215),
            .I(n2426));
    Odrv4 I__5045 (
            .O(N__31212),
            .I(n2426));
    InMux I__5044 (
            .O(N__31207),
            .I(N__31204));
    LocalMux I__5043 (
            .O(N__31204),
            .I(n2480));
    CascadeMux I__5042 (
            .O(N__31201),
            .I(N__31198));
    InMux I__5041 (
            .O(N__31198),
            .I(N__31195));
    LocalMux I__5040 (
            .O(N__31195),
            .I(N__31190));
    InMux I__5039 (
            .O(N__31194),
            .I(N__31187));
    InMux I__5038 (
            .O(N__31193),
            .I(N__31184));
    Odrv4 I__5037 (
            .O(N__31190),
            .I(n2413));
    LocalMux I__5036 (
            .O(N__31187),
            .I(n2413));
    LocalMux I__5035 (
            .O(N__31184),
            .I(n2413));
    CascadeMux I__5034 (
            .O(N__31177),
            .I(N__31174));
    InMux I__5033 (
            .O(N__31174),
            .I(N__31171));
    LocalMux I__5032 (
            .O(N__31171),
            .I(N__31166));
    InMux I__5031 (
            .O(N__31170),
            .I(N__31161));
    InMux I__5030 (
            .O(N__31169),
            .I(N__31161));
    Odrv4 I__5029 (
            .O(N__31166),
            .I(n2512));
    LocalMux I__5028 (
            .O(N__31161),
            .I(n2512));
    CascadeMux I__5027 (
            .O(N__31156),
            .I(N__31153));
    InMux I__5026 (
            .O(N__31153),
            .I(N__31150));
    LocalMux I__5025 (
            .O(N__31150),
            .I(N__31147));
    Span4Mux_v I__5024 (
            .O(N__31147),
            .I(N__31144));
    Span4Mux_h I__5023 (
            .O(N__31144),
            .I(N__31141));
    Odrv4 I__5022 (
            .O(N__31141),
            .I(n2388));
    InMux I__5021 (
            .O(N__31138),
            .I(N__31134));
    CascadeMux I__5020 (
            .O(N__31137),
            .I(N__31131));
    LocalMux I__5019 (
            .O(N__31134),
            .I(N__31128));
    InMux I__5018 (
            .O(N__31131),
            .I(N__31125));
    Span4Mux_h I__5017 (
            .O(N__31128),
            .I(N__31122));
    LocalMux I__5016 (
            .O(N__31125),
            .I(n2420));
    Odrv4 I__5015 (
            .O(N__31122),
            .I(n2420));
    InMux I__5014 (
            .O(N__31117),
            .I(N__31114));
    LocalMux I__5013 (
            .O(N__31114),
            .I(n2487));
    CascadeMux I__5012 (
            .O(N__31111),
            .I(n2420_cascade_));
    InMux I__5011 (
            .O(N__31108),
            .I(N__31104));
    InMux I__5010 (
            .O(N__31107),
            .I(N__31101));
    LocalMux I__5009 (
            .O(N__31104),
            .I(N__31098));
    LocalMux I__5008 (
            .O(N__31101),
            .I(N__31095));
    Span4Mux_h I__5007 (
            .O(N__31098),
            .I(N__31092));
    Span4Mux_h I__5006 (
            .O(N__31095),
            .I(N__31089));
    Odrv4 I__5005 (
            .O(N__31092),
            .I(n2519));
    Odrv4 I__5004 (
            .O(N__31089),
            .I(n2519));
    CascadeMux I__5003 (
            .O(N__31084),
            .I(n2519_cascade_));
    InMux I__5002 (
            .O(N__31081),
            .I(N__31078));
    LocalMux I__5001 (
            .O(N__31078),
            .I(N__31075));
    Span4Mux_v I__5000 (
            .O(N__31075),
            .I(N__31072));
    Odrv4 I__4999 (
            .O(N__31072),
            .I(n2586));
    CascadeMux I__4998 (
            .O(N__31069),
            .I(n2628_cascade_));
    InMux I__4997 (
            .O(N__31066),
            .I(N__31063));
    LocalMux I__4996 (
            .O(N__31063),
            .I(n2585));
    InMux I__4995 (
            .O(N__31060),
            .I(N__31057));
    LocalMux I__4994 (
            .O(N__31057),
            .I(N__31053));
    InMux I__4993 (
            .O(N__31056),
            .I(N__31050));
    Span4Mux_v I__4992 (
            .O(N__31053),
            .I(N__31046));
    LocalMux I__4991 (
            .O(N__31050),
            .I(N__31043));
    InMux I__4990 (
            .O(N__31049),
            .I(N__31040));
    Odrv4 I__4989 (
            .O(N__31046),
            .I(n2518));
    Odrv4 I__4988 (
            .O(N__31043),
            .I(n2518));
    LocalMux I__4987 (
            .O(N__31040),
            .I(n2518));
    InMux I__4986 (
            .O(N__31033),
            .I(N__31029));
    CascadeMux I__4985 (
            .O(N__31032),
            .I(N__31026));
    LocalMux I__4984 (
            .O(N__31029),
            .I(N__31023));
    InMux I__4983 (
            .O(N__31026),
            .I(N__31020));
    Span4Mux_v I__4982 (
            .O(N__31023),
            .I(N__31014));
    LocalMux I__4981 (
            .O(N__31020),
            .I(N__31014));
    InMux I__4980 (
            .O(N__31019),
            .I(N__31011));
    Odrv4 I__4979 (
            .O(N__31014),
            .I(n2417));
    LocalMux I__4978 (
            .O(N__31011),
            .I(n2417));
    InMux I__4977 (
            .O(N__31006),
            .I(N__31003));
    LocalMux I__4976 (
            .O(N__31003),
            .I(n2484));
    CascadeMux I__4975 (
            .O(N__31000),
            .I(N__30997));
    InMux I__4974 (
            .O(N__30997),
            .I(N__30994));
    LocalMux I__4973 (
            .O(N__30994),
            .I(N__30990));
    InMux I__4972 (
            .O(N__30993),
            .I(N__30987));
    Span4Mux_v I__4971 (
            .O(N__30990),
            .I(N__30984));
    LocalMux I__4970 (
            .O(N__30987),
            .I(N__30981));
    Span4Mux_h I__4969 (
            .O(N__30984),
            .I(N__30976));
    Span4Mux_h I__4968 (
            .O(N__30981),
            .I(N__30976));
    Odrv4 I__4967 (
            .O(N__30976),
            .I(n2516));
    InMux I__4966 (
            .O(N__30973),
            .I(N__30968));
    InMux I__4965 (
            .O(N__30972),
            .I(N__30965));
    InMux I__4964 (
            .O(N__30971),
            .I(N__30962));
    LocalMux I__4963 (
            .O(N__30968),
            .I(N__30959));
    LocalMux I__4962 (
            .O(N__30965),
            .I(N__30954));
    LocalMux I__4961 (
            .O(N__30962),
            .I(N__30954));
    Span4Mux_v I__4960 (
            .O(N__30959),
            .I(N__30951));
    Odrv4 I__4959 (
            .O(N__30954),
            .I(n2514));
    Odrv4 I__4958 (
            .O(N__30951),
            .I(n2514));
    CascadeMux I__4957 (
            .O(N__30946),
            .I(n2516_cascade_));
    InMux I__4956 (
            .O(N__30943),
            .I(N__30940));
    LocalMux I__4955 (
            .O(N__30940),
            .I(N__30937));
    Odrv4 I__4954 (
            .O(N__30937),
            .I(n13810));
    CascadeMux I__4953 (
            .O(N__30934),
            .I(n13816_cascade_));
    InMux I__4952 (
            .O(N__30931),
            .I(N__30928));
    LocalMux I__4951 (
            .O(N__30928),
            .I(N__30924));
    InMux I__4950 (
            .O(N__30927),
            .I(N__30921));
    Odrv12 I__4949 (
            .O(N__30924),
            .I(n2511));
    LocalMux I__4948 (
            .O(N__30921),
            .I(n2511));
    InMux I__4947 (
            .O(N__30916),
            .I(N__30913));
    LocalMux I__4946 (
            .O(N__30913),
            .I(N__30910));
    Odrv4 I__4945 (
            .O(N__30910),
            .I(n2582));
    CascadeMux I__4944 (
            .O(N__30907),
            .I(n2544_cascade_));
    CascadeMux I__4943 (
            .O(N__30904),
            .I(N__30901));
    InMux I__4942 (
            .O(N__30901),
            .I(N__30898));
    LocalMux I__4941 (
            .O(N__30898),
            .I(N__30895));
    Odrv4 I__4940 (
            .O(N__30895),
            .I(n2579));
    InMux I__4939 (
            .O(N__30892),
            .I(N__30888));
    CascadeMux I__4938 (
            .O(N__30891),
            .I(N__30885));
    LocalMux I__4937 (
            .O(N__30888),
            .I(N__30881));
    InMux I__4936 (
            .O(N__30885),
            .I(N__30878));
    InMux I__4935 (
            .O(N__30884),
            .I(N__30875));
    Span4Mux_v I__4934 (
            .O(N__30881),
            .I(N__30872));
    LocalMux I__4933 (
            .O(N__30878),
            .I(N__30869));
    LocalMux I__4932 (
            .O(N__30875),
            .I(N__30866));
    Odrv4 I__4931 (
            .O(N__30872),
            .I(n2425));
    Odrv4 I__4930 (
            .O(N__30869),
            .I(n2425));
    Odrv4 I__4929 (
            .O(N__30866),
            .I(n2425));
    InMux I__4928 (
            .O(N__30859),
            .I(N__30856));
    LocalMux I__4927 (
            .O(N__30856),
            .I(n2492));
    CascadeMux I__4926 (
            .O(N__30853),
            .I(N__30849));
    InMux I__4925 (
            .O(N__30852),
            .I(N__30846));
    InMux I__4924 (
            .O(N__30849),
            .I(N__30843));
    LocalMux I__4923 (
            .O(N__30846),
            .I(N__30840));
    LocalMux I__4922 (
            .O(N__30843),
            .I(N__30837));
    Span4Mux_h I__4921 (
            .O(N__30840),
            .I(N__30834));
    Odrv4 I__4920 (
            .O(N__30837),
            .I(n2524));
    Odrv4 I__4919 (
            .O(N__30834),
            .I(n2524));
    InMux I__4918 (
            .O(N__30829),
            .I(N__30826));
    LocalMux I__4917 (
            .O(N__30826),
            .I(n2590));
    InMux I__4916 (
            .O(N__30823),
            .I(N__30820));
    LocalMux I__4915 (
            .O(N__30820),
            .I(N__30817));
    Odrv4 I__4914 (
            .O(N__30817),
            .I(n2592));
    CascadeMux I__4913 (
            .O(N__30814),
            .I(N__30810));
    CascadeMux I__4912 (
            .O(N__30813),
            .I(N__30807));
    InMux I__4911 (
            .O(N__30810),
            .I(N__30804));
    InMux I__4910 (
            .O(N__30807),
            .I(N__30801));
    LocalMux I__4909 (
            .O(N__30804),
            .I(N__30797));
    LocalMux I__4908 (
            .O(N__30801),
            .I(N__30794));
    InMux I__4907 (
            .O(N__30800),
            .I(N__30791));
    Odrv4 I__4906 (
            .O(N__30797),
            .I(n2525));
    Odrv4 I__4905 (
            .O(N__30794),
            .I(n2525));
    LocalMux I__4904 (
            .O(N__30791),
            .I(n2525));
    InMux I__4903 (
            .O(N__30784),
            .I(N__30780));
    CascadeMux I__4902 (
            .O(N__30783),
            .I(N__30777));
    LocalMux I__4901 (
            .O(N__30780),
            .I(N__30774));
    InMux I__4900 (
            .O(N__30777),
            .I(N__30771));
    Span4Mux_v I__4899 (
            .O(N__30774),
            .I(N__30768));
    LocalMux I__4898 (
            .O(N__30771),
            .I(N__30765));
    Odrv4 I__4897 (
            .O(N__30768),
            .I(n2517));
    Odrv4 I__4896 (
            .O(N__30765),
            .I(n2517));
    InMux I__4895 (
            .O(N__30760),
            .I(N__30757));
    LocalMux I__4894 (
            .O(N__30757),
            .I(n2584));
    InMux I__4893 (
            .O(N__30754),
            .I(N__30751));
    LocalMux I__4892 (
            .O(N__30751),
            .I(N__30748));
    Odrv4 I__4891 (
            .O(N__30748),
            .I(n2595));
    CascadeMux I__4890 (
            .O(N__30745),
            .I(N__30741));
    CascadeMux I__4889 (
            .O(N__30744),
            .I(N__30738));
    InMux I__4888 (
            .O(N__30741),
            .I(N__30735));
    InMux I__4887 (
            .O(N__30738),
            .I(N__30732));
    LocalMux I__4886 (
            .O(N__30735),
            .I(N__30729));
    LocalMux I__4885 (
            .O(N__30732),
            .I(N__30725));
    Span4Mux_h I__4884 (
            .O(N__30729),
            .I(N__30722));
    InMux I__4883 (
            .O(N__30728),
            .I(N__30719));
    Odrv4 I__4882 (
            .O(N__30725),
            .I(n2528));
    Odrv4 I__4881 (
            .O(N__30722),
            .I(n2528));
    LocalMux I__4880 (
            .O(N__30719),
            .I(n2528));
    InMux I__4879 (
            .O(N__30712),
            .I(N__30709));
    LocalMux I__4878 (
            .O(N__30709),
            .I(n2491));
    CascadeMux I__4877 (
            .O(N__30706),
            .I(N__30703));
    InMux I__4876 (
            .O(N__30703),
            .I(N__30700));
    LocalMux I__4875 (
            .O(N__30700),
            .I(N__30696));
    CascadeMux I__4874 (
            .O(N__30699),
            .I(N__30693));
    Span4Mux_v I__4873 (
            .O(N__30696),
            .I(N__30690));
    InMux I__4872 (
            .O(N__30693),
            .I(N__30687));
    Span4Mux_h I__4871 (
            .O(N__30690),
            .I(N__30682));
    LocalMux I__4870 (
            .O(N__30687),
            .I(N__30682));
    Span4Mux_h I__4869 (
            .O(N__30682),
            .I(N__30678));
    InMux I__4868 (
            .O(N__30681),
            .I(N__30675));
    Odrv4 I__4867 (
            .O(N__30678),
            .I(n2424));
    LocalMux I__4866 (
            .O(N__30675),
            .I(n2424));
    CascadeMux I__4865 (
            .O(N__30670),
            .I(N__30666));
    CascadeMux I__4864 (
            .O(N__30669),
            .I(N__30662));
    InMux I__4863 (
            .O(N__30666),
            .I(N__30659));
    InMux I__4862 (
            .O(N__30665),
            .I(N__30656));
    InMux I__4861 (
            .O(N__30662),
            .I(N__30653));
    LocalMux I__4860 (
            .O(N__30659),
            .I(N__30650));
    LocalMux I__4859 (
            .O(N__30656),
            .I(N__30647));
    LocalMux I__4858 (
            .O(N__30653),
            .I(n2523));
    Odrv4 I__4857 (
            .O(N__30650),
            .I(n2523));
    Odrv4 I__4856 (
            .O(N__30647),
            .I(n2523));
    InMux I__4855 (
            .O(N__30640),
            .I(N__30637));
    LocalMux I__4854 (
            .O(N__30637),
            .I(N__30634));
    Span4Mux_v I__4853 (
            .O(N__30634),
            .I(N__30631));
    Odrv4 I__4852 (
            .O(N__30631),
            .I(n2583));
    InMux I__4851 (
            .O(N__30628),
            .I(N__30625));
    LocalMux I__4850 (
            .O(N__30625),
            .I(N__30622));
    Odrv4 I__4849 (
            .O(N__30622),
            .I(n2596));
    CascadeMux I__4848 (
            .O(N__30619),
            .I(N__30615));
    InMux I__4847 (
            .O(N__30618),
            .I(N__30612));
    InMux I__4846 (
            .O(N__30615),
            .I(N__30609));
    LocalMux I__4845 (
            .O(N__30612),
            .I(N__30606));
    LocalMux I__4844 (
            .O(N__30609),
            .I(N__30603));
    Span4Mux_h I__4843 (
            .O(N__30606),
            .I(N__30597));
    Span4Mux_v I__4842 (
            .O(N__30603),
            .I(N__30597));
    InMux I__4841 (
            .O(N__30602),
            .I(N__30594));
    Odrv4 I__4840 (
            .O(N__30597),
            .I(n2529));
    LocalMux I__4839 (
            .O(N__30594),
            .I(n2529));
    InMux I__4838 (
            .O(N__30589),
            .I(n12118));
    InMux I__4837 (
            .O(N__30586),
            .I(N__30583));
    LocalMux I__4836 (
            .O(N__30583),
            .I(n1095));
    InMux I__4835 (
            .O(N__30580),
            .I(n12119));
    InMux I__4834 (
            .O(N__30577),
            .I(N__30574));
    LocalMux I__4833 (
            .O(N__30574),
            .I(n1094));
    InMux I__4832 (
            .O(N__30571),
            .I(n12120));
    InMux I__4831 (
            .O(N__30568),
            .I(bfn_6_32_0_));
    InMux I__4830 (
            .O(N__30565),
            .I(N__30562));
    LocalMux I__4829 (
            .O(N__30562),
            .I(n1093));
    CascadeMux I__4828 (
            .O(N__30559),
            .I(N__30556));
    InMux I__4827 (
            .O(N__30556),
            .I(N__30553));
    LocalMux I__4826 (
            .O(N__30553),
            .I(n1096));
    CascadeMux I__4825 (
            .O(N__30550),
            .I(N__30547));
    InMux I__4824 (
            .O(N__30547),
            .I(N__30544));
    LocalMux I__4823 (
            .O(N__30544),
            .I(N__30540));
    CascadeMux I__4822 (
            .O(N__30543),
            .I(N__30537));
    Span4Mux_s2_h I__4821 (
            .O(N__30540),
            .I(N__30533));
    InMux I__4820 (
            .O(N__30537),
            .I(N__30530));
    InMux I__4819 (
            .O(N__30536),
            .I(N__30527));
    Span4Mux_h I__4818 (
            .O(N__30533),
            .I(N__30524));
    LocalMux I__4817 (
            .O(N__30530),
            .I(n1128));
    LocalMux I__4816 (
            .O(N__30527),
            .I(n1128));
    Odrv4 I__4815 (
            .O(N__30524),
            .I(n1128));
    CascadeMux I__4814 (
            .O(N__30517),
            .I(N__30513));
    CascadeMux I__4813 (
            .O(N__30516),
            .I(N__30510));
    InMux I__4812 (
            .O(N__30513),
            .I(N__30506));
    InMux I__4811 (
            .O(N__30510),
            .I(N__30503));
    InMux I__4810 (
            .O(N__30509),
            .I(N__30500));
    LocalMux I__4809 (
            .O(N__30506),
            .I(n1028));
    LocalMux I__4808 (
            .O(N__30503),
            .I(n1028));
    LocalMux I__4807 (
            .O(N__30500),
            .I(n1028));
    CascadeMux I__4806 (
            .O(N__30493),
            .I(N__30489));
    CascadeMux I__4805 (
            .O(N__30492),
            .I(N__30485));
    InMux I__4804 (
            .O(N__30489),
            .I(N__30482));
    InMux I__4803 (
            .O(N__30488),
            .I(N__30479));
    InMux I__4802 (
            .O(N__30485),
            .I(N__30476));
    LocalMux I__4801 (
            .O(N__30482),
            .I(N__30469));
    LocalMux I__4800 (
            .O(N__30479),
            .I(N__30469));
    LocalMux I__4799 (
            .O(N__30476),
            .I(N__30469));
    Odrv4 I__4798 (
            .O(N__30469),
            .I(n1027));
    CascadeMux I__4797 (
            .O(N__30466),
            .I(n1059_cascade_));
    InMux I__4796 (
            .O(N__30463),
            .I(N__30460));
    LocalMux I__4795 (
            .O(N__30460),
            .I(n1099));
    CascadeMux I__4794 (
            .O(N__30457),
            .I(N__30454));
    InMux I__4793 (
            .O(N__30454),
            .I(N__30450));
    CascadeMux I__4792 (
            .O(N__30453),
            .I(N__30446));
    LocalMux I__4791 (
            .O(N__30450),
            .I(N__30443));
    CascadeMux I__4790 (
            .O(N__30449),
            .I(N__30440));
    InMux I__4789 (
            .O(N__30446),
            .I(N__30437));
    Span4Mux_s1_h I__4788 (
            .O(N__30443),
            .I(N__30434));
    InMux I__4787 (
            .O(N__30440),
            .I(N__30431));
    LocalMux I__4786 (
            .O(N__30437),
            .I(N__30428));
    Span4Mux_h I__4785 (
            .O(N__30434),
            .I(N__30425));
    LocalMux I__4784 (
            .O(N__30431),
            .I(n1131));
    Odrv4 I__4783 (
            .O(N__30428),
            .I(n1131));
    Odrv4 I__4782 (
            .O(N__30425),
            .I(n1131));
    CascadeMux I__4781 (
            .O(N__30418),
            .I(N__30414));
    InMux I__4780 (
            .O(N__30417),
            .I(N__30411));
    InMux I__4779 (
            .O(N__30414),
            .I(N__30408));
    LocalMux I__4778 (
            .O(N__30411),
            .I(N__30402));
    LocalMux I__4777 (
            .O(N__30408),
            .I(N__30402));
    InMux I__4776 (
            .O(N__30407),
            .I(N__30399));
    Span4Mux_v I__4775 (
            .O(N__30402),
            .I(N__30396));
    LocalMux I__4774 (
            .O(N__30399),
            .I(encoder0_position_23));
    Odrv4 I__4773 (
            .O(N__30396),
            .I(encoder0_position_23));
    InMux I__4772 (
            .O(N__30391),
            .I(N__30386));
    CascadeMux I__4771 (
            .O(N__30390),
            .I(N__30383));
    InMux I__4770 (
            .O(N__30389),
            .I(N__30380));
    LocalMux I__4769 (
            .O(N__30386),
            .I(N__30377));
    InMux I__4768 (
            .O(N__30383),
            .I(N__30374));
    LocalMux I__4767 (
            .O(N__30380),
            .I(encoder0_position_24));
    Odrv12 I__4766 (
            .O(N__30377),
            .I(encoder0_position_24));
    LocalMux I__4765 (
            .O(N__30374),
            .I(encoder0_position_24));
    CascadeMux I__4764 (
            .O(N__30367),
            .I(N__30364));
    InMux I__4763 (
            .O(N__30364),
            .I(N__30361));
    LocalMux I__4762 (
            .O(N__30361),
            .I(n1101));
    InMux I__4761 (
            .O(N__30358),
            .I(bfn_6_31_0_));
    InMux I__4760 (
            .O(N__30355),
            .I(N__30352));
    LocalMux I__4759 (
            .O(N__30352),
            .I(n1100));
    InMux I__4758 (
            .O(N__30349),
            .I(n12114));
    InMux I__4757 (
            .O(N__30346),
            .I(n12115));
    InMux I__4756 (
            .O(N__30343),
            .I(N__30340));
    LocalMux I__4755 (
            .O(N__30340),
            .I(N__30337));
    Span4Mux_s1_v I__4754 (
            .O(N__30337),
            .I(N__30334));
    Odrv4 I__4753 (
            .O(N__30334),
            .I(n1098));
    InMux I__4752 (
            .O(N__30331),
            .I(n12116));
    InMux I__4751 (
            .O(N__30328),
            .I(N__30325));
    LocalMux I__4750 (
            .O(N__30325),
            .I(n1097));
    InMux I__4749 (
            .O(N__30322),
            .I(n12117));
    InMux I__4748 (
            .O(N__30319),
            .I(N__30314));
    CascadeMux I__4747 (
            .O(N__30318),
            .I(N__30311));
    CascadeMux I__4746 (
            .O(N__30317),
            .I(N__30308));
    LocalMux I__4745 (
            .O(N__30314),
            .I(N__30304));
    InMux I__4744 (
            .O(N__30311),
            .I(N__30301));
    InMux I__4743 (
            .O(N__30308),
            .I(N__30298));
    InMux I__4742 (
            .O(N__30307),
            .I(N__30295));
    Odrv4 I__4741 (
            .O(N__30304),
            .I(n13254));
    LocalMux I__4740 (
            .O(N__30301),
            .I(n13254));
    LocalMux I__4739 (
            .O(N__30298),
            .I(n13254));
    LocalMux I__4738 (
            .O(N__30295),
            .I(n13254));
    InMux I__4737 (
            .O(N__30286),
            .I(N__30283));
    LocalMux I__4736 (
            .O(N__30283),
            .I(n2286));
    CascadeMux I__4735 (
            .O(N__30280),
            .I(n13255_cascade_));
    CascadeMux I__4734 (
            .O(N__30277),
            .I(N__30273));
    InMux I__4733 (
            .O(N__30276),
            .I(N__30268));
    InMux I__4732 (
            .O(N__30273),
            .I(N__30263));
    InMux I__4731 (
            .O(N__30272),
            .I(N__30263));
    InMux I__4730 (
            .O(N__30271),
            .I(N__30260));
    LocalMux I__4729 (
            .O(N__30268),
            .I(N__30255));
    LocalMux I__4728 (
            .O(N__30263),
            .I(N__30255));
    LocalMux I__4727 (
            .O(N__30260),
            .I(encoder0_position_26));
    Odrv4 I__4726 (
            .O(N__30255),
            .I(encoder0_position_26));
    CascadeMux I__4725 (
            .O(N__30250),
            .I(N__30246));
    InMux I__4724 (
            .O(N__30249),
            .I(N__30240));
    InMux I__4723 (
            .O(N__30246),
            .I(N__30240));
    InMux I__4722 (
            .O(N__30245),
            .I(N__30236));
    LocalMux I__4721 (
            .O(N__30240),
            .I(N__30233));
    InMux I__4720 (
            .O(N__30239),
            .I(N__30230));
    LocalMux I__4719 (
            .O(N__30236),
            .I(encoder0_position_30));
    Odrv4 I__4718 (
            .O(N__30233),
            .I(encoder0_position_30));
    LocalMux I__4717 (
            .O(N__30230),
            .I(encoder0_position_30));
    CascadeMux I__4716 (
            .O(N__30223),
            .I(N__30220));
    InMux I__4715 (
            .O(N__30220),
            .I(N__30217));
    LocalMux I__4714 (
            .O(N__30217),
            .I(n403));
    CascadeMux I__4713 (
            .O(N__30214),
            .I(n11712_cascade_));
    CascadeMux I__4712 (
            .O(N__30211),
            .I(n861_cascade_));
    CascadeMux I__4711 (
            .O(N__30208),
            .I(n14170_cascade_));
    InMux I__4710 (
            .O(N__30205),
            .I(N__30202));
    LocalMux I__4709 (
            .O(N__30202),
            .I(n2285));
    CascadeMux I__4708 (
            .O(N__30199),
            .I(N__30196));
    InMux I__4707 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__4706 (
            .O(N__30193),
            .I(n293));
    CascadeMux I__4705 (
            .O(N__30190),
            .I(n293_cascade_));
    InMux I__4704 (
            .O(N__30187),
            .I(N__30184));
    LocalMux I__4703 (
            .O(N__30184),
            .I(n5_adj_697));
    CascadeMux I__4702 (
            .O(N__30181),
            .I(n5_adj_697_cascade_));
    InMux I__4701 (
            .O(N__30178),
            .I(N__30175));
    LocalMux I__4700 (
            .O(N__30175),
            .I(n2290));
    CascadeMux I__4699 (
            .O(N__30172),
            .I(n13254_cascade_));
    InMux I__4698 (
            .O(N__30169),
            .I(N__30166));
    LocalMux I__4697 (
            .O(N__30166),
            .I(n13259));
    InMux I__4696 (
            .O(N__30163),
            .I(N__30160));
    LocalMux I__4695 (
            .O(N__30160),
            .I(n13263));
    CascadeMux I__4694 (
            .O(N__30157),
            .I(N__30154));
    InMux I__4693 (
            .O(N__30154),
            .I(N__30151));
    LocalMux I__4692 (
            .O(N__30151),
            .I(n174));
    InMux I__4691 (
            .O(N__30148),
            .I(\quad_counter0.n12653 ));
    CascadeMux I__4690 (
            .O(N__30145),
            .I(N__30141));
    InMux I__4689 (
            .O(N__30144),
            .I(N__30137));
    InMux I__4688 (
            .O(N__30141),
            .I(N__30134));
    InMux I__4687 (
            .O(N__30140),
            .I(N__30131));
    LocalMux I__4686 (
            .O(N__30137),
            .I(N__30128));
    LocalMux I__4685 (
            .O(N__30134),
            .I(encoder0_position_16));
    LocalMux I__4684 (
            .O(N__30131),
            .I(encoder0_position_16));
    Odrv4 I__4683 (
            .O(N__30128),
            .I(encoder0_position_16));
    InMux I__4682 (
            .O(N__30121),
            .I(N__30117));
    CascadeMux I__4681 (
            .O(N__30120),
            .I(N__30113));
    LocalMux I__4680 (
            .O(N__30117),
            .I(N__30110));
    CascadeMux I__4679 (
            .O(N__30116),
            .I(N__30107));
    InMux I__4678 (
            .O(N__30113),
            .I(N__30103));
    Span4Mux_v I__4677 (
            .O(N__30110),
            .I(N__30100));
    InMux I__4676 (
            .O(N__30107),
            .I(N__30097));
    InMux I__4675 (
            .O(N__30106),
            .I(N__30094));
    LocalMux I__4674 (
            .O(N__30103),
            .I(encoder0_position_27));
    Odrv4 I__4673 (
            .O(N__30100),
            .I(encoder0_position_27));
    LocalMux I__4672 (
            .O(N__30097),
            .I(encoder0_position_27));
    LocalMux I__4671 (
            .O(N__30094),
            .I(encoder0_position_27));
    CascadeMux I__4670 (
            .O(N__30085),
            .I(N__30082));
    InMux I__4669 (
            .O(N__30082),
            .I(N__30079));
    LocalMux I__4668 (
            .O(N__30079),
            .I(n175));
    CascadeMux I__4667 (
            .O(N__30076),
            .I(N__30072));
    CascadeMux I__4666 (
            .O(N__30075),
            .I(N__30069));
    InMux I__4665 (
            .O(N__30072),
            .I(N__30065));
    InMux I__4664 (
            .O(N__30069),
            .I(N__30061));
    InMux I__4663 (
            .O(N__30068),
            .I(N__30058));
    LocalMux I__4662 (
            .O(N__30065),
            .I(N__30055));
    InMux I__4661 (
            .O(N__30064),
            .I(N__30052));
    LocalMux I__4660 (
            .O(N__30061),
            .I(encoder0_position_29));
    LocalMux I__4659 (
            .O(N__30058),
            .I(encoder0_position_29));
    Odrv4 I__4658 (
            .O(N__30055),
            .I(encoder0_position_29));
    LocalMux I__4657 (
            .O(N__30052),
            .I(encoder0_position_29));
    InMux I__4656 (
            .O(N__30043),
            .I(N__30040));
    LocalMux I__4655 (
            .O(N__30040),
            .I(n404));
    InMux I__4654 (
            .O(N__30037),
            .I(N__30030));
    InMux I__4653 (
            .O(N__30036),
            .I(N__30030));
    CascadeMux I__4652 (
            .O(N__30035),
            .I(N__30027));
    LocalMux I__4651 (
            .O(N__30030),
            .I(N__30024));
    InMux I__4650 (
            .O(N__30027),
            .I(N__30021));
    Span4Mux_v I__4649 (
            .O(N__30024),
            .I(N__30018));
    LocalMux I__4648 (
            .O(N__30021),
            .I(encoder0_position_22));
    Odrv4 I__4647 (
            .O(N__30018),
            .I(encoder0_position_22));
    InMux I__4646 (
            .O(N__30013),
            .I(\quad_counter0.n12644 ));
    InMux I__4645 (
            .O(N__30010),
            .I(\quad_counter0.n12645 ));
    InMux I__4644 (
            .O(N__30007),
            .I(bfn_6_26_0_));
    InMux I__4643 (
            .O(N__30004),
            .I(\quad_counter0.n12647 ));
    InMux I__4642 (
            .O(N__30001),
            .I(\quad_counter0.n12648 ));
    InMux I__4641 (
            .O(N__29998),
            .I(\quad_counter0.n12649 ));
    InMux I__4640 (
            .O(N__29995),
            .I(\quad_counter0.n12650 ));
    InMux I__4639 (
            .O(N__29992),
            .I(\quad_counter0.n12651 ));
    InMux I__4638 (
            .O(N__29989),
            .I(\quad_counter0.n12652 ));
    InMux I__4637 (
            .O(N__29986),
            .I(\quad_counter0.n12636 ));
    InMux I__4636 (
            .O(N__29983),
            .I(\quad_counter0.n12637 ));
    InMux I__4635 (
            .O(N__29980),
            .I(bfn_6_25_0_));
    InMux I__4634 (
            .O(N__29977),
            .I(N__29970));
    InMux I__4633 (
            .O(N__29976),
            .I(N__29970));
    InMux I__4632 (
            .O(N__29975),
            .I(N__29967));
    LocalMux I__4631 (
            .O(N__29970),
            .I(N__29964));
    LocalMux I__4630 (
            .O(N__29967),
            .I(encoder0_position_17));
    Odrv4 I__4629 (
            .O(N__29964),
            .I(encoder0_position_17));
    InMux I__4628 (
            .O(N__29959),
            .I(\quad_counter0.n12639 ));
    CascadeMux I__4627 (
            .O(N__29956),
            .I(N__29952));
    InMux I__4626 (
            .O(N__29955),
            .I(N__29948));
    InMux I__4625 (
            .O(N__29952),
            .I(N__29945));
    InMux I__4624 (
            .O(N__29951),
            .I(N__29942));
    LocalMux I__4623 (
            .O(N__29948),
            .I(N__29939));
    LocalMux I__4622 (
            .O(N__29945),
            .I(encoder0_position_18));
    LocalMux I__4621 (
            .O(N__29942),
            .I(encoder0_position_18));
    Odrv4 I__4620 (
            .O(N__29939),
            .I(encoder0_position_18));
    InMux I__4619 (
            .O(N__29932),
            .I(\quad_counter0.n12640 ));
    InMux I__4618 (
            .O(N__29929),
            .I(N__29923));
    InMux I__4617 (
            .O(N__29928),
            .I(N__29923));
    LocalMux I__4616 (
            .O(N__29923),
            .I(N__29919));
    InMux I__4615 (
            .O(N__29922),
            .I(N__29916));
    Span4Mux_v I__4614 (
            .O(N__29919),
            .I(N__29913));
    LocalMux I__4613 (
            .O(N__29916),
            .I(encoder0_position_19));
    Odrv4 I__4612 (
            .O(N__29913),
            .I(encoder0_position_19));
    InMux I__4611 (
            .O(N__29908),
            .I(\quad_counter0.n12641 ));
    InMux I__4610 (
            .O(N__29905),
            .I(N__29902));
    LocalMux I__4609 (
            .O(N__29902),
            .I(N__29898));
    CascadeMux I__4608 (
            .O(N__29901),
            .I(N__29894));
    Span4Mux_h I__4607 (
            .O(N__29898),
            .I(N__29891));
    InMux I__4606 (
            .O(N__29897),
            .I(N__29888));
    InMux I__4605 (
            .O(N__29894),
            .I(N__29885));
    Span4Mux_v I__4604 (
            .O(N__29891),
            .I(N__29880));
    LocalMux I__4603 (
            .O(N__29888),
            .I(N__29880));
    LocalMux I__4602 (
            .O(N__29885),
            .I(encoder0_position_20));
    Odrv4 I__4601 (
            .O(N__29880),
            .I(encoder0_position_20));
    InMux I__4600 (
            .O(N__29875),
            .I(\quad_counter0.n12642 ));
    InMux I__4599 (
            .O(N__29872),
            .I(N__29866));
    InMux I__4598 (
            .O(N__29871),
            .I(N__29866));
    LocalMux I__4597 (
            .O(N__29866),
            .I(N__29862));
    InMux I__4596 (
            .O(N__29865),
            .I(N__29859));
    Span4Mux_v I__4595 (
            .O(N__29862),
            .I(N__29856));
    LocalMux I__4594 (
            .O(N__29859),
            .I(encoder0_position_21));
    Odrv4 I__4593 (
            .O(N__29856),
            .I(encoder0_position_21));
    InMux I__4592 (
            .O(N__29851),
            .I(\quad_counter0.n12643 ));
    InMux I__4591 (
            .O(N__29848),
            .I(\quad_counter0.n12627 ));
    InMux I__4590 (
            .O(N__29845),
            .I(\quad_counter0.n12628 ));
    InMux I__4589 (
            .O(N__29842),
            .I(\quad_counter0.n12629 ));
    InMux I__4588 (
            .O(N__29839),
            .I(bfn_6_24_0_));
    InMux I__4587 (
            .O(N__29836),
            .I(\quad_counter0.n12631 ));
    InMux I__4586 (
            .O(N__29833),
            .I(\quad_counter0.n12632 ));
    InMux I__4585 (
            .O(N__29830),
            .I(\quad_counter0.n12633 ));
    CascadeMux I__4584 (
            .O(N__29827),
            .I(N__29823));
    InMux I__4583 (
            .O(N__29826),
            .I(N__29820));
    InMux I__4582 (
            .O(N__29823),
            .I(N__29816));
    LocalMux I__4581 (
            .O(N__29820),
            .I(N__29813));
    InMux I__4580 (
            .O(N__29819),
            .I(N__29810));
    LocalMux I__4579 (
            .O(N__29816),
            .I(encoder0_position_12));
    Odrv4 I__4578 (
            .O(N__29813),
            .I(encoder0_position_12));
    LocalMux I__4577 (
            .O(N__29810),
            .I(encoder0_position_12));
    InMux I__4576 (
            .O(N__29803),
            .I(\quad_counter0.n12634 ));
    InMux I__4575 (
            .O(N__29800),
            .I(\quad_counter0.n12635 ));
    InMux I__4574 (
            .O(N__29797),
            .I(N__29794));
    LocalMux I__4573 (
            .O(N__29794),
            .I(N__29791));
    Span4Mux_h I__4572 (
            .O(N__29791),
            .I(N__29788));
    Odrv4 I__4571 (
            .O(N__29788),
            .I(n2382));
    CascadeMux I__4570 (
            .O(N__29785),
            .I(n2315_cascade_));
    InMux I__4569 (
            .O(N__29782),
            .I(N__29778));
    InMux I__4568 (
            .O(N__29781),
            .I(N__29775));
    LocalMux I__4567 (
            .O(N__29778),
            .I(N__29772));
    LocalMux I__4566 (
            .O(N__29775),
            .I(N__29767));
    Span4Mux_h I__4565 (
            .O(N__29772),
            .I(N__29767));
    Odrv4 I__4564 (
            .O(N__29767),
            .I(n2414));
    CascadeMux I__4563 (
            .O(N__29764),
            .I(n2414_cascade_));
    InMux I__4562 (
            .O(N__29761),
            .I(N__29758));
    LocalMux I__4561 (
            .O(N__29758),
            .I(N__29755));
    Odrv4 I__4560 (
            .O(N__29755),
            .I(n2481));
    InMux I__4559 (
            .O(N__29752),
            .I(bfn_6_23_0_));
    InMux I__4558 (
            .O(N__29749),
            .I(\quad_counter0.n12623 ));
    InMux I__4557 (
            .O(N__29746),
            .I(\quad_counter0.n12624 ));
    InMux I__4556 (
            .O(N__29743),
            .I(\quad_counter0.n12625 ));
    InMux I__4555 (
            .O(N__29740),
            .I(\quad_counter0.n12626 ));
    CascadeMux I__4554 (
            .O(N__29737),
            .I(n11682_cascade_));
    InMux I__4553 (
            .O(N__29734),
            .I(N__29731));
    LocalMux I__4552 (
            .O(N__29731),
            .I(N__29728));
    Odrv4 I__4551 (
            .O(N__29728),
            .I(n13397));
    InMux I__4550 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__4549 (
            .O(N__29722),
            .I(N__29719));
    Odrv12 I__4548 (
            .O(N__29719),
            .I(n2086));
    CascadeMux I__4547 (
            .O(N__29716),
            .I(N__29713));
    InMux I__4546 (
            .O(N__29713),
            .I(N__29709));
    InMux I__4545 (
            .O(N__29712),
            .I(N__29706));
    LocalMux I__4544 (
            .O(N__29709),
            .I(N__29700));
    LocalMux I__4543 (
            .O(N__29706),
            .I(N__29700));
    InMux I__4542 (
            .O(N__29705),
            .I(N__29697));
    Odrv12 I__4541 (
            .O(N__29700),
            .I(n2019));
    LocalMux I__4540 (
            .O(N__29697),
            .I(n2019));
    InMux I__4539 (
            .O(N__29692),
            .I(N__29688));
    InMux I__4538 (
            .O(N__29691),
            .I(N__29685));
    LocalMux I__4537 (
            .O(N__29688),
            .I(N__29682));
    LocalMux I__4536 (
            .O(N__29685),
            .I(N__29677));
    Span4Mux_s1_h I__4535 (
            .O(N__29682),
            .I(N__29677));
    Span4Mux_h I__4534 (
            .O(N__29677),
            .I(N__29673));
    InMux I__4533 (
            .O(N__29676),
            .I(N__29670));
    Odrv4 I__4532 (
            .O(N__29673),
            .I(n2118));
    LocalMux I__4531 (
            .O(N__29670),
            .I(n2118));
    CascadeMux I__4530 (
            .O(N__29665),
            .I(N__29662));
    InMux I__4529 (
            .O(N__29662),
            .I(N__29658));
    InMux I__4528 (
            .O(N__29661),
            .I(N__29654));
    LocalMux I__4527 (
            .O(N__29658),
            .I(N__29651));
    InMux I__4526 (
            .O(N__29657),
            .I(N__29648));
    LocalMux I__4525 (
            .O(N__29654),
            .I(n2432));
    Odrv4 I__4524 (
            .O(N__29651),
            .I(n2432));
    LocalMux I__4523 (
            .O(N__29648),
            .I(n2432));
    CascadeMux I__4522 (
            .O(N__29641),
            .I(N__29638));
    InMux I__4521 (
            .O(N__29638),
            .I(N__29635));
    LocalMux I__4520 (
            .O(N__29635),
            .I(N__29632));
    Span4Mux_v I__4519 (
            .O(N__29632),
            .I(N__29629));
    Odrv4 I__4518 (
            .O(N__29629),
            .I(n2499));
    InMux I__4517 (
            .O(N__29626),
            .I(N__29622));
    InMux I__4516 (
            .O(N__29625),
            .I(N__29619));
    LocalMux I__4515 (
            .O(N__29622),
            .I(N__29616));
    LocalMux I__4514 (
            .O(N__29619),
            .I(N__29612));
    Span4Mux_v I__4513 (
            .O(N__29616),
            .I(N__29609));
    InMux I__4512 (
            .O(N__29615),
            .I(N__29606));
    Odrv4 I__4511 (
            .O(N__29612),
            .I(n2025));
    Odrv4 I__4510 (
            .O(N__29609),
            .I(n2025));
    LocalMux I__4509 (
            .O(N__29606),
            .I(n2025));
    CascadeMux I__4508 (
            .O(N__29599),
            .I(N__29596));
    InMux I__4507 (
            .O(N__29596),
            .I(N__29593));
    LocalMux I__4506 (
            .O(N__29593),
            .I(N__29590));
    Span4Mux_h I__4505 (
            .O(N__29590),
            .I(N__29587));
    Span4Mux_h I__4504 (
            .O(N__29587),
            .I(N__29584));
    Odrv4 I__4503 (
            .O(N__29584),
            .I(n2092));
    CascadeMux I__4502 (
            .O(N__29581),
            .I(N__29578));
    InMux I__4501 (
            .O(N__29578),
            .I(N__29575));
    LocalMux I__4500 (
            .O(N__29575),
            .I(N__29572));
    Span12Mux_s5_h I__4499 (
            .O(N__29572),
            .I(N__29568));
    InMux I__4498 (
            .O(N__29571),
            .I(N__29565));
    Odrv12 I__4497 (
            .O(N__29568),
            .I(n2124));
    LocalMux I__4496 (
            .O(N__29565),
            .I(n2124));
    InMux I__4495 (
            .O(N__29560),
            .I(N__29557));
    LocalMux I__4494 (
            .O(N__29557),
            .I(N__29554));
    Span4Mux_h I__4493 (
            .O(N__29554),
            .I(N__29551));
    Span4Mux_v I__4492 (
            .O(N__29551),
            .I(N__29548));
    Odrv4 I__4491 (
            .O(N__29548),
            .I(n2191));
    CascadeMux I__4490 (
            .O(N__29545),
            .I(n2124_cascade_));
    CascadeMux I__4489 (
            .O(N__29542),
            .I(n2223_cascade_));
    InMux I__4488 (
            .O(N__29539),
            .I(N__29535));
    InMux I__4487 (
            .O(N__29538),
            .I(N__29532));
    LocalMux I__4486 (
            .O(N__29535),
            .I(N__29527));
    LocalMux I__4485 (
            .O(N__29532),
            .I(N__29527));
    Span4Mux_h I__4484 (
            .O(N__29527),
            .I(N__29524));
    Odrv4 I__4483 (
            .O(N__29524),
            .I(n2315));
    InMux I__4482 (
            .O(N__29521),
            .I(N__29518));
    LocalMux I__4481 (
            .O(N__29518),
            .I(N__29515));
    Span4Mux_h I__4480 (
            .O(N__29515),
            .I(N__29512));
    Span4Mux_h I__4479 (
            .O(N__29512),
            .I(N__29509));
    Odrv4 I__4478 (
            .O(N__29509),
            .I(n2192));
    CascadeMux I__4477 (
            .O(N__29506),
            .I(N__29502));
    InMux I__4476 (
            .O(N__29505),
            .I(N__29498));
    InMux I__4475 (
            .O(N__29502),
            .I(N__29495));
    InMux I__4474 (
            .O(N__29501),
            .I(N__29492));
    LocalMux I__4473 (
            .O(N__29498),
            .I(N__29489));
    LocalMux I__4472 (
            .O(N__29495),
            .I(N__29486));
    LocalMux I__4471 (
            .O(N__29492),
            .I(N__29483));
    Span4Mux_h I__4470 (
            .O(N__29489),
            .I(N__29480));
    Odrv12 I__4469 (
            .O(N__29486),
            .I(n2125));
    Odrv4 I__4468 (
            .O(N__29483),
            .I(n2125));
    Odrv4 I__4467 (
            .O(N__29480),
            .I(n2125));
    CascadeMux I__4466 (
            .O(N__29473),
            .I(n2224_cascade_));
    CascadeMux I__4465 (
            .O(N__29470),
            .I(n14174_cascade_));
    CascadeMux I__4464 (
            .O(N__29467),
            .I(n14178_cascade_));
    InMux I__4463 (
            .O(N__29464),
            .I(N__29461));
    LocalMux I__4462 (
            .O(N__29461),
            .I(N__29458));
    Odrv4 I__4461 (
            .O(N__29458),
            .I(n14184));
    InMux I__4460 (
            .O(N__29455),
            .I(N__29452));
    LocalMux I__4459 (
            .O(N__29452),
            .I(N__29449));
    Odrv12 I__4458 (
            .O(N__29449),
            .I(n2500));
    CascadeMux I__4457 (
            .O(N__29446),
            .I(N__29442));
    CascadeMux I__4456 (
            .O(N__29445),
            .I(N__29439));
    InMux I__4455 (
            .O(N__29442),
            .I(N__29436));
    InMux I__4454 (
            .O(N__29439),
            .I(N__29433));
    LocalMux I__4453 (
            .O(N__29436),
            .I(N__29430));
    LocalMux I__4452 (
            .O(N__29433),
            .I(n2433));
    Odrv4 I__4451 (
            .O(N__29430),
            .I(n2433));
    InMux I__4450 (
            .O(N__29425),
            .I(N__29421));
    CascadeMux I__4449 (
            .O(N__29424),
            .I(N__29418));
    LocalMux I__4448 (
            .O(N__29421),
            .I(N__29415));
    InMux I__4447 (
            .O(N__29418),
            .I(N__29412));
    Span4Mux_v I__4446 (
            .O(N__29415),
            .I(N__29406));
    LocalMux I__4445 (
            .O(N__29412),
            .I(N__29406));
    InMux I__4444 (
            .O(N__29411),
            .I(N__29403));
    Odrv4 I__4443 (
            .O(N__29406),
            .I(n2431));
    LocalMux I__4442 (
            .O(N__29403),
            .I(n2431));
    InMux I__4441 (
            .O(N__29398),
            .I(N__29395));
    LocalMux I__4440 (
            .O(N__29395),
            .I(N__29392));
    Odrv4 I__4439 (
            .O(N__29392),
            .I(n2498));
    InMux I__4438 (
            .O(N__29389),
            .I(N__29386));
    LocalMux I__4437 (
            .O(N__29386),
            .I(N__29383));
    Span4Mux_h I__4436 (
            .O(N__29383),
            .I(N__29380));
    Span4Mux_h I__4435 (
            .O(N__29380),
            .I(N__29377));
    Odrv4 I__4434 (
            .O(N__29377),
            .I(n2194));
    CascadeMux I__4433 (
            .O(N__29374),
            .I(N__29371));
    InMux I__4432 (
            .O(N__29371),
            .I(N__29367));
    InMux I__4431 (
            .O(N__29370),
            .I(N__29363));
    LocalMux I__4430 (
            .O(N__29367),
            .I(N__29360));
    CascadeMux I__4429 (
            .O(N__29366),
            .I(N__29357));
    LocalMux I__4428 (
            .O(N__29363),
            .I(N__29354));
    Span4Mux_h I__4427 (
            .O(N__29360),
            .I(N__29351));
    InMux I__4426 (
            .O(N__29357),
            .I(N__29348));
    Span4Mux_v I__4425 (
            .O(N__29354),
            .I(N__29345));
    Odrv4 I__4424 (
            .O(N__29351),
            .I(n2127));
    LocalMux I__4423 (
            .O(N__29348),
            .I(n2127));
    Odrv4 I__4422 (
            .O(N__29345),
            .I(n2127));
    InMux I__4421 (
            .O(N__29338),
            .I(N__29335));
    LocalMux I__4420 (
            .O(N__29335),
            .I(N__29332));
    Span4Mux_v I__4419 (
            .O(N__29332),
            .I(N__29329));
    Odrv4 I__4418 (
            .O(N__29329),
            .I(n2501));
    CascadeMux I__4417 (
            .O(N__29326),
            .I(n2533_cascade_));
    InMux I__4416 (
            .O(N__29323),
            .I(N__29316));
    InMux I__4415 (
            .O(N__29322),
            .I(N__29316));
    InMux I__4414 (
            .O(N__29321),
            .I(N__29313));
    LocalMux I__4413 (
            .O(N__29316),
            .I(N__29310));
    LocalMux I__4412 (
            .O(N__29313),
            .I(N__29307));
    Span4Mux_h I__4411 (
            .O(N__29310),
            .I(N__29304));
    Odrv12 I__4410 (
            .O(N__29307),
            .I(n2418));
    Odrv4 I__4409 (
            .O(N__29304),
            .I(n2418));
    InMux I__4408 (
            .O(N__29299),
            .I(N__29296));
    LocalMux I__4407 (
            .O(N__29296),
            .I(n2485));
    InMux I__4406 (
            .O(N__29293),
            .I(bfn_6_19_0_));
    InMux I__4405 (
            .O(N__29290),
            .I(n12333));
    InMux I__4404 (
            .O(N__29287),
            .I(n12334));
    CascadeMux I__4403 (
            .O(N__29284),
            .I(N__29281));
    InMux I__4402 (
            .O(N__29281),
            .I(N__29276));
    InMux I__4401 (
            .O(N__29280),
            .I(N__29273));
    InMux I__4400 (
            .O(N__29279),
            .I(N__29270));
    LocalMux I__4399 (
            .O(N__29276),
            .I(n2415));
    LocalMux I__4398 (
            .O(N__29273),
            .I(n2415));
    LocalMux I__4397 (
            .O(N__29270),
            .I(n2415));
    InMux I__4396 (
            .O(N__29263),
            .I(N__29260));
    LocalMux I__4395 (
            .O(N__29260),
            .I(n2482));
    InMux I__4394 (
            .O(N__29257),
            .I(n12335));
    InMux I__4393 (
            .O(N__29254),
            .I(n12336));
    InMux I__4392 (
            .O(N__29251),
            .I(n12337));
    InMux I__4391 (
            .O(N__29248),
            .I(N__29244));
    InMux I__4390 (
            .O(N__29247),
            .I(N__29241));
    LocalMux I__4389 (
            .O(N__29244),
            .I(N__29238));
    LocalMux I__4388 (
            .O(N__29241),
            .I(N__29235));
    Span4Mux_h I__4387 (
            .O(N__29238),
            .I(N__29232));
    Odrv12 I__4386 (
            .O(N__29235),
            .I(n2412));
    Odrv4 I__4385 (
            .O(N__29232),
            .I(n2412));
    InMux I__4384 (
            .O(N__29227),
            .I(n12338));
    CascadeMux I__4383 (
            .O(N__29224),
            .I(N__29220));
    InMux I__4382 (
            .O(N__29223),
            .I(N__29217));
    InMux I__4381 (
            .O(N__29220),
            .I(N__29214));
    LocalMux I__4380 (
            .O(N__29217),
            .I(N__29211));
    LocalMux I__4379 (
            .O(N__29214),
            .I(N__29208));
    Span4Mux_h I__4378 (
            .O(N__29211),
            .I(N__29204));
    Span4Mux_h I__4377 (
            .O(N__29208),
            .I(N__29201));
    InMux I__4376 (
            .O(N__29207),
            .I(N__29198));
    Odrv4 I__4375 (
            .O(N__29204),
            .I(n2421));
    Odrv4 I__4374 (
            .O(N__29201),
            .I(n2421));
    LocalMux I__4373 (
            .O(N__29198),
            .I(n2421));
    CascadeMux I__4372 (
            .O(N__29191),
            .I(N__29188));
    InMux I__4371 (
            .O(N__29188),
            .I(N__29185));
    LocalMux I__4370 (
            .O(N__29185),
            .I(n2488));
    InMux I__4369 (
            .O(N__29182),
            .I(N__29178));
    InMux I__4368 (
            .O(N__29181),
            .I(N__29174));
    LocalMux I__4367 (
            .O(N__29178),
            .I(N__29171));
    CascadeMux I__4366 (
            .O(N__29177),
            .I(N__29168));
    LocalMux I__4365 (
            .O(N__29174),
            .I(N__29165));
    Span4Mux_h I__4364 (
            .O(N__29171),
            .I(N__29162));
    InMux I__4363 (
            .O(N__29168),
            .I(N__29159));
    Span4Mux_v I__4362 (
            .O(N__29165),
            .I(N__29156));
    Odrv4 I__4361 (
            .O(N__29162),
            .I(n2126));
    LocalMux I__4360 (
            .O(N__29159),
            .I(n2126));
    Odrv4 I__4359 (
            .O(N__29156),
            .I(n2126));
    InMux I__4358 (
            .O(N__29149),
            .I(N__29146));
    LocalMux I__4357 (
            .O(N__29146),
            .I(N__29143));
    Span4Mux_h I__4356 (
            .O(N__29143),
            .I(N__29140));
    Span4Mux_h I__4355 (
            .O(N__29140),
            .I(N__29137));
    Odrv4 I__4354 (
            .O(N__29137),
            .I(n2193));
    InMux I__4353 (
            .O(N__29134),
            .I(N__29131));
    LocalMux I__4352 (
            .O(N__29131),
            .I(n2493));
    InMux I__4351 (
            .O(N__29128),
            .I(bfn_6_18_0_));
    InMux I__4350 (
            .O(N__29125),
            .I(n12325));
    InMux I__4349 (
            .O(N__29122),
            .I(n12326));
    InMux I__4348 (
            .O(N__29119),
            .I(N__29116));
    LocalMux I__4347 (
            .O(N__29116),
            .I(n2490));
    InMux I__4346 (
            .O(N__29113),
            .I(n12327));
    CascadeMux I__4345 (
            .O(N__29110),
            .I(N__29107));
    InMux I__4344 (
            .O(N__29107),
            .I(N__29102));
    InMux I__4343 (
            .O(N__29106),
            .I(N__29097));
    InMux I__4342 (
            .O(N__29105),
            .I(N__29097));
    LocalMux I__4341 (
            .O(N__29102),
            .I(n2422));
    LocalMux I__4340 (
            .O(N__29097),
            .I(n2422));
    InMux I__4339 (
            .O(N__29092),
            .I(N__29089));
    LocalMux I__4338 (
            .O(N__29089),
            .I(n2489));
    InMux I__4337 (
            .O(N__29086),
            .I(n12328));
    InMux I__4336 (
            .O(N__29083),
            .I(n12329));
    InMux I__4335 (
            .O(N__29080),
            .I(n12330));
    InMux I__4334 (
            .O(N__29077),
            .I(N__29074));
    LocalMux I__4333 (
            .O(N__29074),
            .I(N__29070));
    CascadeMux I__4332 (
            .O(N__29073),
            .I(N__29066));
    Span4Mux_h I__4331 (
            .O(N__29070),
            .I(N__29063));
    InMux I__4330 (
            .O(N__29069),
            .I(N__29058));
    InMux I__4329 (
            .O(N__29066),
            .I(N__29058));
    Odrv4 I__4328 (
            .O(N__29063),
            .I(n2419));
    LocalMux I__4327 (
            .O(N__29058),
            .I(n2419));
    InMux I__4326 (
            .O(N__29053),
            .I(N__29050));
    LocalMux I__4325 (
            .O(N__29050),
            .I(n2486));
    InMux I__4324 (
            .O(N__29047),
            .I(n12331));
    InMux I__4323 (
            .O(N__29044),
            .I(n12361));
    InMux I__4322 (
            .O(N__29041),
            .I(bfn_6_17_0_));
    InMux I__4321 (
            .O(N__29038),
            .I(n12317));
    InMux I__4320 (
            .O(N__29035),
            .I(n12318));
    InMux I__4319 (
            .O(N__29032),
            .I(n12319));
    CascadeMux I__4318 (
            .O(N__29029),
            .I(N__29026));
    InMux I__4317 (
            .O(N__29026),
            .I(N__29022));
    InMux I__4316 (
            .O(N__29025),
            .I(N__29019));
    LocalMux I__4315 (
            .O(N__29022),
            .I(N__29015));
    LocalMux I__4314 (
            .O(N__29019),
            .I(N__29012));
    InMux I__4313 (
            .O(N__29018),
            .I(N__29009));
    Span4Mux_h I__4312 (
            .O(N__29015),
            .I(N__29006));
    Span4Mux_v I__4311 (
            .O(N__29012),
            .I(N__29001));
    LocalMux I__4310 (
            .O(N__29009),
            .I(N__29001));
    Odrv4 I__4309 (
            .O(N__29006),
            .I(n2430));
    Odrv4 I__4308 (
            .O(N__29001),
            .I(n2430));
    InMux I__4307 (
            .O(N__28996),
            .I(N__28993));
    LocalMux I__4306 (
            .O(N__28993),
            .I(N__28990));
    Odrv4 I__4305 (
            .O(N__28990),
            .I(n2497));
    InMux I__4304 (
            .O(N__28987),
            .I(n12320));
    CascadeMux I__4303 (
            .O(N__28984),
            .I(N__28981));
    InMux I__4302 (
            .O(N__28981),
            .I(N__28977));
    CascadeMux I__4301 (
            .O(N__28980),
            .I(N__28974));
    LocalMux I__4300 (
            .O(N__28977),
            .I(N__28971));
    InMux I__4299 (
            .O(N__28974),
            .I(N__28968));
    Span4Mux_v I__4298 (
            .O(N__28971),
            .I(N__28965));
    LocalMux I__4297 (
            .O(N__28968),
            .I(n2429));
    Odrv4 I__4296 (
            .O(N__28965),
            .I(n2429));
    InMux I__4295 (
            .O(N__28960),
            .I(N__28957));
    LocalMux I__4294 (
            .O(N__28957),
            .I(N__28954));
    Odrv4 I__4293 (
            .O(N__28954),
            .I(n2496));
    InMux I__4292 (
            .O(N__28951),
            .I(n12321));
    CascadeMux I__4291 (
            .O(N__28948),
            .I(N__28945));
    InMux I__4290 (
            .O(N__28945),
            .I(N__28942));
    LocalMux I__4289 (
            .O(N__28942),
            .I(N__28938));
    InMux I__4288 (
            .O(N__28941),
            .I(N__28934));
    Span4Mux_h I__4287 (
            .O(N__28938),
            .I(N__28931));
    InMux I__4286 (
            .O(N__28937),
            .I(N__28928));
    LocalMux I__4285 (
            .O(N__28934),
            .I(n2428));
    Odrv4 I__4284 (
            .O(N__28931),
            .I(n2428));
    LocalMux I__4283 (
            .O(N__28928),
            .I(n2428));
    InMux I__4282 (
            .O(N__28921),
            .I(N__28918));
    LocalMux I__4281 (
            .O(N__28918),
            .I(n2495));
    InMux I__4280 (
            .O(N__28915),
            .I(n12322));
    CascadeMux I__4279 (
            .O(N__28912),
            .I(N__28908));
    CascadeMux I__4278 (
            .O(N__28911),
            .I(N__28905));
    InMux I__4277 (
            .O(N__28908),
            .I(N__28902));
    InMux I__4276 (
            .O(N__28905),
            .I(N__28899));
    LocalMux I__4275 (
            .O(N__28902),
            .I(N__28896));
    LocalMux I__4274 (
            .O(N__28899),
            .I(N__28892));
    Span4Mux_v I__4273 (
            .O(N__28896),
            .I(N__28889));
    InMux I__4272 (
            .O(N__28895),
            .I(N__28886));
    Span4Mux_v I__4271 (
            .O(N__28892),
            .I(N__28883));
    Odrv4 I__4270 (
            .O(N__28889),
            .I(n2427));
    LocalMux I__4269 (
            .O(N__28886),
            .I(n2427));
    Odrv4 I__4268 (
            .O(N__28883),
            .I(n2427));
    InMux I__4267 (
            .O(N__28876),
            .I(N__28873));
    LocalMux I__4266 (
            .O(N__28873),
            .I(n2494));
    InMux I__4265 (
            .O(N__28870),
            .I(n12323));
    InMux I__4264 (
            .O(N__28867),
            .I(n12352));
    InMux I__4263 (
            .O(N__28864),
            .I(n12353));
    InMux I__4262 (
            .O(N__28861),
            .I(bfn_6_16_0_));
    InMux I__4261 (
            .O(N__28858),
            .I(n12355));
    InMux I__4260 (
            .O(N__28855),
            .I(n12356));
    InMux I__4259 (
            .O(N__28852),
            .I(n12357));
    InMux I__4258 (
            .O(N__28849),
            .I(N__28846));
    LocalMux I__4257 (
            .O(N__28846),
            .I(n2581));
    InMux I__4256 (
            .O(N__28843),
            .I(n12358));
    InMux I__4255 (
            .O(N__28840),
            .I(n12359));
    InMux I__4254 (
            .O(N__28837),
            .I(n12360));
    InMux I__4253 (
            .O(N__28834),
            .I(n12343));
    InMux I__4252 (
            .O(N__28831),
            .I(n12344));
    InMux I__4251 (
            .O(N__28828),
            .I(n12345));
    InMux I__4250 (
            .O(N__28825),
            .I(bfn_6_15_0_));
    InMux I__4249 (
            .O(N__28822),
            .I(n12347));
    InMux I__4248 (
            .O(N__28819),
            .I(n12348));
    InMux I__4247 (
            .O(N__28816),
            .I(n12349));
    InMux I__4246 (
            .O(N__28813),
            .I(n12350));
    InMux I__4245 (
            .O(N__28810),
            .I(n12351));
    CascadeMux I__4244 (
            .O(N__28807),
            .I(N__28804));
    InMux I__4243 (
            .O(N__28804),
            .I(N__28801));
    LocalMux I__4242 (
            .O(N__28801),
            .I(N__28797));
    InMux I__4241 (
            .O(N__28800),
            .I(N__28794));
    Odrv12 I__4240 (
            .O(N__28797),
            .I(n1125));
    LocalMux I__4239 (
            .O(N__28794),
            .I(n1125));
    CascadeMux I__4238 (
            .O(N__28789),
            .I(N__28785));
    CascadeMux I__4237 (
            .O(N__28788),
            .I(N__28782));
    InMux I__4236 (
            .O(N__28785),
            .I(N__28779));
    InMux I__4235 (
            .O(N__28782),
            .I(N__28776));
    LocalMux I__4234 (
            .O(N__28779),
            .I(N__28771));
    LocalMux I__4233 (
            .O(N__28776),
            .I(N__28771));
    Odrv12 I__4232 (
            .O(N__28771),
            .I(n1126));
    CascadeMux I__4231 (
            .O(N__28768),
            .I(n1126_cascade_));
    CascadeMux I__4230 (
            .O(N__28765),
            .I(N__28762));
    InMux I__4229 (
            .O(N__28762),
            .I(N__28759));
    LocalMux I__4228 (
            .O(N__28759),
            .I(N__28755));
    InMux I__4227 (
            .O(N__28758),
            .I(N__28751));
    Span4Mux_h I__4226 (
            .O(N__28755),
            .I(N__28748));
    InMux I__4225 (
            .O(N__28754),
            .I(N__28745));
    LocalMux I__4224 (
            .O(N__28751),
            .I(n1127));
    Odrv4 I__4223 (
            .O(N__28748),
            .I(n1127));
    LocalMux I__4222 (
            .O(N__28745),
            .I(n1127));
    InMux I__4221 (
            .O(N__28738),
            .I(N__28735));
    LocalMux I__4220 (
            .O(N__28735),
            .I(n13994));
    InMux I__4219 (
            .O(N__28732),
            .I(bfn_6_14_0_));
    InMux I__4218 (
            .O(N__28729),
            .I(n12339));
    InMux I__4217 (
            .O(N__28726),
            .I(n12340));
    InMux I__4216 (
            .O(N__28723),
            .I(n12341));
    InMux I__4215 (
            .O(N__28720),
            .I(n12342));
    CascadeMux I__4214 (
            .O(N__28717),
            .I(n1228_cascade_));
    CascadeMux I__4213 (
            .O(N__28714),
            .I(N__28710));
    CascadeMux I__4212 (
            .O(N__28713),
            .I(N__28707));
    InMux I__4211 (
            .O(N__28710),
            .I(N__28703));
    InMux I__4210 (
            .O(N__28707),
            .I(N__28698));
    InMux I__4209 (
            .O(N__28706),
            .I(N__28698));
    LocalMux I__4208 (
            .O(N__28703),
            .I(n1226));
    LocalMux I__4207 (
            .O(N__28698),
            .I(n1226));
    InMux I__4206 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__4205 (
            .O(N__28690),
            .I(n14078));
    CascadeMux I__4204 (
            .O(N__28687),
            .I(N__28684));
    InMux I__4203 (
            .O(N__28684),
            .I(N__28679));
    InMux I__4202 (
            .O(N__28683),
            .I(N__28676));
    InMux I__4201 (
            .O(N__28682),
            .I(N__28673));
    LocalMux I__4200 (
            .O(N__28679),
            .I(N__28670));
    LocalMux I__4199 (
            .O(N__28676),
            .I(n1132));
    LocalMux I__4198 (
            .O(N__28673),
            .I(n1132));
    Odrv12 I__4197 (
            .O(N__28670),
            .I(n1132));
    CascadeMux I__4196 (
            .O(N__28663),
            .I(N__28660));
    InMux I__4195 (
            .O(N__28660),
            .I(N__28656));
    CascadeMux I__4194 (
            .O(N__28659),
            .I(N__28653));
    LocalMux I__4193 (
            .O(N__28656),
            .I(N__28650));
    InMux I__4192 (
            .O(N__28653),
            .I(N__28646));
    Span4Mux_s1_h I__4191 (
            .O(N__28650),
            .I(N__28643));
    InMux I__4190 (
            .O(N__28649),
            .I(N__28640));
    LocalMux I__4189 (
            .O(N__28646),
            .I(n1129));
    Odrv4 I__4188 (
            .O(N__28643),
            .I(n1129));
    LocalMux I__4187 (
            .O(N__28640),
            .I(n1129));
    CascadeMux I__4186 (
            .O(N__28633),
            .I(N__28630));
    InMux I__4185 (
            .O(N__28630),
            .I(N__28626));
    CascadeMux I__4184 (
            .O(N__28629),
            .I(N__28623));
    LocalMux I__4183 (
            .O(N__28626),
            .I(N__28619));
    InMux I__4182 (
            .O(N__28623),
            .I(N__28616));
    InMux I__4181 (
            .O(N__28622),
            .I(N__28613));
    Span4Mux_s1_h I__4180 (
            .O(N__28619),
            .I(N__28610));
    LocalMux I__4179 (
            .O(N__28616),
            .I(n1133));
    LocalMux I__4178 (
            .O(N__28613),
            .I(n1133));
    Odrv4 I__4177 (
            .O(N__28610),
            .I(n1133));
    InMux I__4176 (
            .O(N__28603),
            .I(N__28600));
    LocalMux I__4175 (
            .O(N__28600),
            .I(N__28597));
    Odrv12 I__4174 (
            .O(N__28597),
            .I(n1195));
    CascadeMux I__4173 (
            .O(N__28594),
            .I(N__28590));
    CascadeMux I__4172 (
            .O(N__28593),
            .I(N__28587));
    InMux I__4171 (
            .O(N__28590),
            .I(N__28584));
    InMux I__4170 (
            .O(N__28587),
            .I(N__28580));
    LocalMux I__4169 (
            .O(N__28584),
            .I(N__28577));
    InMux I__4168 (
            .O(N__28583),
            .I(N__28574));
    LocalMux I__4167 (
            .O(N__28580),
            .I(n1227));
    Odrv4 I__4166 (
            .O(N__28577),
            .I(n1227));
    LocalMux I__4165 (
            .O(N__28574),
            .I(n1227));
    InMux I__4164 (
            .O(N__28567),
            .I(N__28564));
    LocalMux I__4163 (
            .O(N__28564),
            .I(N__28561));
    Odrv12 I__4162 (
            .O(N__28561),
            .I(n1198));
    CascadeMux I__4161 (
            .O(N__28558),
            .I(N__28554));
    CascadeMux I__4160 (
            .O(N__28557),
            .I(N__28551));
    InMux I__4159 (
            .O(N__28554),
            .I(N__28548));
    InMux I__4158 (
            .O(N__28551),
            .I(N__28545));
    LocalMux I__4157 (
            .O(N__28548),
            .I(N__28542));
    LocalMux I__4156 (
            .O(N__28545),
            .I(n1230));
    Odrv4 I__4155 (
            .O(N__28542),
            .I(n1230));
    CascadeMux I__4154 (
            .O(N__28537),
            .I(N__28533));
    InMux I__4153 (
            .O(N__28536),
            .I(N__28529));
    InMux I__4152 (
            .O(N__28533),
            .I(N__28526));
    InMux I__4151 (
            .O(N__28532),
            .I(N__28523));
    LocalMux I__4150 (
            .O(N__28529),
            .I(n1229));
    LocalMux I__4149 (
            .O(N__28526),
            .I(n1229));
    LocalMux I__4148 (
            .O(N__28523),
            .I(n1229));
    CascadeMux I__4147 (
            .O(N__28516),
            .I(N__28512));
    CascadeMux I__4146 (
            .O(N__28515),
            .I(N__28508));
    InMux I__4145 (
            .O(N__28512),
            .I(N__28505));
    InMux I__4144 (
            .O(N__28511),
            .I(N__28502));
    InMux I__4143 (
            .O(N__28508),
            .I(N__28499));
    LocalMux I__4142 (
            .O(N__28505),
            .I(n1231));
    LocalMux I__4141 (
            .O(N__28502),
            .I(n1231));
    LocalMux I__4140 (
            .O(N__28499),
            .I(n1231));
    CascadeMux I__4139 (
            .O(N__28492),
            .I(n1230_cascade_));
    InMux I__4138 (
            .O(N__28489),
            .I(N__28486));
    LocalMux I__4137 (
            .O(N__28486),
            .I(n11642));
    InMux I__4136 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__4135 (
            .O(N__28480),
            .I(n13318));
    InMux I__4134 (
            .O(N__28477),
            .I(N__28474));
    LocalMux I__4133 (
            .O(N__28474),
            .I(N__28470));
    InMux I__4132 (
            .O(N__28473),
            .I(N__28467));
    Span4Mux_h I__4131 (
            .O(N__28470),
            .I(N__28464));
    LocalMux I__4130 (
            .O(N__28467),
            .I(N__28461));
    IoSpan4Mux I__4129 (
            .O(N__28464),
            .I(N__28458));
    Span4Mux_v I__4128 (
            .O(N__28461),
            .I(N__28455));
    Odrv4 I__4127 (
            .O(N__28458),
            .I(\debounce.reg_A_0 ));
    Odrv4 I__4126 (
            .O(N__28455),
            .I(\debounce.reg_A_0 ));
    CascadeMux I__4125 (
            .O(N__28450),
            .I(N__28447));
    InMux I__4124 (
            .O(N__28447),
            .I(N__28443));
    InMux I__4123 (
            .O(N__28446),
            .I(N__28440));
    LocalMux I__4122 (
            .O(N__28443),
            .I(N__28437));
    LocalMux I__4121 (
            .O(N__28440),
            .I(N__28434));
    Span4Mux_s3_v I__4120 (
            .O(N__28437),
            .I(N__28431));
    Odrv4 I__4119 (
            .O(N__28434),
            .I(reg_B_0));
    Odrv4 I__4118 (
            .O(N__28431),
            .I(reg_B_0));
    InMux I__4117 (
            .O(N__28426),
            .I(N__28423));
    LocalMux I__4116 (
            .O(N__28423),
            .I(n2288));
    InMux I__4115 (
            .O(N__28420),
            .I(N__28417));
    LocalMux I__4114 (
            .O(N__28417),
            .I(N__28414));
    Span4Mux_h I__4113 (
            .O(N__28414),
            .I(N__28411));
    Odrv4 I__4112 (
            .O(N__28411),
            .I(n1293));
    CascadeMux I__4111 (
            .O(N__28408),
            .I(N__28405));
    InMux I__4110 (
            .O(N__28405),
            .I(N__28401));
    InMux I__4109 (
            .O(N__28404),
            .I(N__28398));
    LocalMux I__4108 (
            .O(N__28401),
            .I(N__28395));
    LocalMux I__4107 (
            .O(N__28398),
            .I(n1325));
    Odrv4 I__4106 (
            .O(N__28395),
            .I(n1325));
    InMux I__4105 (
            .O(N__28390),
            .I(N__28386));
    CascadeMux I__4104 (
            .O(N__28389),
            .I(N__28383));
    LocalMux I__4103 (
            .O(N__28386),
            .I(N__28379));
    InMux I__4102 (
            .O(N__28383),
            .I(N__28376));
    InMux I__4101 (
            .O(N__28382),
            .I(N__28373));
    Odrv4 I__4100 (
            .O(N__28379),
            .I(n1326));
    LocalMux I__4099 (
            .O(N__28376),
            .I(n1326));
    LocalMux I__4098 (
            .O(N__28373),
            .I(n1326));
    CascadeMux I__4097 (
            .O(N__28366),
            .I(N__28363));
    InMux I__4096 (
            .O(N__28363),
            .I(N__28359));
    CascadeMux I__4095 (
            .O(N__28362),
            .I(N__28356));
    LocalMux I__4094 (
            .O(N__28359),
            .I(N__28352));
    InMux I__4093 (
            .O(N__28356),
            .I(N__28349));
    InMux I__4092 (
            .O(N__28355),
            .I(N__28346));
    Odrv4 I__4091 (
            .O(N__28352),
            .I(n1327));
    LocalMux I__4090 (
            .O(N__28349),
            .I(n1327));
    LocalMux I__4089 (
            .O(N__28346),
            .I(n1327));
    CascadeMux I__4088 (
            .O(N__28339),
            .I(n1325_cascade_));
    CascadeMux I__4087 (
            .O(N__28336),
            .I(N__28333));
    InMux I__4086 (
            .O(N__28333),
            .I(N__28330));
    LocalMux I__4085 (
            .O(N__28330),
            .I(N__28326));
    CascadeMux I__4084 (
            .O(N__28329),
            .I(N__28323));
    Span4Mux_s3_h I__4083 (
            .O(N__28326),
            .I(N__28319));
    InMux I__4082 (
            .O(N__28323),
            .I(N__28316));
    InMux I__4081 (
            .O(N__28322),
            .I(N__28313));
    Odrv4 I__4080 (
            .O(N__28319),
            .I(n1328));
    LocalMux I__4079 (
            .O(N__28316),
            .I(n1328));
    LocalMux I__4078 (
            .O(N__28313),
            .I(n1328));
    InMux I__4077 (
            .O(N__28306),
            .I(N__28303));
    LocalMux I__4076 (
            .O(N__28303),
            .I(n13734));
    InMux I__4075 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__4074 (
            .O(N__28297),
            .I(N__28293));
    InMux I__4073 (
            .O(N__28296),
            .I(N__28290));
    Span4Mux_s2_v I__4072 (
            .O(N__28293),
            .I(N__28287));
    LocalMux I__4071 (
            .O(N__28290),
            .I(n298));
    Odrv4 I__4070 (
            .O(N__28287),
            .I(n298));
    CascadeMux I__4069 (
            .O(N__28282),
            .I(N__28279));
    InMux I__4068 (
            .O(N__28279),
            .I(N__28275));
    InMux I__4067 (
            .O(N__28278),
            .I(N__28272));
    LocalMux I__4066 (
            .O(N__28275),
            .I(n1233));
    LocalMux I__4065 (
            .O(N__28272),
            .I(n1233));
    CascadeMux I__4064 (
            .O(N__28267),
            .I(n298_cascade_));
    CascadeMux I__4063 (
            .O(N__28264),
            .I(N__28260));
    InMux I__4062 (
            .O(N__28263),
            .I(N__28256));
    InMux I__4061 (
            .O(N__28260),
            .I(N__28253));
    InMux I__4060 (
            .O(N__28259),
            .I(N__28250));
    LocalMux I__4059 (
            .O(N__28256),
            .I(n1232));
    LocalMux I__4058 (
            .O(N__28253),
            .I(n1232));
    LocalMux I__4057 (
            .O(N__28250),
            .I(n1232));
    InMux I__4056 (
            .O(N__28243),
            .I(N__28240));
    LocalMux I__4055 (
            .O(N__28240),
            .I(N__28237));
    Span4Mux_h I__4054 (
            .O(N__28237),
            .I(N__28234));
    Odrv4 I__4053 (
            .O(N__28234),
            .I(n1196));
    CascadeMux I__4052 (
            .O(N__28231),
            .I(N__28228));
    InMux I__4051 (
            .O(N__28228),
            .I(N__28224));
    InMux I__4050 (
            .O(N__28227),
            .I(N__28221));
    LocalMux I__4049 (
            .O(N__28224),
            .I(N__28218));
    LocalMux I__4048 (
            .O(N__28221),
            .I(N__28213));
    Span4Mux_s2_v I__4047 (
            .O(N__28218),
            .I(N__28213));
    Odrv4 I__4046 (
            .O(N__28213),
            .I(n1228));
    InMux I__4045 (
            .O(N__28210),
            .I(N__28207));
    LocalMux I__4044 (
            .O(N__28207),
            .I(n2287));
    InMux I__4043 (
            .O(N__28204),
            .I(n12098));
    InMux I__4042 (
            .O(N__28201),
            .I(n12099));
    CascadeMux I__4041 (
            .O(N__28198),
            .I(N__28195));
    InMux I__4040 (
            .O(N__28195),
            .I(N__28192));
    LocalMux I__4039 (
            .O(N__28192),
            .I(n402));
    InMux I__4038 (
            .O(N__28189),
            .I(n12100));
    InMux I__4037 (
            .O(N__28186),
            .I(N__28183));
    LocalMux I__4036 (
            .O(N__28183),
            .I(n2289));
    CascadeMux I__4035 (
            .O(N__28180),
            .I(n13261_cascade_));
    InMux I__4034 (
            .O(N__28177),
            .I(N__28173));
    InMux I__4033 (
            .O(N__28176),
            .I(N__28170));
    LocalMux I__4032 (
            .O(N__28173),
            .I(N__28166));
    LocalMux I__4031 (
            .O(N__28170),
            .I(N__28163));
    InMux I__4030 (
            .O(N__28169),
            .I(N__28160));
    Span4Mux_s2_v I__4029 (
            .O(N__28166),
            .I(N__28157));
    Span4Mux_h I__4028 (
            .O(N__28163),
            .I(N__28154));
    LocalMux I__4027 (
            .O(N__28160),
            .I(n297));
    Odrv4 I__4026 (
            .O(N__28157),
            .I(n297));
    Odrv4 I__4025 (
            .O(N__28154),
            .I(n297));
    InMux I__4024 (
            .O(N__28147),
            .I(N__28144));
    LocalMux I__4023 (
            .O(N__28144),
            .I(N__28140));
    InMux I__4022 (
            .O(N__28143),
            .I(N__28137));
    Span4Mux_v I__4021 (
            .O(N__28140),
            .I(N__28134));
    LocalMux I__4020 (
            .O(N__28137),
            .I(N__28131));
    Span4Mux_h I__4019 (
            .O(N__28134),
            .I(N__28128));
    IoSpan4Mux I__4018 (
            .O(N__28131),
            .I(N__28125));
    Odrv4 I__4017 (
            .O(N__28128),
            .I(\debounce.reg_A_1 ));
    Odrv4 I__4016 (
            .O(N__28125),
            .I(\debounce.reg_A_1 ));
    InMux I__4015 (
            .O(N__28120),
            .I(N__28116));
    InMux I__4014 (
            .O(N__28119),
            .I(N__28113));
    LocalMux I__4013 (
            .O(N__28116),
            .I(N__28108));
    LocalMux I__4012 (
            .O(N__28113),
            .I(N__28108));
    Span4Mux_s3_v I__4011 (
            .O(N__28108),
            .I(N__28105));
    Odrv4 I__4010 (
            .O(N__28105),
            .I(reg_B_1));
    CascadeMux I__4009 (
            .O(N__28102),
            .I(n13257_cascade_));
    InMux I__4008 (
            .O(N__28099),
            .I(N__28094));
    InMux I__4007 (
            .O(N__28098),
            .I(N__28091));
    InMux I__4006 (
            .O(N__28097),
            .I(N__28088));
    LocalMux I__4005 (
            .O(N__28094),
            .I(N__28085));
    LocalMux I__4004 (
            .O(N__28091),
            .I(N__28080));
    LocalMux I__4003 (
            .O(N__28088),
            .I(N__28080));
    Span4Mux_v I__4002 (
            .O(N__28085),
            .I(N__28077));
    Span4Mux_h I__4001 (
            .O(N__28080),
            .I(N__28074));
    Odrv4 I__4000 (
            .O(N__28077),
            .I(n302));
    Odrv4 I__3999 (
            .O(N__28074),
            .I(n302));
    InMux I__3998 (
            .O(N__28069),
            .I(bfn_5_28_0_));
    InMux I__3997 (
            .O(N__28066),
            .I(n12096));
    InMux I__3996 (
            .O(N__28063),
            .I(n12097));
    InMux I__3995 (
            .O(N__28060),
            .I(N__28057));
    LocalMux I__3994 (
            .O(N__28057),
            .I(N__28054));
    Span4Mux_v I__3993 (
            .O(N__28054),
            .I(N__28051));
    Odrv4 I__3992 (
            .O(N__28051),
            .I(n1801));
    InMux I__3991 (
            .O(N__28048),
            .I(N__28045));
    LocalMux I__3990 (
            .O(N__28045),
            .I(N__28040));
    InMux I__3989 (
            .O(N__28044),
            .I(N__28037));
    InMux I__3988 (
            .O(N__28043),
            .I(N__28034));
    Span4Mux_v I__3987 (
            .O(N__28040),
            .I(N__28031));
    LocalMux I__3986 (
            .O(N__28037),
            .I(n303));
    LocalMux I__3985 (
            .O(N__28034),
            .I(n303));
    Odrv4 I__3984 (
            .O(N__28031),
            .I(n303));
    CascadeMux I__3983 (
            .O(N__28024),
            .I(N__28021));
    InMux I__3982 (
            .O(N__28021),
            .I(N__28016));
    InMux I__3981 (
            .O(N__28020),
            .I(N__28013));
    InMux I__3980 (
            .O(N__28019),
            .I(N__28010));
    LocalMux I__3979 (
            .O(N__28016),
            .I(N__28007));
    LocalMux I__3978 (
            .O(N__28013),
            .I(N__28004));
    LocalMux I__3977 (
            .O(N__28010),
            .I(N__27999));
    Span4Mux_h I__3976 (
            .O(N__28007),
            .I(N__27999));
    Odrv4 I__3975 (
            .O(N__28004),
            .I(n1833));
    Odrv4 I__3974 (
            .O(N__27999),
            .I(n1833));
    InMux I__3973 (
            .O(N__27994),
            .I(N__27990));
    InMux I__3972 (
            .O(N__27993),
            .I(N__27987));
    LocalMux I__3971 (
            .O(N__27990),
            .I(N__27984));
    LocalMux I__3970 (
            .O(N__27987),
            .I(N__27981));
    Span4Mux_v I__3969 (
            .O(N__27984),
            .I(N__27978));
    Span4Mux_v I__3968 (
            .O(N__27981),
            .I(N__27974));
    Span4Mux_v I__3967 (
            .O(N__27978),
            .I(N__27971));
    InMux I__3966 (
            .O(N__27977),
            .I(N__27968));
    Span4Mux_v I__3965 (
            .O(N__27974),
            .I(N__27965));
    Span4Mux_h I__3964 (
            .O(N__27971),
            .I(N__27962));
    LocalMux I__3963 (
            .O(N__27968),
            .I(N__27959));
    Odrv4 I__3962 (
            .O(N__27965),
            .I(n307));
    Odrv4 I__3961 (
            .O(N__27962),
            .I(n307));
    Odrv12 I__3960 (
            .O(N__27959),
            .I(n307));
    InMux I__3959 (
            .O(N__27952),
            .I(N__27949));
    LocalMux I__3958 (
            .O(N__27949),
            .I(N__27946));
    Span4Mux_v I__3957 (
            .O(N__27946),
            .I(N__27940));
    InMux I__3956 (
            .O(N__27945),
            .I(N__27937));
    InMux I__3955 (
            .O(N__27944),
            .I(N__27932));
    InMux I__3954 (
            .O(N__27943),
            .I(N__27932));
    Span4Mux_v I__3953 (
            .O(N__27940),
            .I(N__27925));
    LocalMux I__3952 (
            .O(N__27937),
            .I(N__27925));
    LocalMux I__3951 (
            .O(N__27932),
            .I(N__27925));
    Odrv4 I__3950 (
            .O(N__27925),
            .I(n13490));
    InMux I__3949 (
            .O(N__27922),
            .I(N__27918));
    InMux I__3948 (
            .O(N__27921),
            .I(N__27915));
    LocalMux I__3947 (
            .O(N__27918),
            .I(N__27911));
    LocalMux I__3946 (
            .O(N__27915),
            .I(N__27908));
    InMux I__3945 (
            .O(N__27914),
            .I(N__27905));
    Span4Mux_v I__3944 (
            .O(N__27911),
            .I(N__27902));
    Span4Mux_h I__3943 (
            .O(N__27908),
            .I(N__27897));
    LocalMux I__3942 (
            .O(N__27905),
            .I(N__27897));
    Span4Mux_v I__3941 (
            .O(N__27902),
            .I(N__27894));
    Span4Mux_v I__3940 (
            .O(N__27897),
            .I(N__27891));
    Odrv4 I__3939 (
            .O(N__27894),
            .I(n306));
    Odrv4 I__3938 (
            .O(N__27891),
            .I(n306));
    InMux I__3937 (
            .O(N__27886),
            .I(N__27882));
    CascadeMux I__3936 (
            .O(N__27885),
            .I(N__27879));
    LocalMux I__3935 (
            .O(N__27882),
            .I(N__27876));
    InMux I__3934 (
            .O(N__27879),
            .I(N__27873));
    Span4Mux_v I__3933 (
            .O(N__27876),
            .I(N__27867));
    LocalMux I__3932 (
            .O(N__27873),
            .I(N__27867));
    InMux I__3931 (
            .O(N__27872),
            .I(N__27864));
    Odrv4 I__3930 (
            .O(N__27867),
            .I(n1726));
    LocalMux I__3929 (
            .O(N__27864),
            .I(n1726));
    InMux I__3928 (
            .O(N__27859),
            .I(N__27855));
    CascadeMux I__3927 (
            .O(N__27858),
            .I(N__27852));
    LocalMux I__3926 (
            .O(N__27855),
            .I(N__27849));
    InMux I__3925 (
            .O(N__27852),
            .I(N__27846));
    Span4Mux_v I__3924 (
            .O(N__27849),
            .I(N__27843));
    LocalMux I__3923 (
            .O(N__27846),
            .I(N__27840));
    Odrv4 I__3922 (
            .O(N__27843),
            .I(n1825));
    Odrv12 I__3921 (
            .O(N__27840),
            .I(n1825));
    CascadeMux I__3920 (
            .O(N__27835),
            .I(N__27831));
    CascadeMux I__3919 (
            .O(N__27834),
            .I(N__27828));
    InMux I__3918 (
            .O(N__27831),
            .I(N__27825));
    InMux I__3917 (
            .O(N__27828),
            .I(N__27822));
    LocalMux I__3916 (
            .O(N__27825),
            .I(N__27816));
    LocalMux I__3915 (
            .O(N__27822),
            .I(N__27816));
    InMux I__3914 (
            .O(N__27821),
            .I(N__27813));
    Odrv4 I__3913 (
            .O(N__27816),
            .I(n1827));
    LocalMux I__3912 (
            .O(N__27813),
            .I(n1827));
    CascadeMux I__3911 (
            .O(N__27808),
            .I(N__27805));
    InMux I__3910 (
            .O(N__27805),
            .I(N__27802));
    LocalMux I__3909 (
            .O(N__27802),
            .I(N__27798));
    InMux I__3908 (
            .O(N__27801),
            .I(N__27794));
    Span4Mux_s3_h I__3907 (
            .O(N__27798),
            .I(N__27791));
    InMux I__3906 (
            .O(N__27797),
            .I(N__27788));
    LocalMux I__3905 (
            .O(N__27794),
            .I(n1826));
    Odrv4 I__3904 (
            .O(N__27791),
            .I(n1826));
    LocalMux I__3903 (
            .O(N__27788),
            .I(n1826));
    CascadeMux I__3902 (
            .O(N__27781),
            .I(n1825_cascade_));
    InMux I__3901 (
            .O(N__27778),
            .I(N__27775));
    LocalMux I__3900 (
            .O(N__27775),
            .I(n14122));
    InMux I__3899 (
            .O(N__27772),
            .I(N__27768));
    CascadeMux I__3898 (
            .O(N__27771),
            .I(N__27765));
    LocalMux I__3897 (
            .O(N__27768),
            .I(N__27762));
    InMux I__3896 (
            .O(N__27765),
            .I(N__27759));
    Span4Mux_h I__3895 (
            .O(N__27762),
            .I(N__27754));
    LocalMux I__3894 (
            .O(N__27759),
            .I(N__27754));
    Odrv4 I__3893 (
            .O(N__27754),
            .I(n1729));
    CascadeMux I__3892 (
            .O(N__27751),
            .I(N__27748));
    InMux I__3891 (
            .O(N__27748),
            .I(N__27745));
    LocalMux I__3890 (
            .O(N__27745),
            .I(n1796));
    CascadeMux I__3889 (
            .O(N__27742),
            .I(N__27738));
    InMux I__3888 (
            .O(N__27741),
            .I(N__27735));
    InMux I__3887 (
            .O(N__27738),
            .I(N__27732));
    LocalMux I__3886 (
            .O(N__27735),
            .I(N__27729));
    LocalMux I__3885 (
            .O(N__27732),
            .I(N__27726));
    Span4Mux_v I__3884 (
            .O(N__27729),
            .I(N__27720));
    Span4Mux_h I__3883 (
            .O(N__27726),
            .I(N__27720));
    InMux I__3882 (
            .O(N__27725),
            .I(N__27717));
    Odrv4 I__3881 (
            .O(N__27720),
            .I(n1828));
    LocalMux I__3880 (
            .O(N__27717),
            .I(n1828));
    CascadeMux I__3879 (
            .O(N__27712),
            .I(N__27707));
    CascadeMux I__3878 (
            .O(N__27711),
            .I(N__27704));
    InMux I__3877 (
            .O(N__27710),
            .I(N__27701));
    InMux I__3876 (
            .O(N__27707),
            .I(N__27698));
    InMux I__3875 (
            .O(N__27704),
            .I(N__27695));
    LocalMux I__3874 (
            .O(N__27701),
            .I(N__27692));
    LocalMux I__3873 (
            .O(N__27698),
            .I(n1832));
    LocalMux I__3872 (
            .O(N__27695),
            .I(n1832));
    Odrv12 I__3871 (
            .O(N__27692),
            .I(n1832));
    CascadeMux I__3870 (
            .O(N__27685),
            .I(N__27682));
    InMux I__3869 (
            .O(N__27682),
            .I(N__27677));
    CascadeMux I__3868 (
            .O(N__27681),
            .I(N__27674));
    InMux I__3867 (
            .O(N__27680),
            .I(N__27671));
    LocalMux I__3866 (
            .O(N__27677),
            .I(N__27668));
    InMux I__3865 (
            .O(N__27674),
            .I(N__27665));
    LocalMux I__3864 (
            .O(N__27671),
            .I(n1831));
    Odrv4 I__3863 (
            .O(N__27668),
            .I(n1831));
    LocalMux I__3862 (
            .O(N__27665),
            .I(n1831));
    InMux I__3861 (
            .O(N__27658),
            .I(N__27655));
    LocalMux I__3860 (
            .O(N__27655),
            .I(n11688));
    CascadeMux I__3859 (
            .O(N__27652),
            .I(N__27648));
    InMux I__3858 (
            .O(N__27651),
            .I(N__27645));
    InMux I__3857 (
            .O(N__27648),
            .I(N__27642));
    LocalMux I__3856 (
            .O(N__27645),
            .I(N__27639));
    LocalMux I__3855 (
            .O(N__27642),
            .I(N__27636));
    Span4Mux_v I__3854 (
            .O(N__27639),
            .I(N__27630));
    Span4Mux_s1_h I__3853 (
            .O(N__27636),
            .I(N__27630));
    InMux I__3852 (
            .O(N__27635),
            .I(N__27627));
    Odrv4 I__3851 (
            .O(N__27630),
            .I(n2021));
    LocalMux I__3850 (
            .O(N__27627),
            .I(n2021));
    CascadeMux I__3849 (
            .O(N__27622),
            .I(N__27619));
    InMux I__3848 (
            .O(N__27619),
            .I(N__27616));
    LocalMux I__3847 (
            .O(N__27616),
            .I(N__27613));
    Span4Mux_v I__3846 (
            .O(N__27613),
            .I(N__27610));
    Odrv4 I__3845 (
            .O(N__27610),
            .I(n2088));
    InMux I__3844 (
            .O(N__27607),
            .I(N__27603));
    InMux I__3843 (
            .O(N__27606),
            .I(N__27600));
    LocalMux I__3842 (
            .O(N__27603),
            .I(N__27597));
    LocalMux I__3841 (
            .O(N__27600),
            .I(N__27593));
    Span4Mux_v I__3840 (
            .O(N__27597),
            .I(N__27590));
    InMux I__3839 (
            .O(N__27596),
            .I(N__27587));
    Span4Mux_v I__3838 (
            .O(N__27593),
            .I(N__27582));
    Span4Mux_h I__3837 (
            .O(N__27590),
            .I(N__27582));
    LocalMux I__3836 (
            .O(N__27587),
            .I(N__27579));
    Odrv4 I__3835 (
            .O(N__27582),
            .I(n2120));
    Odrv4 I__3834 (
            .O(N__27579),
            .I(n2120));
    CascadeMux I__3833 (
            .O(N__27574),
            .I(N__27571));
    InMux I__3832 (
            .O(N__27571),
            .I(N__27567));
    InMux I__3831 (
            .O(N__27570),
            .I(N__27564));
    LocalMux I__3830 (
            .O(N__27567),
            .I(N__27558));
    LocalMux I__3829 (
            .O(N__27564),
            .I(N__27558));
    InMux I__3828 (
            .O(N__27563),
            .I(N__27555));
    Span4Mux_h I__3827 (
            .O(N__27558),
            .I(N__27552));
    LocalMux I__3826 (
            .O(N__27555),
            .I(n301));
    Odrv4 I__3825 (
            .O(N__27552),
            .I(n301));
    InMux I__3824 (
            .O(N__27547),
            .I(N__27544));
    LocalMux I__3823 (
            .O(N__27544),
            .I(N__27541));
    Odrv12 I__3822 (
            .O(N__27541),
            .I(n1897));
    CascadeMux I__3821 (
            .O(N__27538),
            .I(N__27534));
    InMux I__3820 (
            .O(N__27537),
            .I(N__27531));
    InMux I__3819 (
            .O(N__27534),
            .I(N__27528));
    LocalMux I__3818 (
            .O(N__27531),
            .I(N__27525));
    LocalMux I__3817 (
            .O(N__27528),
            .I(N__27522));
    Span4Mux_v I__3816 (
            .O(N__27525),
            .I(N__27519));
    Span4Mux_v I__3815 (
            .O(N__27522),
            .I(N__27516));
    Odrv4 I__3814 (
            .O(N__27519),
            .I(n1929));
    Odrv4 I__3813 (
            .O(N__27516),
            .I(n1929));
    CascadeMux I__3812 (
            .O(N__27511),
            .I(n1929_cascade_));
    InMux I__3811 (
            .O(N__27508),
            .I(N__27505));
    LocalMux I__3810 (
            .O(N__27505),
            .I(n14136));
    InMux I__3809 (
            .O(N__27502),
            .I(N__27499));
    LocalMux I__3808 (
            .O(N__27499),
            .I(N__27496));
    Odrv12 I__3807 (
            .O(N__27496),
            .I(n1901));
    CascadeMux I__3806 (
            .O(N__27493),
            .I(N__27490));
    InMux I__3805 (
            .O(N__27490),
            .I(N__27486));
    CascadeMux I__3804 (
            .O(N__27489),
            .I(N__27483));
    LocalMux I__3803 (
            .O(N__27486),
            .I(N__27479));
    InMux I__3802 (
            .O(N__27483),
            .I(N__27476));
    InMux I__3801 (
            .O(N__27482),
            .I(N__27473));
    Span4Mux_h I__3800 (
            .O(N__27479),
            .I(N__27470));
    LocalMux I__3799 (
            .O(N__27476),
            .I(n1933));
    LocalMux I__3798 (
            .O(N__27473),
            .I(n1933));
    Odrv4 I__3797 (
            .O(N__27470),
            .I(n1933));
    InMux I__3796 (
            .O(N__27463),
            .I(N__27460));
    LocalMux I__3795 (
            .O(N__27460),
            .I(N__27457));
    Odrv12 I__3794 (
            .O(N__27457),
            .I(n1898));
    CascadeMux I__3793 (
            .O(N__27454),
            .I(N__27450));
    InMux I__3792 (
            .O(N__27453),
            .I(N__27447));
    InMux I__3791 (
            .O(N__27450),
            .I(N__27444));
    LocalMux I__3790 (
            .O(N__27447),
            .I(N__27439));
    LocalMux I__3789 (
            .O(N__27444),
            .I(N__27439));
    Span4Mux_h I__3788 (
            .O(N__27439),
            .I(N__27435));
    InMux I__3787 (
            .O(N__27438),
            .I(N__27432));
    Odrv4 I__3786 (
            .O(N__27435),
            .I(n1930));
    LocalMux I__3785 (
            .O(N__27432),
            .I(n1930));
    InMux I__3784 (
            .O(N__27427),
            .I(N__27424));
    LocalMux I__3783 (
            .O(N__27424),
            .I(N__27421));
    Span4Mux_h I__3782 (
            .O(N__27421),
            .I(N__27418));
    Odrv4 I__3781 (
            .O(N__27418),
            .I(n1885));
    CascadeMux I__3780 (
            .O(N__27415),
            .I(N__27410));
    CascadeMux I__3779 (
            .O(N__27414),
            .I(N__27407));
    InMux I__3778 (
            .O(N__27413),
            .I(N__27404));
    InMux I__3777 (
            .O(N__27410),
            .I(N__27401));
    InMux I__3776 (
            .O(N__27407),
            .I(N__27398));
    LocalMux I__3775 (
            .O(N__27404),
            .I(N__27395));
    LocalMux I__3774 (
            .O(N__27401),
            .I(N__27392));
    LocalMux I__3773 (
            .O(N__27398),
            .I(N__27389));
    Span4Mux_h I__3772 (
            .O(N__27395),
            .I(N__27386));
    Odrv4 I__3771 (
            .O(N__27392),
            .I(n1818));
    Odrv4 I__3770 (
            .O(N__27389),
            .I(n1818));
    Odrv4 I__3769 (
            .O(N__27386),
            .I(n1818));
    CascadeMux I__3768 (
            .O(N__27379),
            .I(N__27376));
    InMux I__3767 (
            .O(N__27376),
            .I(N__27373));
    LocalMux I__3766 (
            .O(N__27373),
            .I(N__27369));
    InMux I__3765 (
            .O(N__27372),
            .I(N__27366));
    Odrv4 I__3764 (
            .O(N__27369),
            .I(n1917));
    LocalMux I__3763 (
            .O(N__27366),
            .I(n1917));
    InMux I__3762 (
            .O(N__27361),
            .I(N__27358));
    LocalMux I__3761 (
            .O(N__27358),
            .I(n1791));
    CascadeMux I__3760 (
            .O(N__27355),
            .I(N__27352));
    InMux I__3759 (
            .O(N__27352),
            .I(N__27349));
    LocalMux I__3758 (
            .O(N__27349),
            .I(N__27345));
    CascadeMux I__3757 (
            .O(N__27348),
            .I(N__27342));
    Span4Mux_h I__3756 (
            .O(N__27345),
            .I(N__27338));
    InMux I__3755 (
            .O(N__27342),
            .I(N__27335));
    InMux I__3754 (
            .O(N__27341),
            .I(N__27332));
    Odrv4 I__3753 (
            .O(N__27338),
            .I(n1724));
    LocalMux I__3752 (
            .O(N__27335),
            .I(n1724));
    LocalMux I__3751 (
            .O(N__27332),
            .I(n1724));
    InMux I__3750 (
            .O(N__27325),
            .I(N__27321));
    InMux I__3749 (
            .O(N__27324),
            .I(N__27318));
    LocalMux I__3748 (
            .O(N__27321),
            .I(N__27315));
    LocalMux I__3747 (
            .O(N__27318),
            .I(n1823));
    Odrv12 I__3746 (
            .O(N__27315),
            .I(n1823));
    CascadeMux I__3745 (
            .O(N__27310),
            .I(N__27307));
    InMux I__3744 (
            .O(N__27307),
            .I(N__27303));
    InMux I__3743 (
            .O(N__27306),
            .I(N__27299));
    LocalMux I__3742 (
            .O(N__27303),
            .I(N__27296));
    InMux I__3741 (
            .O(N__27302),
            .I(N__27293));
    LocalMux I__3740 (
            .O(N__27299),
            .I(N__27290));
    Span4Mux_s1_h I__3739 (
            .O(N__27296),
            .I(N__27285));
    LocalMux I__3738 (
            .O(N__27293),
            .I(N__27285));
    Odrv4 I__3737 (
            .O(N__27290),
            .I(n1824));
    Odrv4 I__3736 (
            .O(N__27285),
            .I(n1824));
    CascadeMux I__3735 (
            .O(N__27280),
            .I(n1823_cascade_));
    CascadeMux I__3734 (
            .O(N__27277),
            .I(N__27273));
    InMux I__3733 (
            .O(N__27276),
            .I(N__27269));
    InMux I__3732 (
            .O(N__27273),
            .I(N__27266));
    CascadeMux I__3731 (
            .O(N__27272),
            .I(N__27263));
    LocalMux I__3730 (
            .O(N__27269),
            .I(N__27260));
    LocalMux I__3729 (
            .O(N__27266),
            .I(N__27257));
    InMux I__3728 (
            .O(N__27263),
            .I(N__27254));
    Span4Mux_h I__3727 (
            .O(N__27260),
            .I(N__27251));
    Odrv4 I__3726 (
            .O(N__27257),
            .I(n1830));
    LocalMux I__3725 (
            .O(N__27254),
            .I(n1830));
    Odrv4 I__3724 (
            .O(N__27251),
            .I(n1830));
    CascadeMux I__3723 (
            .O(N__27244),
            .I(N__27241));
    InMux I__3722 (
            .O(N__27241),
            .I(N__27237));
    InMux I__3721 (
            .O(N__27240),
            .I(N__27233));
    LocalMux I__3720 (
            .O(N__27237),
            .I(N__27230));
    InMux I__3719 (
            .O(N__27236),
            .I(N__27227));
    LocalMux I__3718 (
            .O(N__27233),
            .I(N__27224));
    Span4Mux_s1_h I__3717 (
            .O(N__27230),
            .I(N__27221));
    LocalMux I__3716 (
            .O(N__27227),
            .I(n1829));
    Odrv4 I__3715 (
            .O(N__27224),
            .I(n1829));
    Odrv4 I__3714 (
            .O(N__27221),
            .I(n1829));
    CascadeMux I__3713 (
            .O(N__27214),
            .I(n14126_cascade_));
    CascadeMux I__3712 (
            .O(N__27211),
            .I(N__27208));
    InMux I__3711 (
            .O(N__27208),
            .I(N__27205));
    LocalMux I__3710 (
            .O(N__27205),
            .I(N__27202));
    Odrv4 I__3709 (
            .O(N__27202),
            .I(n14128));
    InMux I__3708 (
            .O(N__27199),
            .I(N__27196));
    LocalMux I__3707 (
            .O(N__27196),
            .I(n1793));
    InMux I__3706 (
            .O(N__27193),
            .I(N__27190));
    LocalMux I__3705 (
            .O(N__27190),
            .I(N__27187));
    Span4Mux_h I__3704 (
            .O(N__27187),
            .I(N__27184));
    Odrv4 I__3703 (
            .O(N__27184),
            .I(n2000));
    CascadeMux I__3702 (
            .O(N__27181),
            .I(N__27177));
    CascadeMux I__3701 (
            .O(N__27180),
            .I(N__27174));
    InMux I__3700 (
            .O(N__27177),
            .I(N__27171));
    InMux I__3699 (
            .O(N__27174),
            .I(N__27168));
    LocalMux I__3698 (
            .O(N__27171),
            .I(N__27165));
    LocalMux I__3697 (
            .O(N__27168),
            .I(N__27159));
    Span4Mux_h I__3696 (
            .O(N__27165),
            .I(N__27159));
    InMux I__3695 (
            .O(N__27164),
            .I(N__27156));
    Odrv4 I__3694 (
            .O(N__27159),
            .I(n2032));
    LocalMux I__3693 (
            .O(N__27156),
            .I(n2032));
    InMux I__3692 (
            .O(N__27151),
            .I(N__27148));
    LocalMux I__3691 (
            .O(N__27148),
            .I(N__27145));
    Span4Mux_h I__3690 (
            .O(N__27145),
            .I(N__27142));
    Odrv4 I__3689 (
            .O(N__27142),
            .I(n2091));
    CascadeMux I__3688 (
            .O(N__27139),
            .I(N__27136));
    InMux I__3687 (
            .O(N__27136),
            .I(N__27133));
    LocalMux I__3686 (
            .O(N__27133),
            .I(N__27129));
    InMux I__3685 (
            .O(N__27132),
            .I(N__27125));
    Span4Mux_s3_h I__3684 (
            .O(N__27129),
            .I(N__27122));
    InMux I__3683 (
            .O(N__27128),
            .I(N__27119));
    LocalMux I__3682 (
            .O(N__27125),
            .I(n2024));
    Odrv4 I__3681 (
            .O(N__27122),
            .I(n2024));
    LocalMux I__3680 (
            .O(N__27119),
            .I(n2024));
    CascadeMux I__3679 (
            .O(N__27112),
            .I(N__27109));
    InMux I__3678 (
            .O(N__27109),
            .I(N__27106));
    LocalMux I__3677 (
            .O(N__27106),
            .I(N__27102));
    InMux I__3676 (
            .O(N__27105),
            .I(N__27099));
    Span4Mux_h I__3675 (
            .O(N__27102),
            .I(N__27096));
    LocalMux I__3674 (
            .O(N__27099),
            .I(n2123));
    Odrv4 I__3673 (
            .O(N__27096),
            .I(n2123));
    CascadeMux I__3672 (
            .O(N__27091),
            .I(n2123_cascade_));
    InMux I__3671 (
            .O(N__27088),
            .I(N__27084));
    CascadeMux I__3670 (
            .O(N__27087),
            .I(N__27081));
    LocalMux I__3669 (
            .O(N__27084),
            .I(N__27078));
    InMux I__3668 (
            .O(N__27081),
            .I(N__27075));
    Span4Mux_v I__3667 (
            .O(N__27078),
            .I(N__27072));
    LocalMux I__3666 (
            .O(N__27075),
            .I(n2121));
    Odrv4 I__3665 (
            .O(N__27072),
            .I(n2121));
    CascadeMux I__3664 (
            .O(N__27067),
            .I(n13746_cascade_));
    InMux I__3663 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__3662 (
            .O(N__27061),
            .I(n13748));
    InMux I__3661 (
            .O(N__27058),
            .I(N__27054));
    InMux I__3660 (
            .O(N__27057),
            .I(N__27050));
    LocalMux I__3659 (
            .O(N__27054),
            .I(N__27047));
    InMux I__3658 (
            .O(N__27053),
            .I(N__27044));
    LocalMux I__3657 (
            .O(N__27050),
            .I(N__27041));
    Span4Mux_h I__3656 (
            .O(N__27047),
            .I(N__27038));
    LocalMux I__3655 (
            .O(N__27044),
            .I(n2119));
    Odrv4 I__3654 (
            .O(N__27041),
            .I(n2119));
    Odrv4 I__3653 (
            .O(N__27038),
            .I(n2119));
    CascadeMux I__3652 (
            .O(N__27031),
            .I(n13754_cascade_));
    InMux I__3651 (
            .O(N__27028),
            .I(N__27025));
    LocalMux I__3650 (
            .O(N__27025),
            .I(n13382));
    InMux I__3649 (
            .O(N__27022),
            .I(N__27019));
    LocalMux I__3648 (
            .O(N__27019),
            .I(N__27016));
    Span4Mux_h I__3647 (
            .O(N__27016),
            .I(N__27013));
    Odrv4 I__3646 (
            .O(N__27013),
            .I(n13760));
    CascadeMux I__3645 (
            .O(N__27010),
            .I(N__27007));
    InMux I__3644 (
            .O(N__27007),
            .I(N__27003));
    InMux I__3643 (
            .O(N__27006),
            .I(N__27000));
    LocalMux I__3642 (
            .O(N__27003),
            .I(N__26997));
    LocalMux I__3641 (
            .O(N__27000),
            .I(N__26994));
    Span4Mux_s2_h I__3640 (
            .O(N__26997),
            .I(N__26991));
    Odrv4 I__3639 (
            .O(N__26994),
            .I(n1822));
    Odrv4 I__3638 (
            .O(N__26991),
            .I(n1822));
    InMux I__3637 (
            .O(N__26986),
            .I(N__26983));
    LocalMux I__3636 (
            .O(N__26983),
            .I(N__26980));
    Span4Mux_h I__3635 (
            .O(N__26980),
            .I(N__26977));
    Odrv4 I__3634 (
            .O(N__26977),
            .I(n1889));
    InMux I__3633 (
            .O(N__26974),
            .I(N__26970));
    InMux I__3632 (
            .O(N__26973),
            .I(N__26967));
    LocalMux I__3631 (
            .O(N__26970),
            .I(N__26964));
    LocalMux I__3630 (
            .O(N__26967),
            .I(N__26961));
    Span4Mux_v I__3629 (
            .O(N__26964),
            .I(N__26955));
    Span4Mux_v I__3628 (
            .O(N__26961),
            .I(N__26955));
    InMux I__3627 (
            .O(N__26960),
            .I(N__26952));
    Odrv4 I__3626 (
            .O(N__26955),
            .I(n1921));
    LocalMux I__3625 (
            .O(N__26952),
            .I(n1921));
    CascadeMux I__3624 (
            .O(N__26947),
            .I(N__26944));
    InMux I__3623 (
            .O(N__26944),
            .I(N__26941));
    LocalMux I__3622 (
            .O(N__26941),
            .I(N__26938));
    Odrv12 I__3621 (
            .O(N__26938),
            .I(n1900));
    CascadeMux I__3620 (
            .O(N__26935),
            .I(N__26932));
    InMux I__3619 (
            .O(N__26932),
            .I(N__26928));
    CascadeMux I__3618 (
            .O(N__26931),
            .I(N__26925));
    LocalMux I__3617 (
            .O(N__26928),
            .I(N__26922));
    InMux I__3616 (
            .O(N__26925),
            .I(N__26919));
    Span4Mux_h I__3615 (
            .O(N__26922),
            .I(N__26916));
    LocalMux I__3614 (
            .O(N__26919),
            .I(n1932));
    Odrv4 I__3613 (
            .O(N__26916),
            .I(n1932));
    CascadeMux I__3612 (
            .O(N__26911),
            .I(n1932_cascade_));
    CascadeMux I__3611 (
            .O(N__26908),
            .I(N__26905));
    InMux I__3610 (
            .O(N__26905),
            .I(N__26901));
    InMux I__3609 (
            .O(N__26904),
            .I(N__26897));
    LocalMux I__3608 (
            .O(N__26901),
            .I(N__26894));
    InMux I__3607 (
            .O(N__26900),
            .I(N__26891));
    LocalMux I__3606 (
            .O(N__26897),
            .I(N__26888));
    Span4Mux_v I__3605 (
            .O(N__26894),
            .I(N__26883));
    LocalMux I__3604 (
            .O(N__26891),
            .I(N__26883));
    Odrv4 I__3603 (
            .O(N__26888),
            .I(n1931));
    Odrv4 I__3602 (
            .O(N__26883),
            .I(n1931));
    InMux I__3601 (
            .O(N__26878),
            .I(N__26875));
    LocalMux I__3600 (
            .O(N__26875),
            .I(n11686));
    CascadeMux I__3599 (
            .O(N__26872),
            .I(N__26868));
    InMux I__3598 (
            .O(N__26871),
            .I(N__26865));
    InMux I__3597 (
            .O(N__26868),
            .I(N__26862));
    LocalMux I__3596 (
            .O(N__26865),
            .I(N__26856));
    LocalMux I__3595 (
            .O(N__26862),
            .I(N__26856));
    InMux I__3594 (
            .O(N__26861),
            .I(N__26853));
    Span4Mux_h I__3593 (
            .O(N__26856),
            .I(N__26850));
    LocalMux I__3592 (
            .O(N__26853),
            .I(n2332));
    Odrv4 I__3591 (
            .O(N__26850),
            .I(n2332));
    CascadeMux I__3590 (
            .O(N__26845),
            .I(n2333_cascade_));
    InMux I__3589 (
            .O(N__26842),
            .I(N__26838));
    CascadeMux I__3588 (
            .O(N__26841),
            .I(N__26835));
    LocalMux I__3587 (
            .O(N__26838),
            .I(N__26832));
    InMux I__3586 (
            .O(N__26835),
            .I(N__26829));
    Span4Mux_h I__3585 (
            .O(N__26832),
            .I(N__26826));
    LocalMux I__3584 (
            .O(N__26829),
            .I(n2331));
    Odrv4 I__3583 (
            .O(N__26826),
            .I(n2331));
    CascadeMux I__3582 (
            .O(N__26821),
            .I(N__26818));
    InMux I__3581 (
            .O(N__26818),
            .I(N__26815));
    LocalMux I__3580 (
            .O(N__26815),
            .I(n11766));
    CascadeMux I__3579 (
            .O(N__26812),
            .I(N__26809));
    InMux I__3578 (
            .O(N__26809),
            .I(N__26806));
    LocalMux I__3577 (
            .O(N__26806),
            .I(N__26803));
    Span4Mux_v I__3576 (
            .O(N__26803),
            .I(N__26800));
    Odrv4 I__3575 (
            .O(N__26800),
            .I(n2190));
    CascadeMux I__3574 (
            .O(N__26797),
            .I(N__26794));
    InMux I__3573 (
            .O(N__26794),
            .I(N__26790));
    CascadeMux I__3572 (
            .O(N__26793),
            .I(N__26787));
    LocalMux I__3571 (
            .O(N__26790),
            .I(N__26784));
    InMux I__3570 (
            .O(N__26787),
            .I(N__26781));
    Span4Mux_h I__3569 (
            .O(N__26784),
            .I(N__26778));
    LocalMux I__3568 (
            .O(N__26781),
            .I(n2133));
    Odrv4 I__3567 (
            .O(N__26778),
            .I(n2133));
    CascadeMux I__3566 (
            .O(N__26773),
            .I(N__26770));
    InMux I__3565 (
            .O(N__26770),
            .I(N__26766));
    InMux I__3564 (
            .O(N__26769),
            .I(N__26763));
    LocalMux I__3563 (
            .O(N__26766),
            .I(N__26759));
    LocalMux I__3562 (
            .O(N__26763),
            .I(N__26756));
    InMux I__3561 (
            .O(N__26762),
            .I(N__26753));
    Span4Mux_s1_h I__3560 (
            .O(N__26759),
            .I(N__26748));
    Span4Mux_h I__3559 (
            .O(N__26756),
            .I(N__26748));
    LocalMux I__3558 (
            .O(N__26753),
            .I(n2129));
    Odrv4 I__3557 (
            .O(N__26748),
            .I(n2129));
    CascadeMux I__3556 (
            .O(N__26743),
            .I(N__26740));
    InMux I__3555 (
            .O(N__26740),
            .I(N__26736));
    InMux I__3554 (
            .O(N__26739),
            .I(N__26733));
    LocalMux I__3553 (
            .O(N__26736),
            .I(N__26729));
    LocalMux I__3552 (
            .O(N__26733),
            .I(N__26726));
    InMux I__3551 (
            .O(N__26732),
            .I(N__26723));
    Span4Mux_s3_h I__3550 (
            .O(N__26729),
            .I(N__26718));
    Span4Mux_h I__3549 (
            .O(N__26726),
            .I(N__26718));
    LocalMux I__3548 (
            .O(N__26723),
            .I(n2130));
    Odrv4 I__3547 (
            .O(N__26718),
            .I(n2130));
    CascadeMux I__3546 (
            .O(N__26713),
            .I(n11616_cascade_));
    CascadeMux I__3545 (
            .O(N__26710),
            .I(N__26706));
    InMux I__3544 (
            .O(N__26709),
            .I(N__26703));
    InMux I__3543 (
            .O(N__26706),
            .I(N__26700));
    LocalMux I__3542 (
            .O(N__26703),
            .I(N__26697));
    LocalMux I__3541 (
            .O(N__26700),
            .I(N__26694));
    Span4Mux_h I__3540 (
            .O(N__26697),
            .I(N__26688));
    Span4Mux_s3_h I__3539 (
            .O(N__26694),
            .I(N__26688));
    InMux I__3538 (
            .O(N__26693),
            .I(N__26685));
    Odrv4 I__3537 (
            .O(N__26688),
            .I(n2131));
    LocalMux I__3536 (
            .O(N__26685),
            .I(n2131));
    InMux I__3535 (
            .O(N__26680),
            .I(N__26677));
    LocalMux I__3534 (
            .O(N__26677),
            .I(N__26674));
    Odrv12 I__3533 (
            .O(N__26674),
            .I(n2001));
    CascadeMux I__3532 (
            .O(N__26671),
            .I(N__26668));
    InMux I__3531 (
            .O(N__26668),
            .I(N__26665));
    LocalMux I__3530 (
            .O(N__26665),
            .I(N__26662));
    Span4Mux_h I__3529 (
            .O(N__26662),
            .I(N__26658));
    InMux I__3528 (
            .O(N__26661),
            .I(N__26655));
    Odrv4 I__3527 (
            .O(N__26658),
            .I(n2033));
    LocalMux I__3526 (
            .O(N__26655),
            .I(n2033));
    InMux I__3525 (
            .O(N__26650),
            .I(N__26647));
    LocalMux I__3524 (
            .O(N__26647),
            .I(N__26644));
    Span4Mux_v I__3523 (
            .O(N__26644),
            .I(N__26641));
    Odrv4 I__3522 (
            .O(N__26641),
            .I(n2100));
    CascadeMux I__3521 (
            .O(N__26638),
            .I(n2033_cascade_));
    CascadeMux I__3520 (
            .O(N__26635),
            .I(N__26632));
    InMux I__3519 (
            .O(N__26632),
            .I(N__26629));
    LocalMux I__3518 (
            .O(N__26629),
            .I(N__26626));
    Span4Mux_s1_h I__3517 (
            .O(N__26626),
            .I(N__26623));
    Span4Mux_v I__3516 (
            .O(N__26623),
            .I(N__26619));
    InMux I__3515 (
            .O(N__26622),
            .I(N__26616));
    Odrv4 I__3514 (
            .O(N__26619),
            .I(n2132));
    LocalMux I__3513 (
            .O(N__26616),
            .I(n2132));
    InMux I__3512 (
            .O(N__26611),
            .I(N__26608));
    LocalMux I__3511 (
            .O(N__26608),
            .I(N__26605));
    Span4Mux_v I__3510 (
            .O(N__26605),
            .I(N__26602));
    Odrv4 I__3509 (
            .O(N__26602),
            .I(n2199));
    CascadeMux I__3508 (
            .O(N__26599),
            .I(n2132_cascade_));
    InMux I__3507 (
            .O(N__26596),
            .I(N__26593));
    LocalMux I__3506 (
            .O(N__26593),
            .I(N__26589));
    InMux I__3505 (
            .O(N__26592),
            .I(N__26586));
    Odrv4 I__3504 (
            .O(N__26589),
            .I(n2314));
    LocalMux I__3503 (
            .O(N__26586),
            .I(n2314));
    InMux I__3502 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__3501 (
            .O(N__26578),
            .I(N__26575));
    Odrv4 I__3500 (
            .O(N__26575),
            .I(n2381));
    CascadeMux I__3499 (
            .O(N__26572),
            .I(n2314_cascade_));
    CascadeMux I__3498 (
            .O(N__26569),
            .I(n2326_cascade_));
    InMux I__3497 (
            .O(N__26566),
            .I(N__26563));
    LocalMux I__3496 (
            .O(N__26563),
            .I(N__26560));
    Span4Mux_h I__3495 (
            .O(N__26560),
            .I(N__26557));
    Odrv4 I__3494 (
            .O(N__26557),
            .I(n2393));
    InMux I__3493 (
            .O(N__26554),
            .I(N__26551));
    LocalMux I__3492 (
            .O(N__26551),
            .I(N__26548));
    Span4Mux_v I__3491 (
            .O(N__26548),
            .I(N__26545));
    Odrv4 I__3490 (
            .O(N__26545),
            .I(n2400));
    InMux I__3489 (
            .O(N__26542),
            .I(N__26539));
    LocalMux I__3488 (
            .O(N__26539),
            .I(n14194));
    CascadeMux I__3487 (
            .O(N__26536),
            .I(n2247_cascade_));
    CascadeMux I__3486 (
            .O(N__26533),
            .I(N__26530));
    InMux I__3485 (
            .O(N__26530),
            .I(N__26526));
    CascadeMux I__3484 (
            .O(N__26529),
            .I(N__26523));
    LocalMux I__3483 (
            .O(N__26526),
            .I(N__26520));
    InMux I__3482 (
            .O(N__26523),
            .I(N__26517));
    Span4Mux_h I__3481 (
            .O(N__26520),
            .I(N__26514));
    LocalMux I__3480 (
            .O(N__26517),
            .I(n2333));
    Odrv4 I__3479 (
            .O(N__26514),
            .I(n2333));
    CascadeMux I__3478 (
            .O(N__26509),
            .I(n2517_cascade_));
    InMux I__3477 (
            .O(N__26506),
            .I(N__26503));
    LocalMux I__3476 (
            .O(N__26503),
            .I(n13804));
    CascadeMux I__3475 (
            .O(N__26500),
            .I(N__26497));
    InMux I__3474 (
            .O(N__26497),
            .I(N__26494));
    LocalMux I__3473 (
            .O(N__26494),
            .I(N__26491));
    Odrv12 I__3472 (
            .O(N__26491),
            .I(n2185));
    InMux I__3471 (
            .O(N__26488),
            .I(N__26485));
    LocalMux I__3470 (
            .O(N__26485),
            .I(N__26482));
    Span4Mux_h I__3469 (
            .O(N__26482),
            .I(N__26479));
    Odrv4 I__3468 (
            .O(N__26479),
            .I(n2390));
    InMux I__3467 (
            .O(N__26476),
            .I(N__26473));
    LocalMux I__3466 (
            .O(N__26473),
            .I(N__26470));
    Span4Mux_h I__3465 (
            .O(N__26470),
            .I(N__26467));
    Odrv4 I__3464 (
            .O(N__26467),
            .I(n2401));
    CascadeMux I__3463 (
            .O(N__26464),
            .I(n2433_cascade_));
    InMux I__3462 (
            .O(N__26461),
            .I(N__26458));
    LocalMux I__3461 (
            .O(N__26458),
            .I(n11670));
    CascadeMux I__3460 (
            .O(N__26455),
            .I(N__26452));
    InMux I__3459 (
            .O(N__26452),
            .I(N__26449));
    LocalMux I__3458 (
            .O(N__26449),
            .I(N__26446));
    Odrv4 I__3457 (
            .O(N__26446),
            .I(n2383));
    CascadeMux I__3456 (
            .O(N__26443),
            .I(n2527_cascade_));
    InMux I__3455 (
            .O(N__26440),
            .I(N__26437));
    LocalMux I__3454 (
            .O(N__26437),
            .I(n13798));
    CascadeMux I__3453 (
            .O(N__26434),
            .I(n13796_cascade_));
    CascadeMux I__3452 (
            .O(N__26431),
            .I(n14354_cascade_));
    InMux I__3451 (
            .O(N__26428),
            .I(N__26425));
    LocalMux I__3450 (
            .O(N__26425),
            .I(n14220));
    CascadeMux I__3449 (
            .O(N__26422),
            .I(n14224_cascade_));
    CascadeMux I__3448 (
            .O(N__26419),
            .I(n2445_cascade_));
    CascadeMux I__3447 (
            .O(N__26416),
            .I(n1158_cascade_));
    InMux I__3446 (
            .O(N__26413),
            .I(N__26410));
    LocalMux I__3445 (
            .O(N__26410),
            .I(N__26407));
    Odrv4 I__3444 (
            .O(N__26407),
            .I(n1199));
    InMux I__3443 (
            .O(N__26404),
            .I(N__26401));
    LocalMux I__3442 (
            .O(N__26401),
            .I(N__26398));
    Odrv4 I__3441 (
            .O(N__26398),
            .I(n1197));
    CascadeMux I__3440 (
            .O(N__26395),
            .I(N__26392));
    InMux I__3439 (
            .O(N__26392),
            .I(N__26388));
    CascadeMux I__3438 (
            .O(N__26391),
            .I(N__26385));
    LocalMux I__3437 (
            .O(N__26388),
            .I(N__26382));
    InMux I__3436 (
            .O(N__26385),
            .I(N__26379));
    Span4Mux_v I__3435 (
            .O(N__26382),
            .I(N__26376));
    LocalMux I__3434 (
            .O(N__26379),
            .I(n1130));
    Odrv4 I__3433 (
            .O(N__26376),
            .I(n1130));
    CascadeMux I__3432 (
            .O(N__26371),
            .I(n1130_cascade_));
    CascadeMux I__3431 (
            .O(N__26368),
            .I(N__26365));
    InMux I__3430 (
            .O(N__26365),
            .I(N__26362));
    LocalMux I__3429 (
            .O(N__26362),
            .I(n14068));
    InMux I__3428 (
            .O(N__26359),
            .I(N__26356));
    LocalMux I__3427 (
            .O(N__26356),
            .I(n11706));
    CascadeMux I__3426 (
            .O(N__26353),
            .I(N__26349));
    InMux I__3425 (
            .O(N__26352),
            .I(N__26346));
    InMux I__3424 (
            .O(N__26349),
            .I(N__26343));
    LocalMux I__3423 (
            .O(N__26346),
            .I(N__26340));
    LocalMux I__3422 (
            .O(N__26343),
            .I(N__26335));
    Span4Mux_v I__3421 (
            .O(N__26340),
            .I(N__26335));
    Odrv4 I__3420 (
            .O(N__26335),
            .I(n1224));
    CascadeMux I__3419 (
            .O(N__26332),
            .I(n1257_cascade_));
    InMux I__3418 (
            .O(N__26329),
            .I(N__26326));
    LocalMux I__3417 (
            .O(N__26326),
            .I(N__26323));
    Span4Mux_v I__3416 (
            .O(N__26323),
            .I(N__26320));
    Odrv4 I__3415 (
            .O(N__26320),
            .I(n1201));
    InMux I__3414 (
            .O(N__26317),
            .I(N__26314));
    LocalMux I__3413 (
            .O(N__26314),
            .I(n1300));
    CascadeMux I__3412 (
            .O(N__26311),
            .I(n1233_cascade_));
    InMux I__3411 (
            .O(N__26308),
            .I(N__26304));
    CascadeMux I__3410 (
            .O(N__26307),
            .I(N__26301));
    LocalMux I__3409 (
            .O(N__26304),
            .I(N__26297));
    InMux I__3408 (
            .O(N__26301),
            .I(N__26294));
    InMux I__3407 (
            .O(N__26300),
            .I(N__26291));
    Odrv4 I__3406 (
            .O(N__26297),
            .I(n1332));
    LocalMux I__3405 (
            .O(N__26294),
            .I(n1332));
    LocalMux I__3404 (
            .O(N__26291),
            .I(n1332));
    InMux I__3403 (
            .O(N__26284),
            .I(N__26281));
    LocalMux I__3402 (
            .O(N__26281),
            .I(n1296));
    InMux I__3401 (
            .O(N__26278),
            .I(N__26275));
    LocalMux I__3400 (
            .O(N__26275),
            .I(N__26272));
    Odrv12 I__3399 (
            .O(N__26272),
            .I(n1194));
    InMux I__3398 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__3397 (
            .O(N__26266),
            .I(N__26263));
    Odrv12 I__3396 (
            .O(N__26263),
            .I(n1200));
    CascadeMux I__3395 (
            .O(N__26260),
            .I(N__26257));
    InMux I__3394 (
            .O(N__26257),
            .I(N__26253));
    CascadeMux I__3393 (
            .O(N__26256),
            .I(N__26249));
    LocalMux I__3392 (
            .O(N__26253),
            .I(N__26246));
    InMux I__3391 (
            .O(N__26252),
            .I(N__26243));
    InMux I__3390 (
            .O(N__26249),
            .I(N__26240));
    Span4Mux_h I__3389 (
            .O(N__26246),
            .I(N__26237));
    LocalMux I__3388 (
            .O(N__26243),
            .I(n1225));
    LocalMux I__3387 (
            .O(N__26240),
            .I(n1225));
    Odrv4 I__3386 (
            .O(N__26237),
            .I(n1225));
    CascadeMux I__3385 (
            .O(N__26230),
            .I(N__26227));
    InMux I__3384 (
            .O(N__26227),
            .I(N__26224));
    LocalMux I__3383 (
            .O(N__26224),
            .I(n1292));
    InMux I__3382 (
            .O(N__26221),
            .I(N__26217));
    InMux I__3381 (
            .O(N__26220),
            .I(N__26213));
    LocalMux I__3380 (
            .O(N__26217),
            .I(N__26210));
    InMux I__3379 (
            .O(N__26216),
            .I(N__26207));
    LocalMux I__3378 (
            .O(N__26213),
            .I(N__26204));
    Odrv4 I__3377 (
            .O(N__26210),
            .I(n1324));
    LocalMux I__3376 (
            .O(N__26207),
            .I(n1324));
    Odrv4 I__3375 (
            .O(N__26204),
            .I(n1324));
    CascadeMux I__3374 (
            .O(N__26197),
            .I(n11640_cascade_));
    CascadeMux I__3373 (
            .O(N__26194),
            .I(N__26191));
    InMux I__3372 (
            .O(N__26191),
            .I(N__26188));
    LocalMux I__3371 (
            .O(N__26188),
            .I(N__26184));
    CascadeMux I__3370 (
            .O(N__26187),
            .I(N__26180));
    Span4Mux_s2_h I__3369 (
            .O(N__26184),
            .I(N__26177));
    InMux I__3368 (
            .O(N__26183),
            .I(N__26174));
    InMux I__3367 (
            .O(N__26180),
            .I(N__26171));
    Odrv4 I__3366 (
            .O(N__26177),
            .I(n1331));
    LocalMux I__3365 (
            .O(N__26174),
            .I(n1331));
    LocalMux I__3364 (
            .O(N__26171),
            .I(n1331));
    CascadeMux I__3363 (
            .O(N__26164),
            .I(N__26161));
    InMux I__3362 (
            .O(N__26161),
            .I(N__26157));
    InMux I__3361 (
            .O(N__26160),
            .I(N__26154));
    LocalMux I__3360 (
            .O(N__26157),
            .I(N__26149));
    LocalMux I__3359 (
            .O(N__26154),
            .I(N__26149));
    Odrv4 I__3358 (
            .O(N__26149),
            .I(n1323));
    CascadeMux I__3357 (
            .O(N__26146),
            .I(n13315_cascade_));
    CascadeMux I__3356 (
            .O(N__26143),
            .I(n1356_cascade_));
    InMux I__3355 (
            .O(N__26140),
            .I(N__26137));
    LocalMux I__3354 (
            .O(N__26137),
            .I(n1392));
    CascadeMux I__3353 (
            .O(N__26134),
            .I(N__26130));
    InMux I__3352 (
            .O(N__26133),
            .I(N__26125));
    InMux I__3351 (
            .O(N__26130),
            .I(N__26125));
    LocalMux I__3350 (
            .O(N__26125),
            .I(N__26122));
    Span4Mux_v I__3349 (
            .O(N__26122),
            .I(N__26118));
    InMux I__3348 (
            .O(N__26121),
            .I(N__26115));
    Odrv4 I__3347 (
            .O(N__26118),
            .I(n1424));
    LocalMux I__3346 (
            .O(N__26115),
            .I(n1424));
    InMux I__3345 (
            .O(N__26110),
            .I(N__26105));
    InMux I__3344 (
            .O(N__26109),
            .I(N__26102));
    InMux I__3343 (
            .O(N__26108),
            .I(N__26099));
    LocalMux I__3342 (
            .O(N__26105),
            .I(n299));
    LocalMux I__3341 (
            .O(N__26102),
            .I(n299));
    LocalMux I__3340 (
            .O(N__26099),
            .I(n299));
    CascadeMux I__3339 (
            .O(N__26092),
            .I(N__26087));
    InMux I__3338 (
            .O(N__26091),
            .I(N__26082));
    InMux I__3337 (
            .O(N__26090),
            .I(N__26082));
    InMux I__3336 (
            .O(N__26087),
            .I(N__26079));
    LocalMux I__3335 (
            .O(N__26082),
            .I(n1330));
    LocalMux I__3334 (
            .O(N__26079),
            .I(n1330));
    CascadeMux I__3333 (
            .O(N__26074),
            .I(N__26071));
    InMux I__3332 (
            .O(N__26071),
            .I(N__26068));
    LocalMux I__3331 (
            .O(N__26068),
            .I(n1397));
    CascadeMux I__3330 (
            .O(N__26065),
            .I(N__26062));
    InMux I__3329 (
            .O(N__26062),
            .I(N__26058));
    InMux I__3328 (
            .O(N__26061),
            .I(N__26055));
    LocalMux I__3327 (
            .O(N__26058),
            .I(N__26051));
    LocalMux I__3326 (
            .O(N__26055),
            .I(N__26048));
    InMux I__3325 (
            .O(N__26054),
            .I(N__26045));
    Span4Mux_s3_h I__3324 (
            .O(N__26051),
            .I(N__26042));
    Span4Mux_s3_h I__3323 (
            .O(N__26048),
            .I(N__26039));
    LocalMux I__3322 (
            .O(N__26045),
            .I(n1429));
    Odrv4 I__3321 (
            .O(N__26042),
            .I(n1429));
    Odrv4 I__3320 (
            .O(N__26039),
            .I(n1429));
    InMux I__3319 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__3318 (
            .O(N__26029),
            .I(n1297));
    CascadeMux I__3317 (
            .O(N__26026),
            .I(N__26023));
    InMux I__3316 (
            .O(N__26023),
            .I(N__26020));
    LocalMux I__3315 (
            .O(N__26020),
            .I(N__26015));
    InMux I__3314 (
            .O(N__26019),
            .I(N__26012));
    InMux I__3313 (
            .O(N__26018),
            .I(N__26009));
    Odrv4 I__3312 (
            .O(N__26015),
            .I(n1329));
    LocalMux I__3311 (
            .O(N__26012),
            .I(n1329));
    LocalMux I__3310 (
            .O(N__26009),
            .I(n1329));
    InMux I__3309 (
            .O(N__26002),
            .I(N__25999));
    LocalMux I__3308 (
            .O(N__25999),
            .I(n1295));
    InMux I__3307 (
            .O(N__25996),
            .I(N__25993));
    LocalMux I__3306 (
            .O(N__25993),
            .I(n1294));
    InMux I__3305 (
            .O(N__25990),
            .I(N__25987));
    LocalMux I__3304 (
            .O(N__25987),
            .I(N__25984));
    Odrv4 I__3303 (
            .O(N__25984),
            .I(n1393));
    InMux I__3302 (
            .O(N__25981),
            .I(N__25978));
    LocalMux I__3301 (
            .O(N__25978),
            .I(N__25975));
    Odrv4 I__3300 (
            .O(N__25975),
            .I(n1394));
    CascadeMux I__3299 (
            .O(N__25972),
            .I(N__25969));
    InMux I__3298 (
            .O(N__25969),
            .I(N__25965));
    InMux I__3297 (
            .O(N__25968),
            .I(N__25961));
    LocalMux I__3296 (
            .O(N__25965),
            .I(N__25958));
    InMux I__3295 (
            .O(N__25964),
            .I(N__25955));
    LocalMux I__3294 (
            .O(N__25961),
            .I(n1426));
    Odrv4 I__3293 (
            .O(N__25958),
            .I(n1426));
    LocalMux I__3292 (
            .O(N__25955),
            .I(n1426));
    InMux I__3291 (
            .O(N__25948),
            .I(N__25945));
    LocalMux I__3290 (
            .O(N__25945),
            .I(n1399));
    CascadeMux I__3289 (
            .O(N__25942),
            .I(N__25939));
    InMux I__3288 (
            .O(N__25939),
            .I(N__25935));
    InMux I__3287 (
            .O(N__25938),
            .I(N__25931));
    LocalMux I__3286 (
            .O(N__25935),
            .I(N__25928));
    InMux I__3285 (
            .O(N__25934),
            .I(N__25925));
    LocalMux I__3284 (
            .O(N__25931),
            .I(N__25922));
    Span4Mux_s3_h I__3283 (
            .O(N__25928),
            .I(N__25919));
    LocalMux I__3282 (
            .O(N__25925),
            .I(n1431));
    Odrv4 I__3281 (
            .O(N__25922),
            .I(n1431));
    Odrv4 I__3280 (
            .O(N__25919),
            .I(n1431));
    CascadeMux I__3279 (
            .O(N__25912),
            .I(N__25909));
    InMux I__3278 (
            .O(N__25909),
            .I(N__25906));
    LocalMux I__3277 (
            .O(N__25906),
            .I(N__25903));
    Odrv4 I__3276 (
            .O(N__25903),
            .I(n1391));
    CascadeMux I__3275 (
            .O(N__25900),
            .I(N__25897));
    InMux I__3274 (
            .O(N__25897),
            .I(N__25893));
    InMux I__3273 (
            .O(N__25896),
            .I(N__25890));
    LocalMux I__3272 (
            .O(N__25893),
            .I(N__25887));
    LocalMux I__3271 (
            .O(N__25890),
            .I(n1423));
    Odrv4 I__3270 (
            .O(N__25887),
            .I(n1423));
    InMux I__3269 (
            .O(N__25882),
            .I(N__25878));
    InMux I__3268 (
            .O(N__25881),
            .I(N__25875));
    LocalMux I__3267 (
            .O(N__25878),
            .I(N__25872));
    LocalMux I__3266 (
            .O(N__25875),
            .I(N__25869));
    Odrv4 I__3265 (
            .O(N__25872),
            .I(n1422));
    Odrv4 I__3264 (
            .O(N__25869),
            .I(n1422));
    InMux I__3263 (
            .O(N__25864),
            .I(N__25861));
    LocalMux I__3262 (
            .O(N__25861),
            .I(N__25858));
    Odrv4 I__3261 (
            .O(N__25858),
            .I(n13334));
    CascadeMux I__3260 (
            .O(N__25855),
            .I(n1423_cascade_));
    InMux I__3259 (
            .O(N__25852),
            .I(N__25849));
    LocalMux I__3258 (
            .O(N__25849),
            .I(n14094));
    InMux I__3257 (
            .O(N__25846),
            .I(N__25841));
    CascadeMux I__3256 (
            .O(N__25845),
            .I(N__25838));
    InMux I__3255 (
            .O(N__25844),
            .I(N__25835));
    LocalMux I__3254 (
            .O(N__25841),
            .I(N__25832));
    InMux I__3253 (
            .O(N__25838),
            .I(N__25829));
    LocalMux I__3252 (
            .O(N__25835),
            .I(n1425));
    Odrv4 I__3251 (
            .O(N__25832),
            .I(n1425));
    LocalMux I__3250 (
            .O(N__25829),
            .I(n1425));
    CascadeMux I__3249 (
            .O(N__25822),
            .I(n1455_cascade_));
    InMux I__3248 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__3247 (
            .O(N__25816),
            .I(N__25813));
    Odrv12 I__3246 (
            .O(N__25813),
            .I(n1492));
    InMux I__3245 (
            .O(N__25810),
            .I(N__25806));
    CascadeMux I__3244 (
            .O(N__25809),
            .I(N__25803));
    LocalMux I__3243 (
            .O(N__25806),
            .I(N__25799));
    InMux I__3242 (
            .O(N__25803),
            .I(N__25796));
    InMux I__3241 (
            .O(N__25802),
            .I(N__25793));
    Odrv4 I__3240 (
            .O(N__25799),
            .I(n1524));
    LocalMux I__3239 (
            .O(N__25796),
            .I(n1524));
    LocalMux I__3238 (
            .O(N__25793),
            .I(n1524));
    InMux I__3237 (
            .O(N__25786),
            .I(N__25783));
    LocalMux I__3236 (
            .O(N__25783),
            .I(N__25780));
    Odrv4 I__3235 (
            .O(N__25780),
            .I(n1301));
    CascadeMux I__3234 (
            .O(N__25777),
            .I(N__25773));
    InMux I__3233 (
            .O(N__25776),
            .I(N__25770));
    InMux I__3232 (
            .O(N__25773),
            .I(N__25767));
    LocalMux I__3231 (
            .O(N__25770),
            .I(n1333));
    LocalMux I__3230 (
            .O(N__25767),
            .I(n1333));
    CascadeMux I__3229 (
            .O(N__25762),
            .I(n1333_cascade_));
    CascadeMux I__3228 (
            .O(N__25759),
            .I(N__25756));
    InMux I__3227 (
            .O(N__25756),
            .I(N__25753));
    LocalMux I__3226 (
            .O(N__25753),
            .I(N__25750));
    Span4Mux_s3_h I__3225 (
            .O(N__25750),
            .I(N__25747));
    Odrv4 I__3224 (
            .O(N__25747),
            .I(n1592));
    InMux I__3223 (
            .O(N__25744),
            .I(n12172));
    InMux I__3222 (
            .O(N__25741),
            .I(N__25738));
    LocalMux I__3221 (
            .O(N__25738),
            .I(n1591));
    InMux I__3220 (
            .O(N__25735),
            .I(n12173));
    CascadeMux I__3219 (
            .O(N__25732),
            .I(N__25729));
    InMux I__3218 (
            .O(N__25729),
            .I(N__25726));
    LocalMux I__3217 (
            .O(N__25726),
            .I(N__25721));
    InMux I__3216 (
            .O(N__25725),
            .I(N__25718));
    InMux I__3215 (
            .O(N__25724),
            .I(N__25715));
    Span4Mux_h I__3214 (
            .O(N__25721),
            .I(N__25712));
    LocalMux I__3213 (
            .O(N__25718),
            .I(N__25709));
    LocalMux I__3212 (
            .O(N__25715),
            .I(n1523));
    Odrv4 I__3211 (
            .O(N__25712),
            .I(n1523));
    Odrv4 I__3210 (
            .O(N__25709),
            .I(n1523));
    CascadeMux I__3209 (
            .O(N__25702),
            .I(N__25699));
    InMux I__3208 (
            .O(N__25699),
            .I(N__25696));
    LocalMux I__3207 (
            .O(N__25696),
            .I(n1590));
    InMux I__3206 (
            .O(N__25693),
            .I(n12174));
    InMux I__3205 (
            .O(N__25690),
            .I(N__25686));
    InMux I__3204 (
            .O(N__25689),
            .I(N__25683));
    LocalMux I__3203 (
            .O(N__25686),
            .I(n1522));
    LocalMux I__3202 (
            .O(N__25683),
            .I(n1522));
    InMux I__3201 (
            .O(N__25678),
            .I(N__25675));
    LocalMux I__3200 (
            .O(N__25675),
            .I(n1589));
    InMux I__3199 (
            .O(N__25672),
            .I(n12175));
    CascadeMux I__3198 (
            .O(N__25669),
            .I(N__25666));
    InMux I__3197 (
            .O(N__25666),
            .I(N__25663));
    LocalMux I__3196 (
            .O(N__25663),
            .I(N__25659));
    InMux I__3195 (
            .O(N__25662),
            .I(N__25656));
    Span4Mux_h I__3194 (
            .O(N__25659),
            .I(N__25653));
    LocalMux I__3193 (
            .O(N__25656),
            .I(N__25650));
    Odrv4 I__3192 (
            .O(N__25653),
            .I(n1521));
    Odrv4 I__3191 (
            .O(N__25650),
            .I(n1521));
    InMux I__3190 (
            .O(N__25645),
            .I(n12176));
    CascadeMux I__3189 (
            .O(N__25642),
            .I(N__25639));
    InMux I__3188 (
            .O(N__25639),
            .I(N__25635));
    InMux I__3187 (
            .O(N__25638),
            .I(N__25632));
    LocalMux I__3186 (
            .O(N__25635),
            .I(N__25629));
    LocalMux I__3185 (
            .O(N__25632),
            .I(N__25626));
    Odrv4 I__3184 (
            .O(N__25629),
            .I(n1620));
    Odrv4 I__3183 (
            .O(N__25626),
            .I(n1620));
    InMux I__3182 (
            .O(N__25621),
            .I(N__25618));
    LocalMux I__3181 (
            .O(N__25618),
            .I(N__25615));
    Span4Mux_v I__3180 (
            .O(N__25615),
            .I(N__25611));
    InMux I__3179 (
            .O(N__25614),
            .I(N__25608));
    Odrv4 I__3178 (
            .O(N__25611),
            .I(n1427));
    LocalMux I__3177 (
            .O(N__25608),
            .I(n1427));
    CascadeMux I__3176 (
            .O(N__25603),
            .I(N__25600));
    InMux I__3175 (
            .O(N__25600),
            .I(N__25597));
    LocalMux I__3174 (
            .O(N__25597),
            .I(N__25594));
    Odrv4 I__3173 (
            .O(N__25594),
            .I(n1494));
    CascadeMux I__3172 (
            .O(N__25591),
            .I(N__25587));
    CascadeMux I__3171 (
            .O(N__25590),
            .I(N__25584));
    InMux I__3170 (
            .O(N__25587),
            .I(N__25580));
    InMux I__3169 (
            .O(N__25584),
            .I(N__25577));
    InMux I__3168 (
            .O(N__25583),
            .I(N__25574));
    LocalMux I__3167 (
            .O(N__25580),
            .I(n1526));
    LocalMux I__3166 (
            .O(N__25577),
            .I(n1526));
    LocalMux I__3165 (
            .O(N__25574),
            .I(n1526));
    CascadeMux I__3164 (
            .O(N__25567),
            .I(N__25564));
    InMux I__3163 (
            .O(N__25564),
            .I(N__25561));
    LocalMux I__3162 (
            .O(N__25561),
            .I(N__25558));
    Odrv4 I__3161 (
            .O(N__25558),
            .I(n1493));
    InMux I__3160 (
            .O(N__25555),
            .I(N__25552));
    LocalMux I__3159 (
            .O(N__25552),
            .I(N__25548));
    CascadeMux I__3158 (
            .O(N__25551),
            .I(N__25545));
    Span4Mux_s3_h I__3157 (
            .O(N__25548),
            .I(N__25541));
    InMux I__3156 (
            .O(N__25545),
            .I(N__25538));
    InMux I__3155 (
            .O(N__25544),
            .I(N__25535));
    Odrv4 I__3154 (
            .O(N__25541),
            .I(n1525));
    LocalMux I__3153 (
            .O(N__25538),
            .I(n1525));
    LocalMux I__3152 (
            .O(N__25535),
            .I(n1525));
    InMux I__3151 (
            .O(N__25528),
            .I(N__25525));
    LocalMux I__3150 (
            .O(N__25525),
            .I(n1396));
    CascadeMux I__3149 (
            .O(N__25522),
            .I(N__25519));
    InMux I__3148 (
            .O(N__25519),
            .I(N__25516));
    LocalMux I__3147 (
            .O(N__25516),
            .I(N__25511));
    InMux I__3146 (
            .O(N__25515),
            .I(N__25508));
    InMux I__3145 (
            .O(N__25514),
            .I(N__25505));
    Span4Mux_v I__3144 (
            .O(N__25511),
            .I(N__25502));
    LocalMux I__3143 (
            .O(N__25508),
            .I(N__25499));
    LocalMux I__3142 (
            .O(N__25505),
            .I(n1428));
    Odrv4 I__3141 (
            .O(N__25502),
            .I(n1428));
    Odrv12 I__3140 (
            .O(N__25499),
            .I(n1428));
    CascadeMux I__3139 (
            .O(N__25492),
            .I(N__25489));
    InMux I__3138 (
            .O(N__25489),
            .I(N__25484));
    InMux I__3137 (
            .O(N__25488),
            .I(N__25479));
    InMux I__3136 (
            .O(N__25487),
            .I(N__25479));
    LocalMux I__3135 (
            .O(N__25484),
            .I(n1533));
    LocalMux I__3134 (
            .O(N__25479),
            .I(n1533));
    CascadeMux I__3133 (
            .O(N__25474),
            .I(N__25471));
    InMux I__3132 (
            .O(N__25471),
            .I(N__25468));
    LocalMux I__3131 (
            .O(N__25468),
            .I(n1600));
    InMux I__3130 (
            .O(N__25465),
            .I(n12164));
    InMux I__3129 (
            .O(N__25462),
            .I(N__25458));
    CascadeMux I__3128 (
            .O(N__25461),
            .I(N__25455));
    LocalMux I__3127 (
            .O(N__25458),
            .I(N__25451));
    InMux I__3126 (
            .O(N__25455),
            .I(N__25448));
    InMux I__3125 (
            .O(N__25454),
            .I(N__25445));
    Span4Mux_s2_h I__3124 (
            .O(N__25451),
            .I(N__25442));
    LocalMux I__3123 (
            .O(N__25448),
            .I(N__25437));
    LocalMux I__3122 (
            .O(N__25445),
            .I(N__25437));
    Odrv4 I__3121 (
            .O(N__25442),
            .I(n1532));
    Odrv4 I__3120 (
            .O(N__25437),
            .I(n1532));
    CascadeMux I__3119 (
            .O(N__25432),
            .I(N__25429));
    InMux I__3118 (
            .O(N__25429),
            .I(N__25426));
    LocalMux I__3117 (
            .O(N__25426),
            .I(N__25423));
    Odrv4 I__3116 (
            .O(N__25423),
            .I(n1599));
    InMux I__3115 (
            .O(N__25420),
            .I(n12165));
    CascadeMux I__3114 (
            .O(N__25417),
            .I(N__25413));
    InMux I__3113 (
            .O(N__25416),
            .I(N__25410));
    InMux I__3112 (
            .O(N__25413),
            .I(N__25407));
    LocalMux I__3111 (
            .O(N__25410),
            .I(n1531));
    LocalMux I__3110 (
            .O(N__25407),
            .I(n1531));
    InMux I__3109 (
            .O(N__25402),
            .I(N__25399));
    LocalMux I__3108 (
            .O(N__25399),
            .I(N__25396));
    Odrv4 I__3107 (
            .O(N__25396),
            .I(n1598));
    InMux I__3106 (
            .O(N__25393),
            .I(n12166));
    CascadeMux I__3105 (
            .O(N__25390),
            .I(N__25386));
    CascadeMux I__3104 (
            .O(N__25389),
            .I(N__25382));
    InMux I__3103 (
            .O(N__25386),
            .I(N__25379));
    InMux I__3102 (
            .O(N__25385),
            .I(N__25374));
    InMux I__3101 (
            .O(N__25382),
            .I(N__25374));
    LocalMux I__3100 (
            .O(N__25379),
            .I(n1530));
    LocalMux I__3099 (
            .O(N__25374),
            .I(n1530));
    InMux I__3098 (
            .O(N__25369),
            .I(N__25366));
    LocalMux I__3097 (
            .O(N__25366),
            .I(N__25363));
    Odrv4 I__3096 (
            .O(N__25363),
            .I(n1597));
    InMux I__3095 (
            .O(N__25360),
            .I(n12167));
    CascadeMux I__3094 (
            .O(N__25357),
            .I(N__25354));
    InMux I__3093 (
            .O(N__25354),
            .I(N__25349));
    InMux I__3092 (
            .O(N__25353),
            .I(N__25344));
    InMux I__3091 (
            .O(N__25352),
            .I(N__25344));
    LocalMux I__3090 (
            .O(N__25349),
            .I(n1529));
    LocalMux I__3089 (
            .O(N__25344),
            .I(n1529));
    CascadeMux I__3088 (
            .O(N__25339),
            .I(N__25336));
    InMux I__3087 (
            .O(N__25336),
            .I(N__25333));
    LocalMux I__3086 (
            .O(N__25333),
            .I(N__25330));
    Odrv4 I__3085 (
            .O(N__25330),
            .I(n1596));
    InMux I__3084 (
            .O(N__25327),
            .I(n12168));
    CascadeMux I__3083 (
            .O(N__25324),
            .I(N__25320));
    InMux I__3082 (
            .O(N__25323),
            .I(N__25317));
    InMux I__3081 (
            .O(N__25320),
            .I(N__25314));
    LocalMux I__3080 (
            .O(N__25317),
            .I(N__25309));
    LocalMux I__3079 (
            .O(N__25314),
            .I(N__25309));
    Odrv4 I__3078 (
            .O(N__25309),
            .I(n1528));
    InMux I__3077 (
            .O(N__25306),
            .I(N__25303));
    LocalMux I__3076 (
            .O(N__25303),
            .I(n1595));
    InMux I__3075 (
            .O(N__25300),
            .I(n12169));
    CascadeMux I__3074 (
            .O(N__25297),
            .I(N__25293));
    InMux I__3073 (
            .O(N__25296),
            .I(N__25290));
    InMux I__3072 (
            .O(N__25293),
            .I(N__25287));
    LocalMux I__3071 (
            .O(N__25290),
            .I(N__25283));
    LocalMux I__3070 (
            .O(N__25287),
            .I(N__25280));
    InMux I__3069 (
            .O(N__25286),
            .I(N__25277));
    Odrv4 I__3068 (
            .O(N__25283),
            .I(n1527));
    Odrv4 I__3067 (
            .O(N__25280),
            .I(n1527));
    LocalMux I__3066 (
            .O(N__25277),
            .I(n1527));
    InMux I__3065 (
            .O(N__25270),
            .I(N__25267));
    LocalMux I__3064 (
            .O(N__25267),
            .I(N__25264));
    Span4Mux_s2_h I__3063 (
            .O(N__25264),
            .I(N__25261));
    Odrv4 I__3062 (
            .O(N__25261),
            .I(n1594));
    InMux I__3061 (
            .O(N__25258),
            .I(n12170));
    InMux I__3060 (
            .O(N__25255),
            .I(N__25252));
    LocalMux I__3059 (
            .O(N__25252),
            .I(n1593));
    InMux I__3058 (
            .O(N__25249),
            .I(bfn_4_27_0_));
    CascadeMux I__3057 (
            .O(N__25246),
            .I(N__25242));
    InMux I__3056 (
            .O(N__25245),
            .I(N__25238));
    InMux I__3055 (
            .O(N__25242),
            .I(N__25235));
    InMux I__3054 (
            .O(N__25241),
            .I(N__25232));
    LocalMux I__3053 (
            .O(N__25238),
            .I(n1725));
    LocalMux I__3052 (
            .O(N__25235),
            .I(n1725));
    LocalMux I__3051 (
            .O(N__25232),
            .I(n1725));
    InMux I__3050 (
            .O(N__25225),
            .I(N__25222));
    LocalMux I__3049 (
            .O(N__25222),
            .I(n1792));
    InMux I__3048 (
            .O(N__25219),
            .I(n12199));
    InMux I__3047 (
            .O(N__25216),
            .I(n12200));
    CascadeMux I__3046 (
            .O(N__25213),
            .I(N__25208));
    CascadeMux I__3045 (
            .O(N__25212),
            .I(N__25205));
    InMux I__3044 (
            .O(N__25211),
            .I(N__25202));
    InMux I__3043 (
            .O(N__25208),
            .I(N__25199));
    InMux I__3042 (
            .O(N__25205),
            .I(N__25196));
    LocalMux I__3041 (
            .O(N__25202),
            .I(n1723));
    LocalMux I__3040 (
            .O(N__25199),
            .I(n1723));
    LocalMux I__3039 (
            .O(N__25196),
            .I(n1723));
    InMux I__3038 (
            .O(N__25189),
            .I(N__25186));
    LocalMux I__3037 (
            .O(N__25186),
            .I(N__25183));
    Span4Mux_v I__3036 (
            .O(N__25183),
            .I(N__25180));
    Odrv4 I__3035 (
            .O(N__25180),
            .I(n1790));
    InMux I__3034 (
            .O(N__25177),
            .I(n12201));
    CascadeMux I__3033 (
            .O(N__25174),
            .I(N__25170));
    InMux I__3032 (
            .O(N__25173),
            .I(N__25166));
    InMux I__3031 (
            .O(N__25170),
            .I(N__25163));
    InMux I__3030 (
            .O(N__25169),
            .I(N__25160));
    LocalMux I__3029 (
            .O(N__25166),
            .I(n1722));
    LocalMux I__3028 (
            .O(N__25163),
            .I(n1722));
    LocalMux I__3027 (
            .O(N__25160),
            .I(n1722));
    CascadeMux I__3026 (
            .O(N__25153),
            .I(N__25150));
    InMux I__3025 (
            .O(N__25150),
            .I(N__25147));
    LocalMux I__3024 (
            .O(N__25147),
            .I(n1789));
    InMux I__3023 (
            .O(N__25144),
            .I(n12202));
    CascadeMux I__3022 (
            .O(N__25141),
            .I(N__25138));
    InMux I__3021 (
            .O(N__25138),
            .I(N__25135));
    LocalMux I__3020 (
            .O(N__25135),
            .I(N__25130));
    InMux I__3019 (
            .O(N__25134),
            .I(N__25125));
    InMux I__3018 (
            .O(N__25133),
            .I(N__25125));
    Odrv4 I__3017 (
            .O(N__25130),
            .I(n1721));
    LocalMux I__3016 (
            .O(N__25125),
            .I(n1721));
    InMux I__3015 (
            .O(N__25120),
            .I(N__25117));
    LocalMux I__3014 (
            .O(N__25117),
            .I(n1788));
    InMux I__3013 (
            .O(N__25114),
            .I(n12203));
    InMux I__3012 (
            .O(N__25111),
            .I(N__25108));
    LocalMux I__3011 (
            .O(N__25108),
            .I(N__25104));
    InMux I__3010 (
            .O(N__25107),
            .I(N__25101));
    Odrv4 I__3009 (
            .O(N__25104),
            .I(n1720));
    LocalMux I__3008 (
            .O(N__25101),
            .I(n1720));
    InMux I__3007 (
            .O(N__25096),
            .I(N__25093));
    LocalMux I__3006 (
            .O(N__25093),
            .I(N__25090));
    Odrv4 I__3005 (
            .O(N__25090),
            .I(n1787));
    InMux I__3004 (
            .O(N__25087),
            .I(n12204));
    InMux I__3003 (
            .O(N__25084),
            .I(N__25081));
    LocalMux I__3002 (
            .O(N__25081),
            .I(N__25077));
    InMux I__3001 (
            .O(N__25080),
            .I(N__25074));
    Span4Mux_v I__3000 (
            .O(N__25077),
            .I(N__25069));
    LocalMux I__2999 (
            .O(N__25074),
            .I(N__25069));
    Span4Mux_h I__2998 (
            .O(N__25069),
            .I(N__25066));
    Odrv4 I__2997 (
            .O(N__25066),
            .I(n1719));
    InMux I__2996 (
            .O(N__25063),
            .I(n12205));
    InMux I__2995 (
            .O(N__25060),
            .I(N__25057));
    LocalMux I__2994 (
            .O(N__25057),
            .I(N__25054));
    Odrv12 I__2993 (
            .O(N__25054),
            .I(n1601));
    InMux I__2992 (
            .O(N__25051),
            .I(bfn_4_26_0_));
    InMux I__2991 (
            .O(N__25048),
            .I(N__25045));
    LocalMux I__2990 (
            .O(N__25045),
            .I(N__25041));
    InMux I__2989 (
            .O(N__25044),
            .I(N__25038));
    Odrv4 I__2988 (
            .O(N__25041),
            .I(n1733));
    LocalMux I__2987 (
            .O(N__25038),
            .I(n1733));
    InMux I__2986 (
            .O(N__25033),
            .I(N__25030));
    LocalMux I__2985 (
            .O(N__25030),
            .I(N__25027));
    Odrv12 I__2984 (
            .O(N__25027),
            .I(n1800));
    InMux I__2983 (
            .O(N__25024),
            .I(n12191));
    CascadeMux I__2982 (
            .O(N__25021),
            .I(N__25018));
    InMux I__2981 (
            .O(N__25018),
            .I(N__25014));
    CascadeMux I__2980 (
            .O(N__25017),
            .I(N__25011));
    LocalMux I__2979 (
            .O(N__25014),
            .I(N__25008));
    InMux I__2978 (
            .O(N__25011),
            .I(N__25005));
    Span4Mux_v I__2977 (
            .O(N__25008),
            .I(N__24999));
    LocalMux I__2976 (
            .O(N__25005),
            .I(N__24999));
    InMux I__2975 (
            .O(N__25004),
            .I(N__24996));
    Odrv4 I__2974 (
            .O(N__24999),
            .I(n1732));
    LocalMux I__2973 (
            .O(N__24996),
            .I(n1732));
    InMux I__2972 (
            .O(N__24991),
            .I(N__24988));
    LocalMux I__2971 (
            .O(N__24988),
            .I(n1799));
    InMux I__2970 (
            .O(N__24985),
            .I(n12192));
    CascadeMux I__2969 (
            .O(N__24982),
            .I(N__24979));
    InMux I__2968 (
            .O(N__24979),
            .I(N__24975));
    InMux I__2967 (
            .O(N__24978),
            .I(N__24972));
    LocalMux I__2966 (
            .O(N__24975),
            .I(N__24969));
    LocalMux I__2965 (
            .O(N__24972),
            .I(n1731));
    Odrv4 I__2964 (
            .O(N__24969),
            .I(n1731));
    CascadeMux I__2963 (
            .O(N__24964),
            .I(N__24961));
    InMux I__2962 (
            .O(N__24961),
            .I(N__24958));
    LocalMux I__2961 (
            .O(N__24958),
            .I(N__24955));
    Span4Mux_s3_h I__2960 (
            .O(N__24955),
            .I(N__24952));
    Odrv4 I__2959 (
            .O(N__24952),
            .I(n1798));
    InMux I__2958 (
            .O(N__24949),
            .I(n12193));
    CascadeMux I__2957 (
            .O(N__24946),
            .I(N__24942));
    CascadeMux I__2956 (
            .O(N__24945),
            .I(N__24939));
    InMux I__2955 (
            .O(N__24942),
            .I(N__24936));
    InMux I__2954 (
            .O(N__24939),
            .I(N__24933));
    LocalMux I__2953 (
            .O(N__24936),
            .I(N__24928));
    LocalMux I__2952 (
            .O(N__24933),
            .I(N__24928));
    Span4Mux_v I__2951 (
            .O(N__24928),
            .I(N__24924));
    InMux I__2950 (
            .O(N__24927),
            .I(N__24921));
    Odrv4 I__2949 (
            .O(N__24924),
            .I(n1730));
    LocalMux I__2948 (
            .O(N__24921),
            .I(n1730));
    InMux I__2947 (
            .O(N__24916),
            .I(N__24913));
    LocalMux I__2946 (
            .O(N__24913),
            .I(n1797));
    InMux I__2945 (
            .O(N__24910),
            .I(n12194));
    InMux I__2944 (
            .O(N__24907),
            .I(n12195));
    CascadeMux I__2943 (
            .O(N__24904),
            .I(N__24900));
    CascadeMux I__2942 (
            .O(N__24903),
            .I(N__24897));
    InMux I__2941 (
            .O(N__24900),
            .I(N__24894));
    InMux I__2940 (
            .O(N__24897),
            .I(N__24891));
    LocalMux I__2939 (
            .O(N__24894),
            .I(N__24888));
    LocalMux I__2938 (
            .O(N__24891),
            .I(N__24885));
    Span4Mux_v I__2937 (
            .O(N__24888),
            .I(N__24882));
    Span4Mux_h I__2936 (
            .O(N__24885),
            .I(N__24879));
    Odrv4 I__2935 (
            .O(N__24882),
            .I(n1728));
    Odrv4 I__2934 (
            .O(N__24879),
            .I(n1728));
    InMux I__2933 (
            .O(N__24874),
            .I(N__24871));
    LocalMux I__2932 (
            .O(N__24871),
            .I(n1795));
    InMux I__2931 (
            .O(N__24868),
            .I(n12196));
    CascadeMux I__2930 (
            .O(N__24865),
            .I(N__24861));
    InMux I__2929 (
            .O(N__24864),
            .I(N__24858));
    InMux I__2928 (
            .O(N__24861),
            .I(N__24855));
    LocalMux I__2927 (
            .O(N__24858),
            .I(N__24852));
    LocalMux I__2926 (
            .O(N__24855),
            .I(N__24849));
    Span4Mux_h I__2925 (
            .O(N__24852),
            .I(N__24845));
    Span4Mux_h I__2924 (
            .O(N__24849),
            .I(N__24842));
    InMux I__2923 (
            .O(N__24848),
            .I(N__24839));
    Odrv4 I__2922 (
            .O(N__24845),
            .I(n1727));
    Odrv4 I__2921 (
            .O(N__24842),
            .I(n1727));
    LocalMux I__2920 (
            .O(N__24839),
            .I(n1727));
    InMux I__2919 (
            .O(N__24832),
            .I(N__24829));
    LocalMux I__2918 (
            .O(N__24829),
            .I(n1794));
    InMux I__2917 (
            .O(N__24826),
            .I(n12197));
    InMux I__2916 (
            .O(N__24823),
            .I(bfn_4_25_0_));
    CascadeMux I__2915 (
            .O(N__24820),
            .I(n1851_cascade_));
    InMux I__2914 (
            .O(N__24817),
            .I(N__24814));
    LocalMux I__2913 (
            .O(N__24814),
            .I(N__24811));
    Span4Mux_h I__2912 (
            .O(N__24811),
            .I(N__24808));
    Odrv4 I__2911 (
            .O(N__24808),
            .I(n1895));
    CascadeMux I__2910 (
            .O(N__24805),
            .I(N__24802));
    InMux I__2909 (
            .O(N__24802),
            .I(N__24799));
    LocalMux I__2908 (
            .O(N__24799),
            .I(N__24795));
    InMux I__2907 (
            .O(N__24798),
            .I(N__24791));
    Span4Mux_s3_h I__2906 (
            .O(N__24795),
            .I(N__24788));
    InMux I__2905 (
            .O(N__24794),
            .I(N__24785));
    LocalMux I__2904 (
            .O(N__24791),
            .I(n1927));
    Odrv4 I__2903 (
            .O(N__24788),
            .I(n1927));
    LocalMux I__2902 (
            .O(N__24785),
            .I(n1927));
    InMux I__2901 (
            .O(N__24778),
            .I(N__24775));
    LocalMux I__2900 (
            .O(N__24775),
            .I(N__24772));
    Span4Mux_h I__2899 (
            .O(N__24772),
            .I(N__24769));
    Odrv4 I__2898 (
            .O(N__24769),
            .I(n1890));
    InMux I__2897 (
            .O(N__24766),
            .I(N__24762));
    InMux I__2896 (
            .O(N__24765),
            .I(N__24759));
    LocalMux I__2895 (
            .O(N__24762),
            .I(N__24754));
    LocalMux I__2894 (
            .O(N__24759),
            .I(N__24754));
    Span4Mux_v I__2893 (
            .O(N__24754),
            .I(N__24751));
    Odrv4 I__2892 (
            .O(N__24751),
            .I(n1922));
    InMux I__2891 (
            .O(N__24748),
            .I(N__24745));
    LocalMux I__2890 (
            .O(N__24745),
            .I(n13772));
    CascadeMux I__2889 (
            .O(N__24742),
            .I(n1922_cascade_));
    InMux I__2888 (
            .O(N__24739),
            .I(N__24736));
    LocalMux I__2887 (
            .O(N__24736),
            .I(n13770));
    InMux I__2886 (
            .O(N__24733),
            .I(N__24730));
    LocalMux I__2885 (
            .O(N__24730),
            .I(N__24726));
    InMux I__2884 (
            .O(N__24729),
            .I(N__24722));
    Span4Mux_v I__2883 (
            .O(N__24726),
            .I(N__24719));
    InMux I__2882 (
            .O(N__24725),
            .I(N__24716));
    LocalMux I__2881 (
            .O(N__24722),
            .I(N__24713));
    Odrv4 I__2880 (
            .O(N__24719),
            .I(n1920));
    LocalMux I__2879 (
            .O(N__24716),
            .I(n1920));
    Odrv4 I__2878 (
            .O(N__24713),
            .I(n1920));
    CascadeMux I__2877 (
            .O(N__24706),
            .I(n13778_cascade_));
    InMux I__2876 (
            .O(N__24703),
            .I(N__24700));
    LocalMux I__2875 (
            .O(N__24700),
            .I(n13782));
    InMux I__2874 (
            .O(N__24697),
            .I(bfn_4_24_0_));
    CascadeMux I__2873 (
            .O(N__24694),
            .I(N__24690));
    CascadeMux I__2872 (
            .O(N__24693),
            .I(N__24687));
    InMux I__2871 (
            .O(N__24690),
            .I(N__24683));
    InMux I__2870 (
            .O(N__24687),
            .I(N__24680));
    InMux I__2869 (
            .O(N__24686),
            .I(N__24677));
    LocalMux I__2868 (
            .O(N__24683),
            .I(n1928));
    LocalMux I__2867 (
            .O(N__24680),
            .I(n1928));
    LocalMux I__2866 (
            .O(N__24677),
            .I(n1928));
    InMux I__2865 (
            .O(N__24670),
            .I(N__24667));
    LocalMux I__2864 (
            .O(N__24667),
            .I(N__24664));
    Odrv4 I__2863 (
            .O(N__24664),
            .I(n1995));
    CascadeMux I__2862 (
            .O(N__24661),
            .I(N__24657));
    InMux I__2861 (
            .O(N__24660),
            .I(N__24654));
    InMux I__2860 (
            .O(N__24657),
            .I(N__24651));
    LocalMux I__2859 (
            .O(N__24654),
            .I(N__24648));
    LocalMux I__2858 (
            .O(N__24651),
            .I(N__24645));
    Span4Mux_v I__2857 (
            .O(N__24648),
            .I(N__24641));
    Span4Mux_s3_h I__2856 (
            .O(N__24645),
            .I(N__24638));
    InMux I__2855 (
            .O(N__24644),
            .I(N__24635));
    Odrv4 I__2854 (
            .O(N__24641),
            .I(n2027));
    Odrv4 I__2853 (
            .O(N__24638),
            .I(n2027));
    LocalMux I__2852 (
            .O(N__24635),
            .I(n2027));
    InMux I__2851 (
            .O(N__24628),
            .I(N__24625));
    LocalMux I__2850 (
            .O(N__24625),
            .I(N__24621));
    InMux I__2849 (
            .O(N__24624),
            .I(N__24617));
    Span4Mux_v I__2848 (
            .O(N__24621),
            .I(N__24614));
    InMux I__2847 (
            .O(N__24620),
            .I(N__24611));
    LocalMux I__2846 (
            .O(N__24617),
            .I(n2023));
    Odrv4 I__2845 (
            .O(N__24614),
            .I(n2023));
    LocalMux I__2844 (
            .O(N__24611),
            .I(n2023));
    CascadeMux I__2843 (
            .O(N__24604),
            .I(N__24601));
    InMux I__2842 (
            .O(N__24601),
            .I(N__24598));
    LocalMux I__2841 (
            .O(N__24598),
            .I(N__24595));
    Odrv4 I__2840 (
            .O(N__24595),
            .I(n2090));
    CascadeMux I__2839 (
            .O(N__24592),
            .I(N__24589));
    InMux I__2838 (
            .O(N__24589),
            .I(N__24585));
    InMux I__2837 (
            .O(N__24588),
            .I(N__24582));
    LocalMux I__2836 (
            .O(N__24585),
            .I(N__24579));
    LocalMux I__2835 (
            .O(N__24582),
            .I(N__24576));
    Span4Mux_v I__2834 (
            .O(N__24579),
            .I(N__24573));
    Odrv12 I__2833 (
            .O(N__24576),
            .I(n2122));
    Odrv4 I__2832 (
            .O(N__24573),
            .I(n2122));
    CascadeMux I__2831 (
            .O(N__24568),
            .I(N__24565));
    InMux I__2830 (
            .O(N__24565),
            .I(N__24562));
    LocalMux I__2829 (
            .O(N__24562),
            .I(N__24558));
    InMux I__2828 (
            .O(N__24561),
            .I(N__24554));
    Span4Mux_s2_h I__2827 (
            .O(N__24558),
            .I(N__24551));
    InMux I__2826 (
            .O(N__24557),
            .I(N__24548));
    LocalMux I__2825 (
            .O(N__24554),
            .I(n2128));
    Odrv4 I__2824 (
            .O(N__24551),
            .I(n2128));
    LocalMux I__2823 (
            .O(N__24548),
            .I(n2128));
    CascadeMux I__2822 (
            .O(N__24541),
            .I(n2122_cascade_));
    InMux I__2821 (
            .O(N__24538),
            .I(N__24534));
    CascadeMux I__2820 (
            .O(N__24537),
            .I(N__24531));
    LocalMux I__2819 (
            .O(N__24534),
            .I(N__24527));
    InMux I__2818 (
            .O(N__24531),
            .I(N__24522));
    InMux I__2817 (
            .O(N__24530),
            .I(N__24522));
    Span4Mux_h I__2816 (
            .O(N__24527),
            .I(N__24519));
    LocalMux I__2815 (
            .O(N__24522),
            .I(n1918));
    Odrv4 I__2814 (
            .O(N__24519),
            .I(n1918));
    CascadeMux I__2813 (
            .O(N__24514),
            .I(N__24510));
    InMux I__2812 (
            .O(N__24513),
            .I(N__24507));
    InMux I__2811 (
            .O(N__24510),
            .I(N__24504));
    LocalMux I__2810 (
            .O(N__24507),
            .I(n1919));
    LocalMux I__2809 (
            .O(N__24504),
            .I(n1919));
    CascadeMux I__2808 (
            .O(N__24499),
            .I(N__24495));
    InMux I__2807 (
            .O(N__24498),
            .I(N__24491));
    InMux I__2806 (
            .O(N__24495),
            .I(N__24488));
    InMux I__2805 (
            .O(N__24494),
            .I(N__24485));
    LocalMux I__2804 (
            .O(N__24491),
            .I(n1926));
    LocalMux I__2803 (
            .O(N__24488),
            .I(n1926));
    LocalMux I__2802 (
            .O(N__24485),
            .I(n1926));
    CascadeMux I__2801 (
            .O(N__24478),
            .I(n1950_cascade_));
    InMux I__2800 (
            .O(N__24475),
            .I(N__24472));
    LocalMux I__2799 (
            .O(N__24472),
            .I(N__24469));
    Odrv4 I__2798 (
            .O(N__24469),
            .I(n1993));
    InMux I__2797 (
            .O(N__24466),
            .I(N__24463));
    LocalMux I__2796 (
            .O(N__24463),
            .I(N__24460));
    Span4Mux_h I__2795 (
            .O(N__24460),
            .I(N__24457));
    Odrv4 I__2794 (
            .O(N__24457),
            .I(n1999));
    CascadeMux I__2793 (
            .O(N__24454),
            .I(N__24450));
    CascadeMux I__2792 (
            .O(N__24453),
            .I(N__24447));
    InMux I__2791 (
            .O(N__24450),
            .I(N__24444));
    InMux I__2790 (
            .O(N__24447),
            .I(N__24441));
    LocalMux I__2789 (
            .O(N__24444),
            .I(N__24438));
    LocalMux I__2788 (
            .O(N__24441),
            .I(N__24435));
    Span12Mux_s3_h I__2787 (
            .O(N__24438),
            .I(N__24432));
    Odrv4 I__2786 (
            .O(N__24435),
            .I(n2031));
    Odrv12 I__2785 (
            .O(N__24432),
            .I(n2031));
    CascadeMux I__2784 (
            .O(N__24427),
            .I(n2031_cascade_));
    InMux I__2783 (
            .O(N__24424),
            .I(N__24421));
    LocalMux I__2782 (
            .O(N__24421),
            .I(n11680));
    InMux I__2781 (
            .O(N__24418),
            .I(N__24415));
    LocalMux I__2780 (
            .O(N__24415),
            .I(N__24412));
    Odrv4 I__2779 (
            .O(N__24412),
            .I(n1992));
    CascadeMux I__2778 (
            .O(N__24409),
            .I(N__24405));
    CascadeMux I__2777 (
            .O(N__24408),
            .I(N__24402));
    InMux I__2776 (
            .O(N__24405),
            .I(N__24398));
    InMux I__2775 (
            .O(N__24402),
            .I(N__24395));
    InMux I__2774 (
            .O(N__24401),
            .I(N__24392));
    LocalMux I__2773 (
            .O(N__24398),
            .I(n1925));
    LocalMux I__2772 (
            .O(N__24395),
            .I(n1925));
    LocalMux I__2771 (
            .O(N__24392),
            .I(n1925));
    CascadeMux I__2770 (
            .O(N__24385),
            .I(N__24382));
    InMux I__2769 (
            .O(N__24382),
            .I(N__24379));
    LocalMux I__2768 (
            .O(N__24379),
            .I(N__24374));
    InMux I__2767 (
            .O(N__24378),
            .I(N__24371));
    InMux I__2766 (
            .O(N__24377),
            .I(N__24368));
    Span4Mux_s2_h I__2765 (
            .O(N__24374),
            .I(N__24365));
    LocalMux I__2764 (
            .O(N__24371),
            .I(N__24362));
    LocalMux I__2763 (
            .O(N__24368),
            .I(n1819));
    Odrv4 I__2762 (
            .O(N__24365),
            .I(n1819));
    Odrv4 I__2761 (
            .O(N__24362),
            .I(n1819));
    InMux I__2760 (
            .O(N__24355),
            .I(N__24352));
    LocalMux I__2759 (
            .O(N__24352),
            .I(n14134));
    InMux I__2758 (
            .O(N__24349),
            .I(N__24346));
    LocalMux I__2757 (
            .O(N__24346),
            .I(N__24343));
    Span4Mux_h I__2756 (
            .O(N__24343),
            .I(N__24340));
    Odrv4 I__2755 (
            .O(N__24340),
            .I(n2187));
    CascadeMux I__2754 (
            .O(N__24337),
            .I(n2219_cascade_));
    CascadeMux I__2753 (
            .O(N__24334),
            .I(N__24330));
    InMux I__2752 (
            .O(N__24333),
            .I(N__24326));
    InMux I__2751 (
            .O(N__24330),
            .I(N__24321));
    InMux I__2750 (
            .O(N__24329),
            .I(N__24321));
    LocalMux I__2749 (
            .O(N__24326),
            .I(n2318));
    LocalMux I__2748 (
            .O(N__24321),
            .I(n2318));
    CascadeMux I__2747 (
            .O(N__24316),
            .I(N__24313));
    InMux I__2746 (
            .O(N__24313),
            .I(N__24309));
    InMux I__2745 (
            .O(N__24312),
            .I(N__24305));
    LocalMux I__2744 (
            .O(N__24309),
            .I(N__24302));
    InMux I__2743 (
            .O(N__24308),
            .I(N__24299));
    LocalMux I__2742 (
            .O(N__24305),
            .I(N__24294));
    Span4Mux_s3_h I__2741 (
            .O(N__24302),
            .I(N__24294));
    LocalMux I__2740 (
            .O(N__24299),
            .I(n2330));
    Odrv4 I__2739 (
            .O(N__24294),
            .I(n2330));
    InMux I__2738 (
            .O(N__24289),
            .I(N__24286));
    LocalMux I__2737 (
            .O(N__24286),
            .I(N__24283));
    Span4Mux_v I__2736 (
            .O(N__24283),
            .I(N__24280));
    Odrv4 I__2735 (
            .O(N__24280),
            .I(n2099));
    CascadeMux I__2734 (
            .O(N__24277),
            .I(N__24274));
    InMux I__2733 (
            .O(N__24274),
            .I(N__24271));
    LocalMux I__2732 (
            .O(N__24271),
            .I(N__24268));
    Span4Mux_h I__2731 (
            .O(N__24268),
            .I(N__24265));
    Odrv4 I__2730 (
            .O(N__24265),
            .I(n1997));
    InMux I__2729 (
            .O(N__24262),
            .I(N__24258));
    CascadeMux I__2728 (
            .O(N__24261),
            .I(N__24255));
    LocalMux I__2727 (
            .O(N__24258),
            .I(N__24252));
    InMux I__2726 (
            .O(N__24255),
            .I(N__24249));
    Span4Mux_v I__2725 (
            .O(N__24252),
            .I(N__24246));
    LocalMux I__2724 (
            .O(N__24249),
            .I(n2029));
    Odrv4 I__2723 (
            .O(N__24246),
            .I(n2029));
    CascadeMux I__2722 (
            .O(N__24241),
            .I(N__24237));
    InMux I__2721 (
            .O(N__24240),
            .I(N__24234));
    InMux I__2720 (
            .O(N__24237),
            .I(N__24231));
    LocalMux I__2719 (
            .O(N__24234),
            .I(N__24228));
    LocalMux I__2718 (
            .O(N__24231),
            .I(N__24225));
    Span4Mux_v I__2717 (
            .O(N__24228),
            .I(N__24219));
    Span4Mux_s2_h I__2716 (
            .O(N__24225),
            .I(N__24219));
    InMux I__2715 (
            .O(N__24224),
            .I(N__24216));
    Odrv4 I__2714 (
            .O(N__24219),
            .I(n2030));
    LocalMux I__2713 (
            .O(N__24216),
            .I(n2030));
    CascadeMux I__2712 (
            .O(N__24211),
            .I(n2029_cascade_));
    InMux I__2711 (
            .O(N__24208),
            .I(N__24205));
    LocalMux I__2710 (
            .O(N__24205),
            .I(n14154));
    CascadeMux I__2709 (
            .O(N__24202),
            .I(N__24199));
    InMux I__2708 (
            .O(N__24199),
            .I(N__24196));
    LocalMux I__2707 (
            .O(N__24196),
            .I(N__24193));
    Span4Mux_h I__2706 (
            .O(N__24193),
            .I(N__24190));
    Odrv4 I__2705 (
            .O(N__24190),
            .I(n1990));
    InMux I__2704 (
            .O(N__24187),
            .I(N__24184));
    LocalMux I__2703 (
            .O(N__24184),
            .I(N__24180));
    CascadeMux I__2702 (
            .O(N__24183),
            .I(N__24177));
    Span4Mux_h I__2701 (
            .O(N__24180),
            .I(N__24174));
    InMux I__2700 (
            .O(N__24177),
            .I(N__24171));
    Odrv4 I__2699 (
            .O(N__24174),
            .I(n1923));
    LocalMux I__2698 (
            .O(N__24171),
            .I(n1923));
    InMux I__2697 (
            .O(N__24166),
            .I(N__24162));
    CascadeMux I__2696 (
            .O(N__24165),
            .I(N__24159));
    LocalMux I__2695 (
            .O(N__24162),
            .I(N__24156));
    InMux I__2694 (
            .O(N__24159),
            .I(N__24153));
    Span4Mux_v I__2693 (
            .O(N__24156),
            .I(N__24150));
    LocalMux I__2692 (
            .O(N__24153),
            .I(N__24147));
    Odrv4 I__2691 (
            .O(N__24150),
            .I(n2022));
    Odrv4 I__2690 (
            .O(N__24147),
            .I(n2022));
    CascadeMux I__2689 (
            .O(N__24142),
            .I(n2022_cascade_));
    InMux I__2688 (
            .O(N__24139),
            .I(N__24136));
    LocalMux I__2687 (
            .O(N__24136),
            .I(n14146));
    InMux I__2686 (
            .O(N__24133),
            .I(N__24130));
    LocalMux I__2685 (
            .O(N__24130),
            .I(n14152));
    InMux I__2684 (
            .O(N__24127),
            .I(N__24124));
    LocalMux I__2683 (
            .O(N__24124),
            .I(n2384));
    InMux I__2682 (
            .O(N__24121),
            .I(N__24118));
    LocalMux I__2681 (
            .O(N__24118),
            .I(n2385));
    InMux I__2680 (
            .O(N__24115),
            .I(N__24112));
    LocalMux I__2679 (
            .O(N__24112),
            .I(n2389));
    CascadeMux I__2678 (
            .O(N__24109),
            .I(N__24105));
    InMux I__2677 (
            .O(N__24108),
            .I(N__24101));
    InMux I__2676 (
            .O(N__24105),
            .I(N__24096));
    InMux I__2675 (
            .O(N__24104),
            .I(N__24096));
    LocalMux I__2674 (
            .O(N__24101),
            .I(n2317));
    LocalMux I__2673 (
            .O(N__24096),
            .I(n2317));
    InMux I__2672 (
            .O(N__24091),
            .I(N__24088));
    LocalMux I__2671 (
            .O(N__24088),
            .I(N__24085));
    Odrv12 I__2670 (
            .O(N__24085),
            .I(n14410));
    CascadeMux I__2669 (
            .O(N__24082),
            .I(n11774_cascade_));
    CascadeMux I__2668 (
            .O(N__24079),
            .I(n14188_cascade_));
    CascadeMux I__2667 (
            .O(N__24076),
            .I(n2429_cascade_));
    CascadeMux I__2666 (
            .O(N__24073),
            .I(n14210_cascade_));
    CascadeMux I__2665 (
            .O(N__24070),
            .I(n14214_cascade_));
    InMux I__2664 (
            .O(N__24067),
            .I(N__24064));
    LocalMux I__2663 (
            .O(N__24064),
            .I(n13423));
    InMux I__2662 (
            .O(N__24061),
            .I(N__24058));
    LocalMux I__2661 (
            .O(N__24058),
            .I(n2396));
    CascadeMux I__2660 (
            .O(N__24055),
            .I(N__24050));
    CascadeMux I__2659 (
            .O(N__24054),
            .I(N__24047));
    InMux I__2658 (
            .O(N__24053),
            .I(N__24044));
    InMux I__2657 (
            .O(N__24050),
            .I(N__24041));
    InMux I__2656 (
            .O(N__24047),
            .I(N__24038));
    LocalMux I__2655 (
            .O(N__24044),
            .I(N__24035));
    LocalMux I__2654 (
            .O(N__24041),
            .I(n2329));
    LocalMux I__2653 (
            .O(N__24038),
            .I(n2329));
    Odrv4 I__2652 (
            .O(N__24035),
            .I(n2329));
    CascadeMux I__2651 (
            .O(N__24028),
            .I(n14016_cascade_));
    CascadeMux I__2650 (
            .O(N__24025),
            .I(n14022_cascade_));
    InMux I__2649 (
            .O(N__24022),
            .I(N__24019));
    LocalMux I__2648 (
            .O(N__24019),
            .I(N__24016));
    Odrv4 I__2647 (
            .O(N__24016),
            .I(n2395));
    CascadeMux I__2646 (
            .O(N__24013),
            .I(n2346_cascade_));
    InMux I__2645 (
            .O(N__24010),
            .I(N__24007));
    LocalMux I__2644 (
            .O(N__24007),
            .I(N__24004));
    Odrv4 I__2643 (
            .O(N__24004),
            .I(n1193));
    InMux I__2642 (
            .O(N__24001),
            .I(N__23998));
    LocalMux I__2641 (
            .O(N__23998),
            .I(N__23995));
    Odrv4 I__2640 (
            .O(N__23995),
            .I(n2198));
    CascadeMux I__2639 (
            .O(N__23992),
            .I(n2230_cascade_));
    CascadeMux I__2638 (
            .O(N__23989),
            .I(N__23986));
    InMux I__2637 (
            .O(N__23986),
            .I(N__23983));
    LocalMux I__2636 (
            .O(N__23983),
            .I(N__23980));
    Span4Mux_h I__2635 (
            .O(N__23980),
            .I(N__23977));
    Odrv4 I__2634 (
            .O(N__23977),
            .I(n2189));
    CascadeMux I__2633 (
            .O(N__23974),
            .I(n2221_cascade_));
    CascadeMux I__2632 (
            .O(N__23971),
            .I(n2320_cascade_));
    InMux I__2631 (
            .O(N__23968),
            .I(N__23965));
    LocalMux I__2630 (
            .O(N__23965),
            .I(n2387));
    CascadeMux I__2629 (
            .O(N__23962),
            .I(N__23959));
    InMux I__2628 (
            .O(N__23959),
            .I(N__23956));
    LocalMux I__2627 (
            .O(N__23956),
            .I(n2399));
    InMux I__2626 (
            .O(N__23953),
            .I(N__23950));
    LocalMux I__2625 (
            .O(N__23950),
            .I(n2397));
    InMux I__2624 (
            .O(N__23947),
            .I(n12134));
    InMux I__2623 (
            .O(N__23944),
            .I(n12135));
    InMux I__2622 (
            .O(N__23941),
            .I(n12136));
    InMux I__2621 (
            .O(N__23938),
            .I(n12137));
    InMux I__2620 (
            .O(N__23935),
            .I(bfn_3_32_0_));
    InMux I__2619 (
            .O(N__23932),
            .I(n12139));
    InMux I__2618 (
            .O(N__23929),
            .I(n12140));
    InMux I__2617 (
            .O(N__23926),
            .I(N__23920));
    InMux I__2616 (
            .O(N__23925),
            .I(N__23920));
    LocalMux I__2615 (
            .O(N__23920),
            .I(reg_B_2));
    InMux I__2614 (
            .O(N__23917),
            .I(N__23914));
    LocalMux I__2613 (
            .O(N__23914),
            .I(N__23911));
    Odrv4 I__2612 (
            .O(N__23911),
            .I(\debounce.n6 ));
    CascadeMux I__2611 (
            .O(N__23908),
            .I(N__23904));
    InMux I__2610 (
            .O(N__23907),
            .I(N__23901));
    InMux I__2609 (
            .O(N__23904),
            .I(N__23898));
    LocalMux I__2608 (
            .O(N__23901),
            .I(N__23893));
    LocalMux I__2607 (
            .O(N__23898),
            .I(N__23893));
    Span4Mux_s2_v I__2606 (
            .O(N__23893),
            .I(N__23890));
    Odrv4 I__2605 (
            .O(N__23890),
            .I(\debounce.reg_A_2 ));
    SRMux I__2604 (
            .O(N__23887),
            .I(N__23883));
    SRMux I__2603 (
            .O(N__23886),
            .I(N__23880));
    LocalMux I__2602 (
            .O(N__23883),
            .I(N__23877));
    LocalMux I__2601 (
            .O(N__23880),
            .I(N__23874));
    Span4Mux_v I__2600 (
            .O(N__23877),
            .I(N__23869));
    Span4Mux_v I__2599 (
            .O(N__23874),
            .I(N__23869));
    Odrv4 I__2598 (
            .O(N__23869),
            .I(\debounce.cnt_next_9__N_418 ));
    InMux I__2597 (
            .O(N__23866),
            .I(n12150));
    InMux I__2596 (
            .O(N__23863),
            .I(n12151));
    InMux I__2595 (
            .O(N__23860),
            .I(bfn_3_31_0_));
    InMux I__2594 (
            .O(N__23857),
            .I(n12131));
    CascadeMux I__2593 (
            .O(N__23854),
            .I(N__23851));
    InMux I__2592 (
            .O(N__23851),
            .I(N__23848));
    LocalMux I__2591 (
            .O(N__23848),
            .I(n1299));
    InMux I__2590 (
            .O(N__23845),
            .I(n12132));
    InMux I__2589 (
            .O(N__23842),
            .I(N__23839));
    LocalMux I__2588 (
            .O(N__23839),
            .I(n1298));
    InMux I__2587 (
            .O(N__23836),
            .I(n12133));
    CascadeMux I__2586 (
            .O(N__23833),
            .I(N__23830));
    InMux I__2585 (
            .O(N__23830),
            .I(N__23827));
    LocalMux I__2584 (
            .O(N__23827),
            .I(n1400));
    InMux I__2583 (
            .O(N__23824),
            .I(n12141));
    InMux I__2582 (
            .O(N__23821),
            .I(n12142));
    InMux I__2581 (
            .O(N__23818),
            .I(N__23815));
    LocalMux I__2580 (
            .O(N__23815),
            .I(N__23812));
    Span4Mux_s2_h I__2579 (
            .O(N__23812),
            .I(N__23809));
    Odrv4 I__2578 (
            .O(N__23809),
            .I(n1398));
    InMux I__2577 (
            .O(N__23806),
            .I(n12143));
    InMux I__2576 (
            .O(N__23803),
            .I(n12144));
    InMux I__2575 (
            .O(N__23800),
            .I(n12145));
    InMux I__2574 (
            .O(N__23797),
            .I(N__23794));
    LocalMux I__2573 (
            .O(N__23794),
            .I(N__23791));
    Span4Mux_s2_h I__2572 (
            .O(N__23791),
            .I(N__23788));
    Odrv4 I__2571 (
            .O(N__23788),
            .I(n1395));
    InMux I__2570 (
            .O(N__23785),
            .I(n12146));
    InMux I__2569 (
            .O(N__23782),
            .I(n12147));
    InMux I__2568 (
            .O(N__23779),
            .I(bfn_3_30_0_));
    InMux I__2567 (
            .O(N__23776),
            .I(n12149));
    CascadeMux I__2566 (
            .O(N__23773),
            .I(N__23770));
    InMux I__2565 (
            .O(N__23770),
            .I(N__23767));
    LocalMux I__2564 (
            .O(N__23767),
            .I(n1495));
    InMux I__2563 (
            .O(N__23764),
            .I(N__23761));
    LocalMux I__2562 (
            .O(N__23761),
            .I(n1496));
    CascadeMux I__2561 (
            .O(N__23758),
            .I(n1528_cascade_));
    CascadeMux I__2560 (
            .O(N__23755),
            .I(n13978_cascade_));
    InMux I__2559 (
            .O(N__23752),
            .I(N__23749));
    LocalMux I__2558 (
            .O(N__23749),
            .I(N__23746));
    Odrv4 I__2557 (
            .O(N__23746),
            .I(n13984));
    InMux I__2556 (
            .O(N__23743),
            .I(N__23738));
    CascadeMux I__2555 (
            .O(N__23742),
            .I(N__23735));
    InMux I__2554 (
            .O(N__23741),
            .I(N__23732));
    LocalMux I__2553 (
            .O(N__23738),
            .I(N__23729));
    InMux I__2552 (
            .O(N__23735),
            .I(N__23726));
    LocalMux I__2551 (
            .O(N__23732),
            .I(N__23723));
    Odrv4 I__2550 (
            .O(N__23729),
            .I(n1432));
    LocalMux I__2549 (
            .O(N__23726),
            .I(n1432));
    Odrv4 I__2548 (
            .O(N__23723),
            .I(n1432));
    InMux I__2547 (
            .O(N__23716),
            .I(N__23713));
    LocalMux I__2546 (
            .O(N__23713),
            .I(N__23710));
    Odrv4 I__2545 (
            .O(N__23710),
            .I(n14088));
    CascadeMux I__2544 (
            .O(N__23707),
            .I(N__23703));
    CascadeMux I__2543 (
            .O(N__23706),
            .I(N__23700));
    InMux I__2542 (
            .O(N__23703),
            .I(N__23697));
    InMux I__2541 (
            .O(N__23700),
            .I(N__23694));
    LocalMux I__2540 (
            .O(N__23697),
            .I(N__23691));
    LocalMux I__2539 (
            .O(N__23694),
            .I(n1433));
    Odrv4 I__2538 (
            .O(N__23691),
            .I(n1433));
    CascadeMux I__2537 (
            .O(N__23686),
            .I(n1433_cascade_));
    InMux I__2536 (
            .O(N__23683),
            .I(N__23680));
    LocalMux I__2535 (
            .O(N__23680),
            .I(n1500));
    InMux I__2534 (
            .O(N__23677),
            .I(N__23674));
    LocalMux I__2533 (
            .O(N__23674),
            .I(n1401));
    InMux I__2532 (
            .O(N__23671),
            .I(bfn_3_29_0_));
    CascadeMux I__2531 (
            .O(N__23668),
            .I(N__23665));
    InMux I__2530 (
            .O(N__23665),
            .I(N__23660));
    CascadeMux I__2529 (
            .O(N__23664),
            .I(N__23657));
    InMux I__2528 (
            .O(N__23663),
            .I(N__23654));
    LocalMux I__2527 (
            .O(N__23660),
            .I(N__23651));
    InMux I__2526 (
            .O(N__23657),
            .I(N__23648));
    LocalMux I__2525 (
            .O(N__23654),
            .I(n1627));
    Odrv4 I__2524 (
            .O(N__23651),
            .I(n1627));
    LocalMux I__2523 (
            .O(N__23648),
            .I(n1627));
    InMux I__2522 (
            .O(N__23641),
            .I(N__23638));
    LocalMux I__2521 (
            .O(N__23638),
            .I(N__23635));
    Span4Mux_h I__2520 (
            .O(N__23635),
            .I(N__23631));
    InMux I__2519 (
            .O(N__23634),
            .I(N__23628));
    Odrv4 I__2518 (
            .O(N__23631),
            .I(n1430));
    LocalMux I__2517 (
            .O(N__23628),
            .I(n1430));
    InMux I__2516 (
            .O(N__23623),
            .I(N__23620));
    LocalMux I__2515 (
            .O(N__23620),
            .I(n1497));
    InMux I__2514 (
            .O(N__23617),
            .I(N__23614));
    LocalMux I__2513 (
            .O(N__23614),
            .I(n1498));
    InMux I__2512 (
            .O(N__23611),
            .I(N__23608));
    LocalMux I__2511 (
            .O(N__23608),
            .I(N__23605));
    Span4Mux_v I__2510 (
            .O(N__23605),
            .I(N__23600));
    InMux I__2509 (
            .O(N__23604),
            .I(N__23597));
    InMux I__2508 (
            .O(N__23603),
            .I(N__23594));
    Span4Mux_s1_h I__2507 (
            .O(N__23600),
            .I(N__23591));
    LocalMux I__2506 (
            .O(N__23597),
            .I(N__23588));
    LocalMux I__2505 (
            .O(N__23594),
            .I(N__23585));
    Odrv4 I__2504 (
            .O(N__23591),
            .I(n1622));
    Odrv4 I__2503 (
            .O(N__23588),
            .I(n1622));
    Odrv4 I__2502 (
            .O(N__23585),
            .I(n1622));
    InMux I__2501 (
            .O(N__23578),
            .I(N__23574));
    InMux I__2500 (
            .O(N__23577),
            .I(N__23571));
    LocalMux I__2499 (
            .O(N__23574),
            .I(N__23568));
    LocalMux I__2498 (
            .O(N__23571),
            .I(N__23563));
    Span4Mux_v I__2497 (
            .O(N__23568),
            .I(N__23563));
    Odrv4 I__2496 (
            .O(N__23563),
            .I(n300));
    InMux I__2495 (
            .O(N__23560),
            .I(N__23557));
    LocalMux I__2494 (
            .O(N__23557),
            .I(n1501));
    CascadeMux I__2493 (
            .O(N__23554),
            .I(n300_cascade_));
    InMux I__2492 (
            .O(N__23551),
            .I(N__23548));
    LocalMux I__2491 (
            .O(N__23548),
            .I(N__23545));
    Odrv4 I__2490 (
            .O(N__23545),
            .I(n1490));
    CascadeMux I__2489 (
            .O(N__23542),
            .I(n1522_cascade_));
    CascadeMux I__2488 (
            .O(N__23539),
            .I(N__23536));
    InMux I__2487 (
            .O(N__23536),
            .I(N__23533));
    LocalMux I__2486 (
            .O(N__23533),
            .I(N__23528));
    InMux I__2485 (
            .O(N__23532),
            .I(N__23525));
    InMux I__2484 (
            .O(N__23531),
            .I(N__23522));
    Span4Mux_v I__2483 (
            .O(N__23528),
            .I(N__23519));
    LocalMux I__2482 (
            .O(N__23525),
            .I(N__23516));
    LocalMux I__2481 (
            .O(N__23522),
            .I(N__23513));
    Odrv4 I__2480 (
            .O(N__23519),
            .I(n1621));
    Odrv4 I__2479 (
            .O(N__23516),
            .I(n1621));
    Odrv12 I__2478 (
            .O(N__23513),
            .I(n1621));
    CascadeMux I__2477 (
            .O(N__23506),
            .I(N__23503));
    InMux I__2476 (
            .O(N__23503),
            .I(N__23498));
    InMux I__2475 (
            .O(N__23502),
            .I(N__23493));
    InMux I__2474 (
            .O(N__23501),
            .I(N__23493));
    LocalMux I__2473 (
            .O(N__23498),
            .I(n1626));
    LocalMux I__2472 (
            .O(N__23493),
            .I(n1626));
    CascadeMux I__2471 (
            .O(N__23488),
            .I(N__23485));
    InMux I__2470 (
            .O(N__23485),
            .I(N__23482));
    LocalMux I__2469 (
            .O(N__23482),
            .I(N__23479));
    Span4Mux_h I__2468 (
            .O(N__23479),
            .I(N__23476));
    Odrv4 I__2467 (
            .O(N__23476),
            .I(n1693));
    CascadeMux I__2466 (
            .O(N__23473),
            .I(N__23469));
    InMux I__2465 (
            .O(N__23472),
            .I(N__23466));
    InMux I__2464 (
            .O(N__23469),
            .I(N__23463));
    LocalMux I__2463 (
            .O(N__23466),
            .I(N__23460));
    LocalMux I__2462 (
            .O(N__23463),
            .I(N__23457));
    Odrv4 I__2461 (
            .O(N__23460),
            .I(n1632));
    Odrv4 I__2460 (
            .O(N__23457),
            .I(n1632));
    CascadeMux I__2459 (
            .O(N__23452),
            .I(n1632_cascade_));
    InMux I__2458 (
            .O(N__23449),
            .I(N__23445));
    CascadeMux I__2457 (
            .O(N__23448),
            .I(N__23442));
    LocalMux I__2456 (
            .O(N__23445),
            .I(N__23438));
    InMux I__2455 (
            .O(N__23442),
            .I(N__23435));
    InMux I__2454 (
            .O(N__23441),
            .I(N__23432));
    Odrv4 I__2453 (
            .O(N__23438),
            .I(n1633));
    LocalMux I__2452 (
            .O(N__23435),
            .I(n1633));
    LocalMux I__2451 (
            .O(N__23432),
            .I(n1633));
    InMux I__2450 (
            .O(N__23425),
            .I(N__23422));
    LocalMux I__2449 (
            .O(N__23422),
            .I(n11634));
    CascadeMux I__2448 (
            .O(N__23419),
            .I(N__23416));
    InMux I__2447 (
            .O(N__23416),
            .I(N__23413));
    LocalMux I__2446 (
            .O(N__23413),
            .I(N__23410));
    Span4Mux_s2_h I__2445 (
            .O(N__23410),
            .I(N__23405));
    InMux I__2444 (
            .O(N__23409),
            .I(N__23400));
    InMux I__2443 (
            .O(N__23408),
            .I(N__23400));
    Odrv4 I__2442 (
            .O(N__23405),
            .I(n1625));
    LocalMux I__2441 (
            .O(N__23400),
            .I(n1625));
    CascadeMux I__2440 (
            .O(N__23395),
            .I(N__23392));
    InMux I__2439 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__2438 (
            .O(N__23389),
            .I(N__23384));
    InMux I__2437 (
            .O(N__23388),
            .I(N__23381));
    InMux I__2436 (
            .O(N__23387),
            .I(N__23378));
    Span4Mux_s2_h I__2435 (
            .O(N__23384),
            .I(N__23373));
    LocalMux I__2434 (
            .O(N__23381),
            .I(N__23373));
    LocalMux I__2433 (
            .O(N__23378),
            .I(n1623));
    Odrv4 I__2432 (
            .O(N__23373),
            .I(n1623));
    CascadeMux I__2431 (
            .O(N__23368),
            .I(N__23365));
    InMux I__2430 (
            .O(N__23365),
            .I(N__23362));
    LocalMux I__2429 (
            .O(N__23362),
            .I(n1499));
    CascadeMux I__2428 (
            .O(N__23359),
            .I(n1531_cascade_));
    InMux I__2427 (
            .O(N__23356),
            .I(N__23353));
    LocalMux I__2426 (
            .O(N__23353),
            .I(n11698));
    CascadeMux I__2425 (
            .O(N__23350),
            .I(n14110_cascade_));
    CascadeMux I__2424 (
            .O(N__23347),
            .I(n1653_cascade_));
    InMux I__2423 (
            .O(N__23344),
            .I(N__23341));
    LocalMux I__2422 (
            .O(N__23341),
            .I(N__23338));
    Span4Mux_h I__2421 (
            .O(N__23338),
            .I(N__23335));
    Odrv4 I__2420 (
            .O(N__23335),
            .I(n1691));
    InMux I__2419 (
            .O(N__23332),
            .I(N__23329));
    LocalMux I__2418 (
            .O(N__23329),
            .I(n13962));
    InMux I__2417 (
            .O(N__23326),
            .I(N__23323));
    LocalMux I__2416 (
            .O(N__23323),
            .I(n11694));
    CascadeMux I__2415 (
            .O(N__23320),
            .I(n13968_cascade_));
    InMux I__2414 (
            .O(N__23317),
            .I(N__23314));
    LocalMux I__2413 (
            .O(N__23314),
            .I(n14116));
    CascadeMux I__2412 (
            .O(N__23311),
            .I(N__23308));
    InMux I__2411 (
            .O(N__23308),
            .I(N__23305));
    LocalMux I__2410 (
            .O(N__23305),
            .I(n13972));
    InMux I__2409 (
            .O(N__23302),
            .I(N__23299));
    LocalMux I__2408 (
            .O(N__23299),
            .I(N__23296));
    Span4Mux_v I__2407 (
            .O(N__23296),
            .I(N__23293));
    Odrv4 I__2406 (
            .O(N__23293),
            .I(n1690));
    CascadeMux I__2405 (
            .O(N__23290),
            .I(N__23286));
    CascadeMux I__2404 (
            .O(N__23289),
            .I(N__23283));
    InMux I__2403 (
            .O(N__23286),
            .I(N__23279));
    InMux I__2402 (
            .O(N__23283),
            .I(N__23276));
    InMux I__2401 (
            .O(N__23282),
            .I(N__23273));
    LocalMux I__2400 (
            .O(N__23279),
            .I(n1628));
    LocalMux I__2399 (
            .O(N__23276),
            .I(n1628));
    LocalMux I__2398 (
            .O(N__23273),
            .I(n1628));
    InMux I__2397 (
            .O(N__23266),
            .I(N__23263));
    LocalMux I__2396 (
            .O(N__23263),
            .I(n14104));
    CascadeMux I__2395 (
            .O(N__23260),
            .I(N__23257));
    InMux I__2394 (
            .O(N__23257),
            .I(N__23254));
    LocalMux I__2393 (
            .O(N__23254),
            .I(N__23250));
    CascadeMux I__2392 (
            .O(N__23253),
            .I(N__23246));
    Span4Mux_s2_h I__2391 (
            .O(N__23250),
            .I(N__23243));
    InMux I__2390 (
            .O(N__23249),
            .I(N__23238));
    InMux I__2389 (
            .O(N__23246),
            .I(N__23238));
    Odrv4 I__2388 (
            .O(N__23243),
            .I(n1624));
    LocalMux I__2387 (
            .O(N__23238),
            .I(n1624));
    CascadeMux I__2386 (
            .O(N__23233),
            .I(N__23230));
    InMux I__2385 (
            .O(N__23230),
            .I(N__23227));
    LocalMux I__2384 (
            .O(N__23227),
            .I(N__23224));
    Span4Mux_h I__2383 (
            .O(N__23224),
            .I(N__23221));
    Odrv4 I__2382 (
            .O(N__23221),
            .I(n1692));
    InMux I__2381 (
            .O(N__23218),
            .I(N__23215));
    LocalMux I__2380 (
            .O(N__23215),
            .I(N__23212));
    Odrv4 I__2379 (
            .O(N__23212),
            .I(n1894));
    InMux I__2378 (
            .O(N__23209),
            .I(N__23206));
    LocalMux I__2377 (
            .O(N__23206),
            .I(N__23203));
    Span4Mux_h I__2376 (
            .O(N__23203),
            .I(N__23200));
    Odrv4 I__2375 (
            .O(N__23200),
            .I(n1688));
    CascadeMux I__2374 (
            .O(N__23197),
            .I(n1720_cascade_));
    InMux I__2373 (
            .O(N__23194),
            .I(N__23190));
    CascadeMux I__2372 (
            .O(N__23193),
            .I(N__23187));
    LocalMux I__2371 (
            .O(N__23190),
            .I(N__23184));
    InMux I__2370 (
            .O(N__23187),
            .I(N__23181));
    Span4Mux_v I__2369 (
            .O(N__23184),
            .I(N__23177));
    LocalMux I__2368 (
            .O(N__23181),
            .I(N__23174));
    InMux I__2367 (
            .O(N__23180),
            .I(N__23171));
    Odrv4 I__2366 (
            .O(N__23177),
            .I(n1820));
    Odrv4 I__2365 (
            .O(N__23174),
            .I(n1820));
    LocalMux I__2364 (
            .O(N__23171),
            .I(n1820));
    CascadeMux I__2363 (
            .O(N__23164),
            .I(n1752_cascade_));
    CascadeMux I__2362 (
            .O(N__23161),
            .I(N__23157));
    CascadeMux I__2361 (
            .O(N__23160),
            .I(N__23154));
    InMux I__2360 (
            .O(N__23157),
            .I(N__23151));
    InMux I__2359 (
            .O(N__23154),
            .I(N__23147));
    LocalMux I__2358 (
            .O(N__23151),
            .I(N__23144));
    InMux I__2357 (
            .O(N__23150),
            .I(N__23141));
    LocalMux I__2356 (
            .O(N__23147),
            .I(n1821));
    Odrv4 I__2355 (
            .O(N__23144),
            .I(n1821));
    LocalMux I__2354 (
            .O(N__23141),
            .I(n1821));
    InMux I__2353 (
            .O(N__23134),
            .I(N__23131));
    LocalMux I__2352 (
            .O(N__23131),
            .I(n13343));
    CascadeMux I__2351 (
            .O(N__23128),
            .I(N__23125));
    InMux I__2350 (
            .O(N__23125),
            .I(N__23122));
    LocalMux I__2349 (
            .O(N__23122),
            .I(N__23119));
    Span4Mux_h I__2348 (
            .O(N__23119),
            .I(N__23116));
    Odrv4 I__2347 (
            .O(N__23116),
            .I(n1892));
    CascadeMux I__2346 (
            .O(N__23113),
            .I(N__23109));
    CascadeMux I__2345 (
            .O(N__23112),
            .I(N__23106));
    InMux I__2344 (
            .O(N__23109),
            .I(N__23103));
    InMux I__2343 (
            .O(N__23106),
            .I(N__23100));
    LocalMux I__2342 (
            .O(N__23103),
            .I(n1924));
    LocalMux I__2341 (
            .O(N__23100),
            .I(n1924));
    CascadeMux I__2340 (
            .O(N__23095),
            .I(n1924_cascade_));
    InMux I__2339 (
            .O(N__23092),
            .I(N__23089));
    LocalMux I__2338 (
            .O(N__23089),
            .I(N__23086));
    Span4Mux_h I__2337 (
            .O(N__23086),
            .I(N__23083));
    Odrv4 I__2336 (
            .O(N__23083),
            .I(n1893));
    CascadeMux I__2335 (
            .O(N__23080),
            .I(N__23077));
    InMux I__2334 (
            .O(N__23077),
            .I(N__23074));
    LocalMux I__2333 (
            .O(N__23074),
            .I(N__23071));
    Span4Mux_v I__2332 (
            .O(N__23071),
            .I(N__23068));
    Odrv4 I__2331 (
            .O(N__23068),
            .I(n1891));
    CascadeMux I__2330 (
            .O(N__23065),
            .I(n1923_cascade_));
    CascadeMux I__2329 (
            .O(N__23062),
            .I(N__23059));
    InMux I__2328 (
            .O(N__23059),
            .I(N__23056));
    LocalMux I__2327 (
            .O(N__23056),
            .I(N__23053));
    Span4Mux_h I__2326 (
            .O(N__23053),
            .I(N__23050));
    Odrv4 I__2325 (
            .O(N__23050),
            .I(n1896));
    InMux I__2324 (
            .O(N__23047),
            .I(N__23044));
    LocalMux I__2323 (
            .O(N__23044),
            .I(N__23041));
    Odrv4 I__2322 (
            .O(N__23041),
            .I(n1899));
    CascadeMux I__2321 (
            .O(N__23038),
            .I(n1822_cascade_));
    CascadeMux I__2320 (
            .O(N__23035),
            .I(N__23031));
    CascadeMux I__2319 (
            .O(N__23034),
            .I(N__23028));
    InMux I__2318 (
            .O(N__23031),
            .I(N__23025));
    InMux I__2317 (
            .O(N__23028),
            .I(N__23022));
    LocalMux I__2316 (
            .O(N__23025),
            .I(N__23018));
    LocalMux I__2315 (
            .O(N__23022),
            .I(N__23015));
    InMux I__2314 (
            .O(N__23021),
            .I(N__23012));
    Odrv4 I__2313 (
            .O(N__23018),
            .I(n2028));
    Odrv4 I__2312 (
            .O(N__23015),
            .I(n2028));
    LocalMux I__2311 (
            .O(N__23012),
            .I(n2028));
    CascadeMux I__2310 (
            .O(N__23005),
            .I(N__23002));
    InMux I__2309 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__2308 (
            .O(N__22999),
            .I(n1989));
    InMux I__2307 (
            .O(N__22996),
            .I(N__22993));
    LocalMux I__2306 (
            .O(N__22993),
            .I(n1998));
    CascadeMux I__2305 (
            .O(N__22990),
            .I(N__22987));
    InMux I__2304 (
            .O(N__22987),
            .I(N__22984));
    LocalMux I__2303 (
            .O(N__22984),
            .I(n1994));
    CascadeMux I__2302 (
            .O(N__22981),
            .I(N__22977));
    CascadeMux I__2301 (
            .O(N__22980),
            .I(N__22973));
    InMux I__2300 (
            .O(N__22977),
            .I(N__22970));
    CascadeMux I__2299 (
            .O(N__22976),
            .I(N__22967));
    InMux I__2298 (
            .O(N__22973),
            .I(N__22964));
    LocalMux I__2297 (
            .O(N__22970),
            .I(N__22961));
    InMux I__2296 (
            .O(N__22967),
            .I(N__22958));
    LocalMux I__2295 (
            .O(N__22964),
            .I(n2026));
    Odrv4 I__2294 (
            .O(N__22961),
            .I(n2026));
    LocalMux I__2293 (
            .O(N__22958),
            .I(n2026));
    InMux I__2292 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__2291 (
            .O(N__22948),
            .I(N__22945));
    Span4Mux_h I__2290 (
            .O(N__22945),
            .I(N__22942));
    Odrv4 I__2289 (
            .O(N__22942),
            .I(n1887));
    InMux I__2288 (
            .O(N__22939),
            .I(N__22936));
    LocalMux I__2287 (
            .O(N__22936),
            .I(n1986));
    CascadeMux I__2286 (
            .O(N__22933),
            .I(n1919_cascade_));
    InMux I__2285 (
            .O(N__22930),
            .I(N__22926));
    InMux I__2284 (
            .O(N__22929),
            .I(N__22923));
    LocalMux I__2283 (
            .O(N__22926),
            .I(N__22919));
    LocalMux I__2282 (
            .O(N__22923),
            .I(N__22916));
    InMux I__2281 (
            .O(N__22922),
            .I(N__22913));
    Span4Mux_v I__2280 (
            .O(N__22919),
            .I(N__22910));
    Span4Mux_s3_h I__2279 (
            .O(N__22916),
            .I(N__22907));
    LocalMux I__2278 (
            .O(N__22913),
            .I(n2018));
    Odrv4 I__2277 (
            .O(N__22910),
            .I(n2018));
    Odrv4 I__2276 (
            .O(N__22907),
            .I(n2018));
    InMux I__2275 (
            .O(N__22900),
            .I(N__22897));
    LocalMux I__2274 (
            .O(N__22897),
            .I(n1988));
    CascadeMux I__2273 (
            .O(N__22894),
            .I(N__22891));
    InMux I__2272 (
            .O(N__22891),
            .I(N__22886));
    CascadeMux I__2271 (
            .O(N__22890),
            .I(N__22883));
    InMux I__2270 (
            .O(N__22889),
            .I(N__22880));
    LocalMux I__2269 (
            .O(N__22886),
            .I(N__22877));
    InMux I__2268 (
            .O(N__22883),
            .I(N__22874));
    LocalMux I__2267 (
            .O(N__22880),
            .I(n2020));
    Odrv4 I__2266 (
            .O(N__22877),
            .I(n2020));
    LocalMux I__2265 (
            .O(N__22874),
            .I(n2020));
    CascadeMux I__2264 (
            .O(N__22867),
            .I(N__22864));
    InMux I__2263 (
            .O(N__22864),
            .I(N__22861));
    LocalMux I__2262 (
            .O(N__22861),
            .I(n1987));
    InMux I__2261 (
            .O(N__22858),
            .I(N__22855));
    LocalMux I__2260 (
            .O(N__22855),
            .I(n1991));
    InMux I__2259 (
            .O(N__22852),
            .I(N__22849));
    LocalMux I__2258 (
            .O(N__22849),
            .I(N__22846));
    Span4Mux_h I__2257 (
            .O(N__22846),
            .I(N__22843));
    Odrv4 I__2256 (
            .O(N__22843),
            .I(n2098));
    CascadeMux I__2255 (
            .O(N__22840),
            .I(N__22837));
    InMux I__2254 (
            .O(N__22837),
            .I(N__22834));
    LocalMux I__2253 (
            .O(N__22834),
            .I(n2392));
    InMux I__2252 (
            .O(N__22831),
            .I(N__22828));
    LocalMux I__2251 (
            .O(N__22828),
            .I(N__22825));
    Odrv4 I__2250 (
            .O(N__22825),
            .I(n2096));
    CascadeMux I__2249 (
            .O(N__22822),
            .I(N__22819));
    InMux I__2248 (
            .O(N__22819),
            .I(N__22816));
    LocalMux I__2247 (
            .O(N__22816),
            .I(N__22813));
    Span4Mux_h I__2246 (
            .O(N__22813),
            .I(N__22810));
    Odrv4 I__2245 (
            .O(N__22810),
            .I(n2197));
    InMux I__2244 (
            .O(N__22807),
            .I(N__22804));
    LocalMux I__2243 (
            .O(N__22804),
            .I(n1996));
    CascadeMux I__2242 (
            .O(N__22801),
            .I(N__22798));
    InMux I__2241 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__2240 (
            .O(N__22795),
            .I(N__22792));
    Span4Mux_h I__2239 (
            .O(N__22792),
            .I(N__22789));
    Odrv4 I__2238 (
            .O(N__22789),
            .I(n2196));
    InMux I__2237 (
            .O(N__22786),
            .I(N__22783));
    LocalMux I__2236 (
            .O(N__22783),
            .I(N__22780));
    Span4Mux_v I__2235 (
            .O(N__22780),
            .I(N__22777));
    Odrv4 I__2234 (
            .O(N__22777),
            .I(n2201));
    InMux I__2233 (
            .O(N__22774),
            .I(N__22771));
    LocalMux I__2232 (
            .O(N__22771),
            .I(n14160));
    InMux I__2231 (
            .O(N__22768),
            .I(N__22765));
    LocalMux I__2230 (
            .O(N__22765),
            .I(N__22762));
    Span4Mux_h I__2229 (
            .O(N__22762),
            .I(N__22759));
    Odrv4 I__2228 (
            .O(N__22759),
            .I(n2186));
    InMux I__2227 (
            .O(N__22756),
            .I(n12308));
    InMux I__2226 (
            .O(N__22753),
            .I(n12309));
    InMux I__2225 (
            .O(N__22750),
            .I(N__22747));
    LocalMux I__2224 (
            .O(N__22747),
            .I(n2386));
    InMux I__2223 (
            .O(N__22744),
            .I(n12310));
    InMux I__2222 (
            .O(N__22741),
            .I(bfn_3_19_0_));
    InMux I__2221 (
            .O(N__22738),
            .I(n12312));
    InMux I__2220 (
            .O(N__22735),
            .I(n12313));
    InMux I__2219 (
            .O(N__22732),
            .I(n12314));
    InMux I__2218 (
            .O(N__22729),
            .I(n12315));
    InMux I__2217 (
            .O(N__22726),
            .I(n12316));
    InMux I__2216 (
            .O(N__22723),
            .I(n12299));
    InMux I__2215 (
            .O(N__22720),
            .I(n12300));
    InMux I__2214 (
            .O(N__22717),
            .I(n12301));
    InMux I__2213 (
            .O(N__22714),
            .I(n12302));
    InMux I__2212 (
            .O(N__22711),
            .I(bfn_3_18_0_));
    InMux I__2211 (
            .O(N__22708),
            .I(n12304));
    InMux I__2210 (
            .O(N__22705),
            .I(n12305));
    InMux I__2209 (
            .O(N__22702),
            .I(n12306));
    InMux I__2208 (
            .O(N__22699),
            .I(n12307));
    InMux I__2207 (
            .O(N__22696),
            .I(n12739));
    InMux I__2206 (
            .O(N__22693),
            .I(bfn_2_32_0_));
    InMux I__2205 (
            .O(N__22690),
            .I(n12741));
    InMux I__2204 (
            .O(N__22687),
            .I(N__22683));
    InMux I__2203 (
            .O(N__22686),
            .I(N__22680));
    LocalMux I__2202 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__2201 (
            .O(N__22680),
            .I(\debounce.cnt_reg_4 ));
    Odrv4 I__2200 (
            .O(N__22677),
            .I(\debounce.cnt_reg_4 ));
    InMux I__2199 (
            .O(N__22672),
            .I(N__22668));
    InMux I__2198 (
            .O(N__22671),
            .I(N__22665));
    LocalMux I__2197 (
            .O(N__22668),
            .I(N__22662));
    LocalMux I__2196 (
            .O(N__22665),
            .I(\debounce.cnt_reg_6 ));
    Odrv4 I__2195 (
            .O(N__22662),
            .I(\debounce.cnt_reg_6 ));
    CascadeMux I__2194 (
            .O(N__22657),
            .I(N__22654));
    InMux I__2193 (
            .O(N__22654),
            .I(N__22651));
    LocalMux I__2192 (
            .O(N__22651),
            .I(N__22647));
    InMux I__2191 (
            .O(N__22650),
            .I(N__22644));
    Span4Mux_s1_v I__2190 (
            .O(N__22647),
            .I(N__22641));
    LocalMux I__2189 (
            .O(N__22644),
            .I(\debounce.cnt_reg_0 ));
    Odrv4 I__2188 (
            .O(N__22641),
            .I(\debounce.cnt_reg_0 ));
    InMux I__2187 (
            .O(N__22636),
            .I(N__22632));
    InMux I__2186 (
            .O(N__22635),
            .I(N__22629));
    LocalMux I__2185 (
            .O(N__22632),
            .I(N__22626));
    LocalMux I__2184 (
            .O(N__22629),
            .I(\debounce.cnt_reg_7 ));
    Odrv4 I__2183 (
            .O(N__22626),
            .I(\debounce.cnt_reg_7 ));
    InMux I__2182 (
            .O(N__22621),
            .I(N__22618));
    LocalMux I__2181 (
            .O(N__22618),
            .I(\debounce.n13 ));
    InMux I__2180 (
            .O(N__22615),
            .I(bfn_3_17_0_));
    InMux I__2179 (
            .O(N__22612),
            .I(n12296));
    InMux I__2178 (
            .O(N__22609),
            .I(n12297));
    InMux I__2177 (
            .O(N__22606),
            .I(N__22603));
    LocalMux I__2176 (
            .O(N__22603),
            .I(n2398));
    InMux I__2175 (
            .O(N__22600),
            .I(n12298));
    InMux I__2174 (
            .O(N__22597),
            .I(N__22594));
    LocalMux I__2173 (
            .O(N__22594),
            .I(n11_adj_663));
    InMux I__2172 (
            .O(N__22591),
            .I(n12731));
    InMux I__2171 (
            .O(N__22588),
            .I(N__22585));
    LocalMux I__2170 (
            .O(N__22585),
            .I(n10_adj_662));
    InMux I__2169 (
            .O(N__22582),
            .I(bfn_2_31_0_));
    InMux I__2168 (
            .O(N__22579),
            .I(N__22576));
    LocalMux I__2167 (
            .O(N__22576),
            .I(n9_adj_661));
    InMux I__2166 (
            .O(N__22573),
            .I(n12733));
    InMux I__2165 (
            .O(N__22570),
            .I(N__22567));
    LocalMux I__2164 (
            .O(N__22567),
            .I(n8_adj_660));
    InMux I__2163 (
            .O(N__22564),
            .I(n12734));
    InMux I__2162 (
            .O(N__22561),
            .I(N__22558));
    LocalMux I__2161 (
            .O(N__22558),
            .I(n7_adj_659));
    InMux I__2160 (
            .O(N__22555),
            .I(n12735));
    InMux I__2159 (
            .O(N__22552),
            .I(N__22549));
    LocalMux I__2158 (
            .O(N__22549),
            .I(n6_adj_658));
    InMux I__2157 (
            .O(N__22546),
            .I(n12736));
    InMux I__2156 (
            .O(N__22543),
            .I(n12737));
    InMux I__2155 (
            .O(N__22540),
            .I(n12738));
    InMux I__2154 (
            .O(N__22537),
            .I(N__22534));
    LocalMux I__2153 (
            .O(N__22534),
            .I(n20_adj_672));
    InMux I__2152 (
            .O(N__22531),
            .I(n12722));
    InMux I__2151 (
            .O(N__22528),
            .I(N__22525));
    LocalMux I__2150 (
            .O(N__22525),
            .I(n19_adj_671));
    InMux I__2149 (
            .O(N__22522),
            .I(n12723));
    InMux I__2148 (
            .O(N__22519),
            .I(N__22516));
    LocalMux I__2147 (
            .O(N__22516),
            .I(n18_adj_670));
    InMux I__2146 (
            .O(N__22513),
            .I(bfn_2_30_0_));
    InMux I__2145 (
            .O(N__22510),
            .I(N__22507));
    LocalMux I__2144 (
            .O(N__22507),
            .I(n17_adj_669));
    InMux I__2143 (
            .O(N__22504),
            .I(n12725));
    InMux I__2142 (
            .O(N__22501),
            .I(N__22498));
    LocalMux I__2141 (
            .O(N__22498),
            .I(n16_adj_668));
    InMux I__2140 (
            .O(N__22495),
            .I(n12726));
    InMux I__2139 (
            .O(N__22492),
            .I(N__22489));
    LocalMux I__2138 (
            .O(N__22489),
            .I(n15_adj_667));
    InMux I__2137 (
            .O(N__22486),
            .I(n12727));
    InMux I__2136 (
            .O(N__22483),
            .I(N__22480));
    LocalMux I__2135 (
            .O(N__22480),
            .I(n14_adj_666));
    InMux I__2134 (
            .O(N__22477),
            .I(n12728));
    InMux I__2133 (
            .O(N__22474),
            .I(N__22471));
    LocalMux I__2132 (
            .O(N__22471),
            .I(n13_adj_665));
    InMux I__2131 (
            .O(N__22468),
            .I(n12729));
    InMux I__2130 (
            .O(N__22465),
            .I(N__22462));
    LocalMux I__2129 (
            .O(N__22462),
            .I(n12_adj_664));
    InMux I__2128 (
            .O(N__22459),
            .I(n12730));
    InMux I__2127 (
            .O(N__22456),
            .I(N__22453));
    LocalMux I__2126 (
            .O(N__22453),
            .I(n1491));
    InMux I__2125 (
            .O(N__22450),
            .I(N__22447));
    LocalMux I__2124 (
            .O(N__22447),
            .I(n26_adj_678));
    InMux I__2123 (
            .O(N__22444),
            .I(bfn_2_29_0_));
    InMux I__2122 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__2121 (
            .O(N__22438),
            .I(n25_adj_677));
    InMux I__2120 (
            .O(N__22435),
            .I(n12717));
    InMux I__2119 (
            .O(N__22432),
            .I(N__22429));
    LocalMux I__2118 (
            .O(N__22429),
            .I(n24_adj_676));
    InMux I__2117 (
            .O(N__22426),
            .I(n12718));
    InMux I__2116 (
            .O(N__22423),
            .I(N__22420));
    LocalMux I__2115 (
            .O(N__22420),
            .I(n23_adj_675));
    InMux I__2114 (
            .O(N__22417),
            .I(n12719));
    InMux I__2113 (
            .O(N__22414),
            .I(N__22411));
    LocalMux I__2112 (
            .O(N__22411),
            .I(n22_adj_674));
    InMux I__2111 (
            .O(N__22408),
            .I(n12720));
    InMux I__2110 (
            .O(N__22405),
            .I(N__22402));
    LocalMux I__2109 (
            .O(N__22402),
            .I(n21_adj_673));
    InMux I__2108 (
            .O(N__22399),
            .I(n12721));
    InMux I__2107 (
            .O(N__22396),
            .I(n12154));
    InMux I__2106 (
            .O(N__22393),
            .I(n12155));
    InMux I__2105 (
            .O(N__22390),
            .I(n12156));
    InMux I__2104 (
            .O(N__22387),
            .I(n12157));
    InMux I__2103 (
            .O(N__22384),
            .I(n12158));
    InMux I__2102 (
            .O(N__22381),
            .I(bfn_2_28_0_));
    InMux I__2101 (
            .O(N__22378),
            .I(n12160));
    InMux I__2100 (
            .O(N__22375),
            .I(n12161));
    InMux I__2099 (
            .O(N__22372),
            .I(n12162));
    InMux I__2098 (
            .O(N__22369),
            .I(n12163));
    CascadeMux I__2097 (
            .O(N__22366),
            .I(n13986_cascade_));
    CascadeMux I__2096 (
            .O(N__22363),
            .I(n1554_cascade_));
    CascadeMux I__2095 (
            .O(N__22360),
            .I(N__22356));
    CascadeMux I__2094 (
            .O(N__22359),
            .I(N__22352));
    InMux I__2093 (
            .O(N__22356),
            .I(N__22349));
    InMux I__2092 (
            .O(N__22355),
            .I(N__22344));
    InMux I__2091 (
            .O(N__22352),
            .I(N__22344));
    LocalMux I__2090 (
            .O(N__22349),
            .I(n1629));
    LocalMux I__2089 (
            .O(N__22344),
            .I(n1629));
    CascadeMux I__2088 (
            .O(N__22339),
            .I(N__22336));
    InMux I__2087 (
            .O(N__22336),
            .I(N__22331));
    InMux I__2086 (
            .O(N__22335),
            .I(N__22326));
    InMux I__2085 (
            .O(N__22334),
            .I(N__22326));
    LocalMux I__2084 (
            .O(N__22331),
            .I(n1631));
    LocalMux I__2083 (
            .O(N__22326),
            .I(n1631));
    InMux I__2082 (
            .O(N__22321),
            .I(bfn_2_27_0_));
    InMux I__2081 (
            .O(N__22318),
            .I(n12152));
    InMux I__2080 (
            .O(N__22315),
            .I(n12153));
    InMux I__2079 (
            .O(N__22312),
            .I(N__22309));
    LocalMux I__2078 (
            .O(N__22309),
            .I(n1698));
    CascadeMux I__2077 (
            .O(N__22306),
            .I(N__22303));
    InMux I__2076 (
            .O(N__22303),
            .I(N__22300));
    LocalMux I__2075 (
            .O(N__22300),
            .I(n1696));
    CascadeMux I__2074 (
            .O(N__22297),
            .I(n1728_cascade_));
    InMux I__2073 (
            .O(N__22294),
            .I(N__22291));
    LocalMux I__2072 (
            .O(N__22291),
            .I(n1695));
    CascadeMux I__2071 (
            .O(N__22288),
            .I(N__22285));
    InMux I__2070 (
            .O(N__22285),
            .I(N__22282));
    LocalMux I__2069 (
            .O(N__22282),
            .I(n1694));
    InMux I__2068 (
            .O(N__22279),
            .I(N__22276));
    LocalMux I__2067 (
            .O(N__22276),
            .I(N__22273));
    Span4Mux_h I__2066 (
            .O(N__22273),
            .I(N__22270));
    Odrv4 I__2065 (
            .O(N__22270),
            .I(n1689));
    CascadeMux I__2064 (
            .O(N__22267),
            .I(N__22264));
    InMux I__2063 (
            .O(N__22264),
            .I(N__22260));
    CascadeMux I__2062 (
            .O(N__22263),
            .I(N__22257));
    LocalMux I__2061 (
            .O(N__22260),
            .I(N__22253));
    InMux I__2060 (
            .O(N__22257),
            .I(N__22250));
    InMux I__2059 (
            .O(N__22256),
            .I(N__22247));
    Odrv12 I__2058 (
            .O(N__22253),
            .I(n1630));
    LocalMux I__2057 (
            .O(N__22250),
            .I(n1630));
    LocalMux I__2056 (
            .O(N__22247),
            .I(n1630));
    CascadeMux I__2055 (
            .O(N__22240),
            .I(N__22237));
    InMux I__2054 (
            .O(N__22237),
            .I(N__22234));
    LocalMux I__2053 (
            .O(N__22234),
            .I(N__22231));
    Odrv4 I__2052 (
            .O(N__22231),
            .I(n1700));
    InMux I__2051 (
            .O(N__22228),
            .I(N__22225));
    LocalMux I__2050 (
            .O(N__22225),
            .I(N__22222));
    Odrv4 I__2049 (
            .O(N__22222),
            .I(n1699));
    CascadeMux I__2048 (
            .O(N__22219),
            .I(n1731_cascade_));
    InMux I__2047 (
            .O(N__22216),
            .I(N__22213));
    LocalMux I__2046 (
            .O(N__22213),
            .I(N__22210));
    Odrv4 I__2045 (
            .O(N__22210),
            .I(n1697));
    CascadeMux I__2044 (
            .O(N__22207),
            .I(n1729_cascade_));
    InMux I__2043 (
            .O(N__22204),
            .I(N__22201));
    LocalMux I__2042 (
            .O(N__22201),
            .I(N__22198));
    Odrv4 I__2041 (
            .O(N__22198),
            .I(n1701));
    CascadeMux I__2040 (
            .O(N__22195),
            .I(n1733_cascade_));
    CascadeMux I__2039 (
            .O(N__22192),
            .I(N__22189));
    InMux I__2038 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__2037 (
            .O(N__22186),
            .I(n1886));
    InMux I__2036 (
            .O(N__22183),
            .I(n12233));
    InMux I__2035 (
            .O(N__22180),
            .I(n12234));
    InMux I__2034 (
            .O(N__22177),
            .I(n12235));
    InMux I__2033 (
            .O(N__22174),
            .I(n12236));
    InMux I__2032 (
            .O(N__22171),
            .I(bfn_2_23_0_));
    InMux I__2031 (
            .O(N__22168),
            .I(n12238));
    CascadeMux I__2030 (
            .O(N__22165),
            .I(N__22162));
    InMux I__2029 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__2028 (
            .O(N__22159),
            .I(N__22155));
    InMux I__2027 (
            .O(N__22158),
            .I(N__22152));
    Span4Mux_s2_h I__2026 (
            .O(N__22155),
            .I(N__22149));
    LocalMux I__2025 (
            .O(N__22152),
            .I(n2016));
    Odrv4 I__2024 (
            .O(N__22149),
            .I(n2016));
    InMux I__2023 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__2022 (
            .O(N__22141),
            .I(n1888));
    InMux I__2021 (
            .O(N__22138),
            .I(N__22135));
    LocalMux I__2020 (
            .O(N__22135),
            .I(n1985));
    CascadeMux I__2019 (
            .O(N__22132),
            .I(N__22129));
    InMux I__2018 (
            .O(N__22129),
            .I(N__22126));
    LocalMux I__2017 (
            .O(N__22126),
            .I(N__22122));
    InMux I__2016 (
            .O(N__22125),
            .I(N__22118));
    Span4Mux_v I__2015 (
            .O(N__22122),
            .I(N__22115));
    InMux I__2014 (
            .O(N__22121),
            .I(N__22112));
    LocalMux I__2013 (
            .O(N__22118),
            .I(N__22109));
    Odrv4 I__2012 (
            .O(N__22115),
            .I(n2017));
    LocalMux I__2011 (
            .O(N__22112),
            .I(n2017));
    Odrv12 I__2010 (
            .O(N__22109),
            .I(n2017));
    InMux I__2009 (
            .O(N__22102),
            .I(n12223));
    InMux I__2008 (
            .O(N__22099),
            .I(n12224));
    InMux I__2007 (
            .O(N__22096),
            .I(n12225));
    InMux I__2006 (
            .O(N__22093),
            .I(n12226));
    InMux I__2005 (
            .O(N__22090),
            .I(n12227));
    InMux I__2004 (
            .O(N__22087),
            .I(n12228));
    InMux I__2003 (
            .O(N__22084),
            .I(bfn_2_22_0_));
    InMux I__2002 (
            .O(N__22081),
            .I(n12230));
    InMux I__2001 (
            .O(N__22078),
            .I(n12231));
    InMux I__2000 (
            .O(N__22075),
            .I(n12232));
    InMux I__1999 (
            .O(N__22072),
            .I(N__22069));
    LocalMux I__1998 (
            .O(N__22069),
            .I(N__22066));
    Odrv4 I__1997 (
            .O(N__22066),
            .I(n2084));
    CascadeMux I__1996 (
            .O(N__22063),
            .I(N__22060));
    InMux I__1995 (
            .O(N__22060),
            .I(N__22056));
    InMux I__1994 (
            .O(N__22059),
            .I(N__22053));
    LocalMux I__1993 (
            .O(N__22056),
            .I(n2116));
    LocalMux I__1992 (
            .O(N__22053),
            .I(n2116));
    CascadeMux I__1991 (
            .O(N__22048),
            .I(N__22045));
    InMux I__1990 (
            .O(N__22045),
            .I(N__22041));
    InMux I__1989 (
            .O(N__22044),
            .I(N__22038));
    LocalMux I__1988 (
            .O(N__22041),
            .I(N__22033));
    LocalMux I__1987 (
            .O(N__22038),
            .I(N__22033));
    Odrv4 I__1986 (
            .O(N__22033),
            .I(n2115));
    CascadeMux I__1985 (
            .O(N__22030),
            .I(n2116_cascade_));
    CascadeMux I__1984 (
            .O(N__22027),
            .I(n2148_cascade_));
    InMux I__1983 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__1982 (
            .O(N__22021),
            .I(N__22018));
    Odrv4 I__1981 (
            .O(N__22018),
            .I(n2195));
    InMux I__1980 (
            .O(N__22015),
            .I(N__22012));
    LocalMux I__1979 (
            .O(N__22012),
            .I(n2087));
    InMux I__1978 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__1977 (
            .O(N__22006),
            .I(n2093));
    InMux I__1976 (
            .O(N__22003),
            .I(N__22000));
    LocalMux I__1975 (
            .O(N__22000),
            .I(N__21997));
    Span4Mux_v I__1974 (
            .O(N__21997),
            .I(N__21994));
    Odrv4 I__1973 (
            .O(N__21994),
            .I(n2085));
    InMux I__1972 (
            .O(N__21991),
            .I(N__21986));
    InMux I__1971 (
            .O(N__21990),
            .I(N__21981));
    InMux I__1970 (
            .O(N__21989),
            .I(N__21981));
    LocalMux I__1969 (
            .O(N__21986),
            .I(n2117));
    LocalMux I__1968 (
            .O(N__21981),
            .I(n2117));
    InMux I__1967 (
            .O(N__21976),
            .I(bfn_2_21_0_));
    InMux I__1966 (
            .O(N__21973),
            .I(n12222));
    CascadeMux I__1965 (
            .O(N__21970),
            .I(n2331_cascade_));
    CascadeMux I__1964 (
            .O(N__21967),
            .I(N__21964));
    InMux I__1963 (
            .O(N__21964),
            .I(N__21961));
    LocalMux I__1962 (
            .O(N__21961),
            .I(N__21958));
    Odrv4 I__1961 (
            .O(N__21958),
            .I(n2089));
    InMux I__1960 (
            .O(N__21955),
            .I(N__21952));
    LocalMux I__1959 (
            .O(N__21952),
            .I(n2188));
    CascadeMux I__1958 (
            .O(N__21949),
            .I(n2121_cascade_));
    CascadeMux I__1957 (
            .O(N__21946),
            .I(n2220_cascade_));
    CascadeMux I__1956 (
            .O(N__21943),
            .I(n2319_cascade_));
    InMux I__1955 (
            .O(N__21940),
            .I(N__21937));
    LocalMux I__1954 (
            .O(N__21937),
            .I(n2097));
    CascadeMux I__1953 (
            .O(N__21934),
            .I(n2049_cascade_));
    InMux I__1952 (
            .O(N__21931),
            .I(N__21928));
    LocalMux I__1951 (
            .O(N__21928),
            .I(n2183));
    InMux I__1950 (
            .O(N__21925),
            .I(N__21922));
    LocalMux I__1949 (
            .O(N__21922),
            .I(n2184));
    InMux I__1948 (
            .O(N__21919),
            .I(N__21915));
    InMux I__1947 (
            .O(N__21918),
            .I(N__21912));
    LocalMux I__1946 (
            .O(N__21915),
            .I(N__21909));
    LocalMux I__1945 (
            .O(N__21912),
            .I(\debounce.cnt_reg_3 ));
    Odrv4 I__1944 (
            .O(N__21909),
            .I(\debounce.cnt_reg_3 ));
    InMux I__1943 (
            .O(N__21904),
            .I(N__21900));
    InMux I__1942 (
            .O(N__21903),
            .I(N__21897));
    LocalMux I__1941 (
            .O(N__21900),
            .I(N__21894));
    LocalMux I__1940 (
            .O(N__21897),
            .I(\debounce.cnt_reg_9 ));
    Odrv4 I__1939 (
            .O(N__21894),
            .I(\debounce.cnt_reg_9 ));
    CascadeMux I__1938 (
            .O(N__21889),
            .I(N__21886));
    InMux I__1937 (
            .O(N__21886),
            .I(N__21882));
    InMux I__1936 (
            .O(N__21885),
            .I(N__21879));
    LocalMux I__1935 (
            .O(N__21882),
            .I(N__21876));
    LocalMux I__1934 (
            .O(N__21879),
            .I(\debounce.cnt_reg_5 ));
    Odrv4 I__1933 (
            .O(N__21876),
            .I(\debounce.cnt_reg_5 ));
    InMux I__1932 (
            .O(N__21871),
            .I(N__21867));
    InMux I__1931 (
            .O(N__21870),
            .I(N__21864));
    LocalMux I__1930 (
            .O(N__21867),
            .I(N__21861));
    LocalMux I__1929 (
            .O(N__21864),
            .I(\debounce.cnt_reg_8 ));
    Odrv4 I__1928 (
            .O(N__21861),
            .I(\debounce.cnt_reg_8 ));
    InMux I__1927 (
            .O(N__21856),
            .I(N__21852));
    InMux I__1926 (
            .O(N__21855),
            .I(N__21849));
    LocalMux I__1925 (
            .O(N__21852),
            .I(N__21846));
    LocalMux I__1924 (
            .O(N__21849),
            .I(\debounce.cnt_reg_1 ));
    Odrv12 I__1923 (
            .O(N__21846),
            .I(\debounce.cnt_reg_1 ));
    InMux I__1922 (
            .O(N__21841),
            .I(N__21837));
    InMux I__1921 (
            .O(N__21840),
            .I(N__21834));
    LocalMux I__1920 (
            .O(N__21837),
            .I(N__21831));
    LocalMux I__1919 (
            .O(N__21834),
            .I(\debounce.cnt_reg_2 ));
    Odrv4 I__1918 (
            .O(N__21831),
            .I(\debounce.cnt_reg_2 ));
    CascadeMux I__1917 (
            .O(N__21826),
            .I(\debounce.n14472_cascade_ ));
    InMux I__1916 (
            .O(N__21823),
            .I(N__21820));
    LocalMux I__1915 (
            .O(N__21820),
            .I(N__21817));
    Odrv4 I__1914 (
            .O(N__21817),
            .I(n2095));
    InMux I__1913 (
            .O(N__21814),
            .I(N__21811));
    LocalMux I__1912 (
            .O(N__21811),
            .I(N__21808));
    Span4Mux_v I__1911 (
            .O(N__21808),
            .I(N__21805));
    Odrv4 I__1910 (
            .O(N__21805),
            .I(n2094));
    InMux I__1909 (
            .O(N__21802),
            .I(N__21799));
    LocalMux I__1908 (
            .O(N__21799),
            .I(N__21796));
    Odrv4 I__1907 (
            .O(N__21796),
            .I(n2101));
    InMux I__1906 (
            .O(N__21793),
            .I(N__21790));
    LocalMux I__1905 (
            .O(N__21790),
            .I(n2200));
    CascadeMux I__1904 (
            .O(N__21787),
            .I(n2133_cascade_));
    CascadeMux I__1903 (
            .O(N__21784),
            .I(n2232_cascade_));
    InMux I__1902 (
            .O(N__21781),
            .I(n12122));
    InMux I__1901 (
            .O(N__21778),
            .I(n12123));
    InMux I__1900 (
            .O(N__21775),
            .I(n12124));
    InMux I__1899 (
            .O(N__21772),
            .I(n12125));
    InMux I__1898 (
            .O(N__21769),
            .I(n12126));
    InMux I__1897 (
            .O(N__21766),
            .I(n12127));
    InMux I__1896 (
            .O(N__21763),
            .I(n12128));
    InMux I__1895 (
            .O(N__21760),
            .I(bfn_1_32_0_));
    InMux I__1894 (
            .O(N__21757),
            .I(n12130));
    InMux I__1893 (
            .O(N__21754),
            .I(\debounce.n12655 ));
    InMux I__1892 (
            .O(N__21751),
            .I(\debounce.n12656 ));
    InMux I__1891 (
            .O(N__21748),
            .I(\debounce.n12657 ));
    InMux I__1890 (
            .O(N__21745),
            .I(\debounce.n12658 ));
    InMux I__1889 (
            .O(N__21742),
            .I(\debounce.n12659 ));
    InMux I__1888 (
            .O(N__21739),
            .I(\debounce.n12660 ));
    InMux I__1887 (
            .O(N__21736),
            .I(bfn_1_30_0_));
    InMux I__1886 (
            .O(N__21733),
            .I(\debounce.n12662 ));
    InMux I__1885 (
            .O(N__21730),
            .I(bfn_1_31_0_));
    InMux I__1884 (
            .O(N__21727),
            .I(n12188));
    InMux I__1883 (
            .O(N__21724),
            .I(n12189));
    InMux I__1882 (
            .O(N__21721),
            .I(n12190));
    CascadeMux I__1881 (
            .O(N__21718),
            .I(n1427_cascade_));
    CascadeMux I__1880 (
            .O(N__21715),
            .I(n1430_cascade_));
    InMux I__1879 (
            .O(N__21712),
            .I(N__21709));
    LocalMux I__1878 (
            .O(N__21709),
            .I(n11638));
    InMux I__1877 (
            .O(N__21706),
            .I(bfn_1_29_0_));
    InMux I__1876 (
            .O(N__21703),
            .I(\debounce.n12654 ));
    InMux I__1875 (
            .O(N__21700),
            .I(n12179));
    InMux I__1874 (
            .O(N__21697),
            .I(n12180));
    InMux I__1873 (
            .O(N__21694),
            .I(n12181));
    InMux I__1872 (
            .O(N__21691),
            .I(n12182));
    InMux I__1871 (
            .O(N__21688),
            .I(n12183));
    InMux I__1870 (
            .O(N__21685),
            .I(bfn_1_27_0_));
    InMux I__1869 (
            .O(N__21682),
            .I(n12185));
    InMux I__1868 (
            .O(N__21679),
            .I(n12186));
    InMux I__1867 (
            .O(N__21676),
            .I(n12187));
    InMux I__1866 (
            .O(N__21673),
            .I(n12216));
    InMux I__1865 (
            .O(N__21670),
            .I(n12217));
    InMux I__1864 (
            .O(N__21667),
            .I(n12218));
    InMux I__1863 (
            .O(N__21664),
            .I(n12219));
    InMux I__1862 (
            .O(N__21661),
            .I(n12220));
    InMux I__1861 (
            .O(N__21658),
            .I(bfn_1_25_0_));
    InMux I__1860 (
            .O(N__21655),
            .I(bfn_1_26_0_));
    InMux I__1859 (
            .O(N__21652),
            .I(n12177));
    InMux I__1858 (
            .O(N__21649),
            .I(n12178));
    InMux I__1857 (
            .O(N__21646),
            .I(n12207));
    InMux I__1856 (
            .O(N__21643),
            .I(n12208));
    InMux I__1855 (
            .O(N__21640),
            .I(n12209));
    InMux I__1854 (
            .O(N__21637),
            .I(n12210));
    InMux I__1853 (
            .O(N__21634),
            .I(n12211));
    InMux I__1852 (
            .O(N__21631),
            .I(n12212));
    InMux I__1851 (
            .O(N__21628),
            .I(bfn_1_24_0_));
    InMux I__1850 (
            .O(N__21625),
            .I(n12214));
    InMux I__1849 (
            .O(N__21622),
            .I(n12215));
    InMux I__1848 (
            .O(N__21619),
            .I(n12250));
    InMux I__1847 (
            .O(N__21616),
            .I(n12251));
    InMux I__1846 (
            .O(N__21613),
            .I(n12252));
    InMux I__1845 (
            .O(N__21610),
            .I(n12253));
    InMux I__1844 (
            .O(N__21607),
            .I(bfn_1_22_0_));
    InMux I__1843 (
            .O(N__21604),
            .I(n12255));
    InMux I__1842 (
            .O(N__21601),
            .I(n12256));
    InMux I__1841 (
            .O(N__21598),
            .I(bfn_1_23_0_));
    InMux I__1840 (
            .O(N__21595),
            .I(n12206));
    InMux I__1839 (
            .O(N__21592),
            .I(n12241));
    InMux I__1838 (
            .O(N__21589),
            .I(n12242));
    InMux I__1837 (
            .O(N__21586),
            .I(n12243));
    InMux I__1836 (
            .O(N__21583),
            .I(n12244));
    InMux I__1835 (
            .O(N__21580),
            .I(n12245));
    InMux I__1834 (
            .O(N__21577),
            .I(bfn_1_21_0_));
    InMux I__1833 (
            .O(N__21574),
            .I(n12247));
    InMux I__1832 (
            .O(N__21571),
            .I(n12248));
    InMux I__1831 (
            .O(N__21568),
            .I(n12249));
    InMux I__1830 (
            .O(N__21565),
            .I(n12271));
    InMux I__1829 (
            .O(N__21562),
            .I(bfn_1_19_0_));
    InMux I__1828 (
            .O(N__21559),
            .I(n12273));
    InMux I__1827 (
            .O(N__21556),
            .I(n12274));
    InMux I__1826 (
            .O(N__21553),
            .I(n12275));
    InMux I__1825 (
            .O(N__21550),
            .I(bfn_1_20_0_));
    InMux I__1824 (
            .O(N__21547),
            .I(n12239));
    InMux I__1823 (
            .O(N__21544),
            .I(n12240));
    InMux I__1822 (
            .O(N__21541),
            .I(n12262));
    InMux I__1821 (
            .O(N__21538),
            .I(n12263));
    InMux I__1820 (
            .O(N__21535),
            .I(bfn_1_18_0_));
    InMux I__1819 (
            .O(N__21532),
            .I(n12265));
    InMux I__1818 (
            .O(N__21529),
            .I(n12266));
    InMux I__1817 (
            .O(N__21526),
            .I(n12267));
    InMux I__1816 (
            .O(N__21523),
            .I(n12268));
    InMux I__1815 (
            .O(N__21520),
            .I(n12269));
    InMux I__1814 (
            .O(N__21517),
            .I(n12270));
    InMux I__1813 (
            .O(N__21514),
            .I(bfn_1_17_0_));
    InMux I__1812 (
            .O(N__21511),
            .I(n12257));
    InMux I__1811 (
            .O(N__21508),
            .I(n12258));
    InMux I__1810 (
            .O(N__21505),
            .I(n12259));
    InMux I__1809 (
            .O(N__21502),
            .I(n12260));
    InMux I__1808 (
            .O(N__21499),
            .I(n12261));
    IoInMux I__1807 (
            .O(N__21496),
            .I(N__21493));
    LocalMux I__1806 (
            .O(N__21493),
            .I(N__21490));
    IoSpan4Mux I__1805 (
            .O(N__21490),
            .I(N__21487));
    IoSpan4Mux I__1804 (
            .O(N__21487),
            .I(N__21484));
    IoSpan4Mux I__1803 (
            .O(N__21484),
            .I(N__21481));
    Odrv4 I__1802 (
            .O(N__21481),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(n12528),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(n12536),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(n12544),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_28_0_));
    defparam IN_MUX_bfv_13_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_29_0_ (
            .carryinitin(n12057),
            .carryinitout(bfn_13_29_0_));
    defparam IN_MUX_bfv_13_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_30_0_ (
            .carryinitin(n12065),
            .carryinitout(bfn_13_30_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(n12613),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(n12621),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(\quad_counter0.n12630 ),
            .carryinitout(bfn_6_24_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(\quad_counter0.n12638 ),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_6_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_26_0_ (
            .carryinitin(\quad_counter0.n12646 ),
            .carryinitout(bfn_6_26_0_));
    defparam IN_MUX_bfv_16_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_26_0_));
    defparam IN_MUX_bfv_16_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_27_0_ (
            .carryinitin(n12670),
            .carryinitout(bfn_16_27_0_));
    defparam IN_MUX_bfv_16_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_28_0_ (
            .carryinitin(n12678),
            .carryinitout(bfn_16_28_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(n12080),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(n12088),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(n12582),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(n12590),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(n12598),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_27_0_));
    defparam IN_MUX_bfv_2_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_28_0_ (
            .carryinitin(n12159),
            .carryinitout(bfn_2_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_3_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_30_0_ (
            .carryinitin(n12148),
            .carryinitout(bfn_3_30_0_));
    defparam IN_MUX_bfv_3_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_31_0_));
    defparam IN_MUX_bfv_3_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_32_0_ (
            .carryinitin(n12138),
            .carryinitout(bfn_3_32_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(n12129),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_6_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_31_0_));
    defparam IN_MUX_bfv_6_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_32_0_ (
            .carryinitin(n12121),
            .carryinitout(bfn_6_32_0_));
    defparam IN_MUX_bfv_7_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_30_0_));
    defparam IN_MUX_bfv_7_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_29_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(n12499),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(n12507),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(n12515),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(n12471),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(n12479),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(n12487),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(n12444),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(n12452),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(n12460),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(n12418),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(n12426),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(n12434),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(n12393),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(n12401),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(n12409),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(n12369),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(n12377),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(n12385),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(n12346),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(n12354),
            .carryinitout(bfn_6_16_0_));
    defparam IN_MUX_bfv_6_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_17_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(n12324),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_6_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_19_0_ (
            .carryinitin(n12332),
            .carryinitout(bfn_6_19_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(n12303),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(n12311),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(n12283),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(n12291),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(n12264),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(n12272),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(n12246),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(n12254),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(n12229),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(n12237),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(n12213),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(n12221),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_4_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_25_0_ (
            .carryinitin(n12198),
            .carryinitout(bfn_4_25_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_1_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_27_0_ (
            .carryinitin(n12184),
            .carryinitout(bfn_1_27_0_));
    defparam IN_MUX_bfv_4_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_26_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(n12171),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(\debounce.n12661 ),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(n12724),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_2_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_31_0_ (
            .carryinitin(n12732),
            .carryinitout(bfn_2_31_0_));
    defparam IN_MUX_bfv_2_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_32_0_ (
            .carryinitin(n12740),
            .carryinitout(bfn_2_32_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(n12559),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(n12567),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_5_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_28_0_));
    defparam IN_MUX_bfv_11_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_29_0_));
    defparam IN_MUX_bfv_11_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_30_0_ (
            .carryinitin(\PWM.n12693 ),
            .carryinitout(bfn_11_30_0_));
    defparam IN_MUX_bfv_11_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_31_0_ (
            .carryinitin(\PWM.n12701 ),
            .carryinitout(bfn_11_31_0_));
    defparam IN_MUX_bfv_11_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_32_0_ (
            .carryinitin(\PWM.n12709 ),
            .carryinitout(bfn_11_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21496),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_1_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_1_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_1_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_2_lut_LC_1_17_0 (
            .in0(_gnd_net_),
            .in1(N__27994),
            .in2(_gnd_net_),
            .in3(N__21514),
            .lcout(n2201),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(n12257),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_1_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_1_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_1_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_3_lut_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(N__53827),
            .in2(N__26793),
            .in3(N__21511),
            .lcout(n2200),
            .ltout(),
            .carryin(n12257),
            .carryout(n12258),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_1_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_1_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_1_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_4_lut_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26635),
            .in3(N__21508),
            .lcout(n2199),
            .ltout(),
            .carryin(n12258),
            .carryout(n12259),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_1_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_1_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_1_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_5_lut_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(N__53828),
            .in2(N__26710),
            .in3(N__21505),
            .lcout(n2198),
            .ltout(),
            .carryin(n12259),
            .carryout(n12260),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_1_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_1_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_1_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_6_lut_LC_1_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26743),
            .in3(N__21502),
            .lcout(n2197),
            .ltout(),
            .carryin(n12260),
            .carryout(n12261),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_1_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_1_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_1_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_7_lut_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26773),
            .in3(N__21499),
            .lcout(n2196),
            .ltout(),
            .carryin(n12261),
            .carryout(n12262),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_1_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_1_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_1_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_8_lut_LC_1_17_6 (
            .in0(_gnd_net_),
            .in1(N__53830),
            .in2(N__24568),
            .in3(N__21541),
            .lcout(n2195),
            .ltout(),
            .carryin(n12262),
            .carryout(n12263),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_1_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_1_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_1_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_9_lut_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(N__53829),
            .in2(N__29366),
            .in3(N__21538),
            .lcout(n2194),
            .ltout(),
            .carryin(n12263),
            .carryout(n12264),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_1_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_1_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_1_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_10_lut_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(N__53611),
            .in2(N__29177),
            .in3(N__21535),
            .lcout(n2193),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(n12265),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_1_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_1_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_1_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_11_lut_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(N__29501),
            .in2(N__53990),
            .in3(N__21532),
            .lcout(n2192),
            .ltout(),
            .carryin(n12265),
            .carryout(n12266),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_1_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_1_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_1_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_12_lut_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(N__53615),
            .in2(N__29581),
            .in3(N__21529),
            .lcout(n2191),
            .ltout(),
            .carryin(n12266),
            .carryout(n12267),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_1_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_1_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_1_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_13_lut_LC_1_18_3 (
            .in0(_gnd_net_),
            .in1(N__53620),
            .in2(N__27112),
            .in3(N__21526),
            .lcout(n2190),
            .ltout(),
            .carryin(n12267),
            .carryout(n12268),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_1_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_1_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_1_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_14_lut_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(N__53616),
            .in2(N__24592),
            .in3(N__21523),
            .lcout(n2189),
            .ltout(),
            .carryin(n12268),
            .carryout(n12269),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_1_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_1_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_1_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_15_lut_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(N__53621),
            .in2(N__27087),
            .in3(N__21520),
            .lcout(n2188),
            .ltout(),
            .carryin(n12269),
            .carryout(n12270),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_1_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_1_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_1_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_16_lut_LC_1_18_6 (
            .in0(_gnd_net_),
            .in1(N__27607),
            .in2(N__53992),
            .in3(N__21517),
            .lcout(n2187),
            .ltout(),
            .carryin(n12270),
            .carryout(n12271),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_1_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_1_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_1_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_17_lut_LC_1_18_7 (
            .in0(_gnd_net_),
            .in1(N__27057),
            .in2(N__53991),
            .in3(N__21565),
            .lcout(n2186),
            .ltout(),
            .carryin(n12271),
            .carryout(n12272),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_1_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_1_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_1_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_18_lut_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(N__29692),
            .in2(N__54920),
            .in3(N__21562),
            .lcout(n2185),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(n12273),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_1_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_1_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_19_lut_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(N__21991),
            .in2(N__54925),
            .in3(N__21559),
            .lcout(n2184),
            .ltout(),
            .carryin(n12273),
            .carryout(n12274),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_1_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_1_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_1_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_20_lut_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(N__22059),
            .in2(N__54921),
            .in3(N__21556),
            .lcout(n2183),
            .ltout(),
            .carryin(n12274),
            .carryout(n12275),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_1_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_1_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_1_19_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1436_21_lut_LC_1_19_3 (
            .in0(N__54517),
            .in1(N__36222),
            .in2(N__22048),
            .in3(N__21553),
            .lcout(n2214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12563_1_lut_LC_1_19_7.C_ON=1'b0;
    defparam i12563_1_lut_LC_1_19_7.SEQ_MODE=4'b0000;
    defparam i12563_1_lut_LC_1_19_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12563_1_lut_LC_1_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35994),
            .lcout(n15035),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_1_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_1_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_1_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_2_lut_LC_1_20_0 (
            .in0(_gnd_net_),
            .in1(N__27922),
            .in2(_gnd_net_),
            .in3(N__21550),
            .lcout(n2101),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(n12239),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_1_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_1_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_1_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_3_lut_LC_1_20_1 (
            .in0(_gnd_net_),
            .in1(N__54518),
            .in2(N__26671),
            .in3(N__21547),
            .lcout(n2100),
            .ltout(),
            .carryin(n12239),
            .carryout(n12240),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_1_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_1_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_1_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_4_lut_LC_1_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27181),
            .in3(N__21544),
            .lcout(n2099),
            .ltout(),
            .carryin(n12240),
            .carryout(n12241),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_1_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_1_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_1_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_5_lut_LC_1_20_3 (
            .in0(_gnd_net_),
            .in1(N__54519),
            .in2(N__24454),
            .in3(N__21592),
            .lcout(n2098),
            .ltout(),
            .carryin(n12241),
            .carryout(n12242),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_1_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_1_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_1_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_6_lut_LC_1_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24241),
            .in3(N__21589),
            .lcout(n2097),
            .ltout(),
            .carryin(n12242),
            .carryout(n12243),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_1_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_1_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_1_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_7_lut_LC_1_20_5 (
            .in0(_gnd_net_),
            .in1(N__24262),
            .in2(_gnd_net_),
            .in3(N__21586),
            .lcout(n2096),
            .ltout(),
            .carryin(n12243),
            .carryout(n12244),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_1_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_1_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_1_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_8_lut_LC_1_20_6 (
            .in0(_gnd_net_),
            .in1(N__54521),
            .in2(N__23034),
            .in3(N__21583),
            .lcout(n2095),
            .ltout(),
            .carryin(n12244),
            .carryout(n12245),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_1_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_1_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_1_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_9_lut_LC_1_20_7 (
            .in0(_gnd_net_),
            .in1(N__54520),
            .in2(N__24661),
            .in3(N__21580),
            .lcout(n2094),
            .ltout(),
            .carryin(n12245),
            .carryout(n12246),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_1_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_1_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_1_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_10_lut_LC_1_21_0 (
            .in0(_gnd_net_),
            .in1(N__54501),
            .in2(N__22981),
            .in3(N__21577),
            .lcout(n2093),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(n12247),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_1_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_1_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_1_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_11_lut_LC_1_21_1 (
            .in0(_gnd_net_),
            .in1(N__29626),
            .in2(N__54922),
            .in3(N__21574),
            .lcout(n2092),
            .ltout(),
            .carryin(n12247),
            .carryout(n12248),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_1_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_1_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_1_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_12_lut_LC_1_21_2 (
            .in0(_gnd_net_),
            .in1(N__54505),
            .in2(N__27139),
            .in3(N__21571),
            .lcout(n2091),
            .ltout(),
            .carryin(n12248),
            .carryout(n12249),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_1_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_1_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_1_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_13_lut_LC_1_21_3 (
            .in0(_gnd_net_),
            .in1(N__24628),
            .in2(N__54923),
            .in3(N__21568),
            .lcout(n2090),
            .ltout(),
            .carryin(n12249),
            .carryout(n12250),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_1_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_1_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_1_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_14_lut_LC_1_21_4 (
            .in0(_gnd_net_),
            .in1(N__54509),
            .in2(N__24165),
            .in3(N__21619),
            .lcout(n2089),
            .ltout(),
            .carryin(n12250),
            .carryout(n12251),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_1_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_1_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_1_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_15_lut_LC_1_21_5 (
            .in0(_gnd_net_),
            .in1(N__54531),
            .in2(N__27652),
            .in3(N__21616),
            .lcout(n2088),
            .ltout(),
            .carryin(n12251),
            .carryout(n12252),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_1_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_1_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_1_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_16_lut_LC_1_21_6 (
            .in0(_gnd_net_),
            .in1(N__54510),
            .in2(N__22894),
            .in3(N__21613),
            .lcout(n2087),
            .ltout(),
            .carryin(n12252),
            .carryout(n12253),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_1_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_1_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_1_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_17_lut_LC_1_21_7 (
            .in0(_gnd_net_),
            .in1(N__29712),
            .in2(N__54924),
            .in3(N__21610),
            .lcout(n2086),
            .ltout(),
            .carryin(n12253),
            .carryout(n12254),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_1_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_1_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_18_lut_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__22930),
            .in2(N__54934),
            .in3(N__21607),
            .lcout(n2085),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n12255),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_1_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_1_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_19_lut_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__22121),
            .in2(N__54935),
            .in3(N__21604),
            .lcout(n2084),
            .ltout(),
            .carryin(n12255),
            .carryout(n12256),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_1_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_1_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_1_22_2.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1369_20_lut_LC_1_22_2 (
            .in0(N__54535),
            .in1(N__22158),
            .in2(N__36072),
            .in3(N__21601),
            .lcout(n2115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_1_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_1_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_1_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_2_lut_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__32694),
            .in2(_gnd_net_),
            .in3(N__21598),
            .lcout(n1901),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(n12206),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_1_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_1_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_1_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_3_lut_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__54936),
            .in2(N__28024),
            .in3(N__21595),
            .lcout(n1900),
            .ltout(),
            .carryin(n12206),
            .carryout(n12207),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_1_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_1_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_1_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_4_lut_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27711),
            .in3(N__21646),
            .lcout(n1899),
            .ltout(),
            .carryin(n12207),
            .carryout(n12208),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_1_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_1_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_1_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_5_lut_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__54937),
            .in2(N__27685),
            .in3(N__21643),
            .lcout(n1898),
            .ltout(),
            .carryin(n12208),
            .carryout(n12209),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_1_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_1_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_1_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_6_lut_LC_1_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27272),
            .in3(N__21640),
            .lcout(n1897),
            .ltout(),
            .carryin(n12209),
            .carryout(n12210),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_1_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_1_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_1_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_7_lut_LC_1_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27244),
            .in3(N__21637),
            .lcout(n1896),
            .ltout(),
            .carryin(n12210),
            .carryout(n12211),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_1_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_1_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_1_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_8_lut_LC_1_23_6 (
            .in0(_gnd_net_),
            .in1(N__54939),
            .in2(N__27742),
            .in3(N__21634),
            .lcout(n1895),
            .ltout(),
            .carryin(n12211),
            .carryout(n12212),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_1_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_1_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_1_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_9_lut_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(N__54938),
            .in2(N__27834),
            .in3(N__21631),
            .lcout(n1894),
            .ltout(),
            .carryin(n12212),
            .carryout(n12213),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_1_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_1_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_1_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_10_lut_LC_1_24_0 (
            .in0(_gnd_net_),
            .in1(N__54940),
            .in2(N__27808),
            .in3(N__21628),
            .lcout(n1893),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(n12214),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_1_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_1_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_1_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_11_lut_LC_1_24_1 (
            .in0(_gnd_net_),
            .in1(N__54947),
            .in2(N__27858),
            .in3(N__21625),
            .lcout(n1892),
            .ltout(),
            .carryin(n12214),
            .carryout(n12215),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_1_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_1_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_1_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_12_lut_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__54941),
            .in2(N__27310),
            .in3(N__21622),
            .lcout(n1891),
            .ltout(),
            .carryin(n12215),
            .carryout(n12216),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_1_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_1_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_1_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_13_lut_LC_1_24_3 (
            .in0(_gnd_net_),
            .in1(N__27325),
            .in2(N__55134),
            .in3(N__21673),
            .lcout(n1890),
            .ltout(),
            .carryin(n12216),
            .carryout(n12217),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_1_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_1_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_1_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_14_lut_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__54945),
            .in2(N__27010),
            .in3(N__21670),
            .lcout(n1889),
            .ltout(),
            .carryin(n12217),
            .carryout(n12218),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_1_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_1_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_1_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_15_lut_LC_1_24_5 (
            .in0(_gnd_net_),
            .in1(N__54948),
            .in2(N__23161),
            .in3(N__21667),
            .lcout(n1888),
            .ltout(),
            .carryin(n12218),
            .carryout(n12219),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_1_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_1_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_1_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_16_lut_LC_1_24_6 (
            .in0(_gnd_net_),
            .in1(N__54946),
            .in2(N__23193),
            .in3(N__21664),
            .lcout(n1887),
            .ltout(),
            .carryin(n12219),
            .carryout(n12220),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_1_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_1_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_1_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_17_lut_LC_1_24_7 (
            .in0(_gnd_net_),
            .in1(N__54949),
            .in2(N__24385),
            .in3(N__21661),
            .lcout(n1886),
            .ltout(),
            .carryin(n12220),
            .carryout(n12221),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_1_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_1_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_1_25_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 encoder0_position_31__I_0_add_1235_18_lut_LC_1_25_0 (
            .in0(N__54950),
            .in1(_gnd_net_),
            .in2(N__27414),
            .in3(N__21658),
            .lcout(n1885),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_1_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_1_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_1_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_2_lut_LC_1_26_0 (
            .in0(_gnd_net_),
            .in1(N__28098),
            .in2(_gnd_net_),
            .in3(N__21655),
            .lcout(n1701),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(n12177),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_1_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_1_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_1_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_3_lut_LC_1_26_1 (
            .in0(_gnd_net_),
            .in1(N__54581),
            .in2(N__23448),
            .in3(N__21652),
            .lcout(n1700),
            .ltout(),
            .carryin(n12177),
            .carryout(n12178),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_1_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_1_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_1_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_4_lut_LC_1_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23473),
            .in3(N__21649),
            .lcout(n1699),
            .ltout(),
            .carryin(n12178),
            .carryout(n12179),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_1_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_1_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_1_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_5_lut_LC_1_26_3 (
            .in0(_gnd_net_),
            .in1(N__54582),
            .in2(N__22339),
            .in3(N__21700),
            .lcout(n1698),
            .ltout(),
            .carryin(n12179),
            .carryout(n12180),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_1_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_1_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_1_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_6_lut_LC_1_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22263),
            .in3(N__21697),
            .lcout(n1697),
            .ltout(),
            .carryin(n12180),
            .carryout(n12181),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_1_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_1_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_1_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_7_lut_LC_1_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22360),
            .in3(N__21694),
            .lcout(n1696),
            .ltout(),
            .carryin(n12181),
            .carryout(n12182),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_1_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_1_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_1_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_8_lut_LC_1_26_6 (
            .in0(_gnd_net_),
            .in1(N__54951),
            .in2(N__23289),
            .in3(N__21691),
            .lcout(n1695),
            .ltout(),
            .carryin(n12182),
            .carryout(n12183),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_1_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_1_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_1_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_9_lut_LC_1_26_7 (
            .in0(_gnd_net_),
            .in1(N__54583),
            .in2(N__23668),
            .in3(N__21688),
            .lcout(n1694),
            .ltout(),
            .carryin(n12183),
            .carryout(n12184),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_1_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_1_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_1_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_10_lut_LC_1_27_0 (
            .in0(_gnd_net_),
            .in1(N__55135),
            .in2(N__23506),
            .in3(N__21685),
            .lcout(n1693),
            .ltout(),
            .carryin(bfn_1_27_0_),
            .carryout(n12185),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_1_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_1_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_1_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_11_lut_LC_1_27_1 (
            .in0(_gnd_net_),
            .in1(N__55140),
            .in2(N__23419),
            .in3(N__21682),
            .lcout(n1692),
            .ltout(),
            .carryin(n12185),
            .carryout(n12186),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_1_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_1_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_1_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_12_lut_LC_1_27_2 (
            .in0(_gnd_net_),
            .in1(N__55136),
            .in2(N__23260),
            .in3(N__21679),
            .lcout(n1691),
            .ltout(),
            .carryin(n12186),
            .carryout(n12187),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_1_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_1_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_1_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_13_lut_LC_1_27_3 (
            .in0(_gnd_net_),
            .in1(N__55141),
            .in2(N__23395),
            .in3(N__21676),
            .lcout(n1690),
            .ltout(),
            .carryin(n12187),
            .carryout(n12188),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_1_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_1_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_1_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_14_lut_LC_1_27_4 (
            .in0(_gnd_net_),
            .in1(N__23604),
            .in2(N__55219),
            .in3(N__21727),
            .lcout(n1689),
            .ltout(),
            .carryin(n12188),
            .carryout(n12189),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_1_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_1_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_1_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_15_lut_LC_1_27_5 (
            .in0(_gnd_net_),
            .in1(N__23532),
            .in2(N__55218),
            .in3(N__21724),
            .lcout(n1688),
            .ltout(),
            .carryin(n12189),
            .carryout(n12190),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_1_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_1_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_1_27_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1101_16_lut_LC_1_27_6 (
            .in0(N__55145),
            .in1(N__35520),
            .in2(N__25642),
            .in3(N__21721),
            .lcout(n1719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i907_3_lut_LC_1_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_1_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_1_28_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i907_3_lut_LC_1_28_0 (
            .in0(_gnd_net_),
            .in1(N__23797),
            .in2(N__28336),
            .in3(N__36743),
            .lcout(n1427),
            .ltout(n1427_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_73_LC_1_28_1.C_ON=1'b0;
    defparam i1_2_lut_adj_73_LC_1_28_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_73_LC_1_28_1.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_73_LC_1_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21718),
            .in3(N__25515),
            .lcout(n14088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i910_3_lut_LC_1_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_1_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_1_28_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i910_3_lut_LC_1_28_4 (
            .in0(_gnd_net_),
            .in1(N__23818),
            .in2(N__26194),
            .in3(N__36744),
            .lcout(n1430),
            .ltout(n1430_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_74_LC_1_28_5.C_ON=1'b0;
    defparam i1_4_lut_adj_74_LC_1_28_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_74_LC_1_28_5.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_74_LC_1_28_5 (
            .in0(N__25938),
            .in1(N__26061),
            .in2(N__21715),
            .in3(N__21712),
            .lcout(n13334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9924_3_lut_LC_1_28_6.C_ON=1'b0;
    defparam i9924_3_lut_LC_1_28_6.SEQ_MODE=4'b0000;
    defparam i9924_3_lut_LC_1_28_6.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9924_3_lut_LC_1_28_6 (
            .in0(_gnd_net_),
            .in1(N__23578),
            .in2(N__23707),
            .in3(N__23741),
            .lcout(n11638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.cnt_reg_636__i0_LC_1_29_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i0_LC_1_29_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i0_LC_1_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i0_LC_1_29_0  (
            .in0(_gnd_net_),
            .in1(N__22650),
            .in2(_gnd_net_),
            .in3(N__21706),
            .lcout(\debounce.cnt_reg_0 ),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(\debounce.n12654 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i1_LC_1_29_1 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i1_LC_1_29_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i1_LC_1_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i1_LC_1_29_1  (
            .in0(_gnd_net_),
            .in1(N__21855),
            .in2(_gnd_net_),
            .in3(N__21703),
            .lcout(\debounce.cnt_reg_1 ),
            .ltout(),
            .carryin(\debounce.n12654 ),
            .carryout(\debounce.n12655 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i2_LC_1_29_2 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i2_LC_1_29_2 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i2_LC_1_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i2_LC_1_29_2  (
            .in0(_gnd_net_),
            .in1(N__21840),
            .in2(_gnd_net_),
            .in3(N__21754),
            .lcout(\debounce.cnt_reg_2 ),
            .ltout(),
            .carryin(\debounce.n12655 ),
            .carryout(\debounce.n12656 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i3_LC_1_29_3 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i3_LC_1_29_3 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i3_LC_1_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i3_LC_1_29_3  (
            .in0(_gnd_net_),
            .in1(N__21918),
            .in2(_gnd_net_),
            .in3(N__21751),
            .lcout(\debounce.cnt_reg_3 ),
            .ltout(),
            .carryin(\debounce.n12656 ),
            .carryout(\debounce.n12657 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i4_LC_1_29_4 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i4_LC_1_29_4 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i4_LC_1_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i4_LC_1_29_4  (
            .in0(_gnd_net_),
            .in1(N__22686),
            .in2(_gnd_net_),
            .in3(N__21748),
            .lcout(\debounce.cnt_reg_4 ),
            .ltout(),
            .carryin(\debounce.n12657 ),
            .carryout(\debounce.n12658 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i5_LC_1_29_5 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i5_LC_1_29_5 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i5_LC_1_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i5_LC_1_29_5  (
            .in0(_gnd_net_),
            .in1(N__21885),
            .in2(_gnd_net_),
            .in3(N__21745),
            .lcout(\debounce.cnt_reg_5 ),
            .ltout(),
            .carryin(\debounce.n12658 ),
            .carryout(\debounce.n12659 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i6_LC_1_29_6 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i6_LC_1_29_6 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i6_LC_1_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i6_LC_1_29_6  (
            .in0(_gnd_net_),
            .in1(N__22671),
            .in2(_gnd_net_),
            .in3(N__21742),
            .lcout(\debounce.cnt_reg_6 ),
            .ltout(),
            .carryin(\debounce.n12659 ),
            .carryout(\debounce.n12660 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i7_LC_1_29_7 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i7_LC_1_29_7 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i7_LC_1_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i7_LC_1_29_7  (
            .in0(_gnd_net_),
            .in1(N__22635),
            .in2(_gnd_net_),
            .in3(N__21739),
            .lcout(\debounce.cnt_reg_7 ),
            .ltout(),
            .carryin(\debounce.n12660 ),
            .carryout(\debounce.n12661 ),
            .clk(N__56042),
            .ce(),
            .sr(N__23887));
    defparam \debounce.cnt_reg_636__i8_LC_1_30_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_636__i8_LC_1_30_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i8_LC_1_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i8_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(N__21870),
            .in2(_gnd_net_),
            .in3(N__21736),
            .lcout(\debounce.cnt_reg_8 ),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(\debounce.n12662 ),
            .clk(N__56044),
            .ce(),
            .sr(N__23886));
    defparam \debounce.cnt_reg_636__i9_LC_1_30_1 .C_ON=1'b0;
    defparam \debounce.cnt_reg_636__i9_LC_1_30_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_636__i9_LC_1_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_636__i9_LC_1_30_1  (
            .in0(_gnd_net_),
            .in1(N__21903),
            .in2(_gnd_net_),
            .in3(N__21733),
            .lcout(\debounce.cnt_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56044),
            .ce(),
            .sr(N__23886));
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_1_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_1_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_1_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_2_lut_LC_1_31_0 (
            .in0(_gnd_net_),
            .in1(N__28176),
            .in2(_gnd_net_),
            .in3(N__21730),
            .lcout(n1201),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(n12122),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_1_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_1_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_1_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_3_lut_LC_1_31_1 (
            .in0(_gnd_net_),
            .in1(N__55220),
            .in2(N__28633),
            .in3(N__21781),
            .lcout(n1200),
            .ltout(),
            .carryin(n12122),
            .carryout(n12123),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_1_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_1_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_1_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_4_lut_LC_1_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28687),
            .in3(N__21778),
            .lcout(n1199),
            .ltout(),
            .carryin(n12123),
            .carryout(n12124),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_1_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_1_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_1_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_5_lut_LC_1_31_3 (
            .in0(_gnd_net_),
            .in1(N__55221),
            .in2(N__30457),
            .in3(N__21775),
            .lcout(n1198),
            .ltout(),
            .carryin(n12124),
            .carryout(n12125),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_1_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_1_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_1_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_6_lut_LC_1_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26395),
            .in3(N__21772),
            .lcout(n1197),
            .ltout(),
            .carryin(n12125),
            .carryout(n12126),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_1_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_1_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_1_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_7_lut_LC_1_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28663),
            .in3(N__21769),
            .lcout(n1196),
            .ltout(),
            .carryin(n12126),
            .carryout(n12127),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_1_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_1_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_1_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_8_lut_LC_1_31_6 (
            .in0(_gnd_net_),
            .in1(N__55223),
            .in2(N__30550),
            .in3(N__21766),
            .lcout(n1195),
            .ltout(),
            .carryin(n12127),
            .carryout(n12128),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_1_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_1_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_1_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_9_lut_LC_1_31_7 (
            .in0(_gnd_net_),
            .in1(N__55222),
            .in2(N__28765),
            .in3(N__21763),
            .lcout(n1194),
            .ltout(),
            .carryin(n12128),
            .carryout(n12129),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_1_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_1_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_1_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_10_lut_LC_1_32_0 (
            .in0(_gnd_net_),
            .in1(N__55224),
            .in2(N__28788),
            .in3(N__21760),
            .lcout(n1193),
            .ltout(),
            .carryin(bfn_1_32_0_),
            .carryout(n12130),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_1_32_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_1_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_1_32_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_766_11_lut_LC_1_32_1 (
            .in0(N__55225),
            .in1(N__36570),
            .in2(N__28807),
            .in3(N__21757),
            .lcout(n1224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i12061_4_lut_LC_1_32_2 .C_ON=1'b0;
    defparam \debounce.i12061_4_lut_LC_1_32_2 .SEQ_MODE=4'b0000;
    defparam \debounce.i12061_4_lut_LC_1_32_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \debounce.i12061_4_lut_LC_1_32_2  (
            .in0(N__21919),
            .in1(N__21904),
            .in2(N__21889),
            .in3(N__21871),
            .lcout(),
            .ltout(\debounce.n14472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i2_4_lut_LC_1_32_3 .C_ON=1'b0;
    defparam \debounce.i2_4_lut_LC_1_32_3 .SEQ_MODE=4'b0000;
    defparam \debounce.i2_4_lut_LC_1_32_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \debounce.i2_4_lut_LC_1_32_3  (
            .in0(N__21856),
            .in1(N__21841),
            .in2(N__21826),
            .in3(N__22621),
            .lcout(n13490),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_2_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_2_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_2_18_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1383_3_lut_LC_2_18_0 (
            .in0(_gnd_net_),
            .in1(N__21823),
            .in2(N__23035),
            .in3(N__35987),
            .lcout(n2127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_2_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_2_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_2_18_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1382_3_lut_LC_2_18_1 (
            .in0(_gnd_net_),
            .in1(N__21814),
            .in2(N__36017),
            .in3(N__24660),
            .lcout(n2126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_2_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_2_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_2_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_2_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37554),
            .lcout(n23_adj_647),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_2_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_2_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_2_18_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1389_3_lut_LC_2_18_4 (
            .in0(N__21802),
            .in1(N__27921),
            .in2(_gnd_net_),
            .in3(N__35986),
            .lcout(n2133),
            .ltout(n2133_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_2_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_2_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_2_18_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1456_3_lut_LC_2_18_5 (
            .in0(N__21793),
            .in1(_gnd_net_),
            .in2(N__21787),
            .in3(N__36168),
            .lcout(n2232),
            .ltout(n2232_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_2_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_2_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_2_18_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1523_3_lut_LC_2_18_6 (
            .in0(N__31456),
            .in1(_gnd_net_),
            .in2(N__21784),
            .in3(N__39145),
            .lcout(n2331),
            .ltout(n2331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_2_18_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1590_3_lut_LC_2_18_7 (
            .in0(_gnd_net_),
            .in1(N__22606),
            .in2(N__21970),
            .in3(N__34929),
            .lcout(n2430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12587_1_lut_LC_2_19_0.C_ON=1'b0;
    defparam i12587_1_lut_LC_2_19_0.SEQ_MODE=4'b0000;
    defparam i12587_1_lut_LC_2_19_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12587_1_lut_LC_2_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36158),
            .lcout(n15059),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_2_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_2_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_2_19_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1377_3_lut_LC_2_19_1 (
            .in0(_gnd_net_),
            .in1(N__24166),
            .in2(N__21967),
            .in3(N__35993),
            .lcout(n2121),
            .ltout(n2121_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_2_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_2_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_2_19_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1444_3_lut_LC_2_19_2 (
            .in0(_gnd_net_),
            .in1(N__21955),
            .in2(N__21949),
            .in3(N__36157),
            .lcout(n2220),
            .ltout(n2220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_2_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_2_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_2_19_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1511_3_lut_LC_2_19_3 (
            .in0(_gnd_net_),
            .in1(N__31642),
            .in2(N__21946),
            .in3(N__39134),
            .lcout(n2319),
            .ltout(n2319_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_2_19_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1578_3_lut_LC_2_19_4 (
            .in0(_gnd_net_),
            .in1(N__22750),
            .in2(N__21943),
            .in3(N__34935),
            .lcout(n2418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12566_4_lut_LC_2_19_6.C_ON=1'b0;
    defparam i12566_4_lut_LC_2_19_6.SEQ_MODE=4'b0000;
    defparam i12566_4_lut_LC_2_19_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12566_4_lut_LC_2_19_6 (
            .in0(N__22125),
            .in1(N__22929),
            .in2(N__22165),
            .in3(N__22774),
            .lcout(n2049),
            .ltout(n2049_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_2_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_2_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_2_19_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1385_3_lut_LC_2_19_7 (
            .in0(N__21940),
            .in1(_gnd_net_),
            .in2(N__21934),
            .in3(N__24240),
            .lcout(n2129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_2_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_2_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_2_20_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1439_3_lut_LC_2_20_0 (
            .in0(_gnd_net_),
            .in1(N__21931),
            .in2(N__22063),
            .in3(N__36159),
            .lcout(n2215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_2_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_2_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_2_20_1.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1440_3_lut_LC_2_20_1 (
            .in0(N__21990),
            .in1(N__21925),
            .in2(N__36193),
            .in3(_gnd_net_),
            .lcout(n2216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_2_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_2_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_2_20_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1372_3_lut_LC_2_20_2 (
            .in0(_gnd_net_),
            .in1(N__22072),
            .in2(N__22132),
            .in3(N__35985),
            .lcout(n2116),
            .ltout(n2116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12590_4_lut_LC_2_20_3.C_ON=1'b0;
    defparam i12590_4_lut_LC_2_20_3.SEQ_MODE=4'b0000;
    defparam i12590_4_lut_LC_2_20_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12590_4_lut_LC_2_20_3 (
            .in0(N__21989),
            .in1(N__22044),
            .in2(N__22030),
            .in3(N__27022),
            .lcout(n2148),
            .ltout(n2148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_2_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_2_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_2_20_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1451_3_lut_LC_2_20_4 (
            .in0(_gnd_net_),
            .in1(N__24561),
            .in2(N__22027),
            .in3(N__22024),
            .lcout(n2227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_2_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_2_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_2_20_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1375_3_lut_LC_2_20_5 (
            .in0(N__22015),
            .in1(_gnd_net_),
            .in2(N__36015),
            .in3(N__22889),
            .lcout(n2119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_2_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_2_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_2_20_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1381_3_lut_LC_2_20_6 (
            .in0(_gnd_net_),
            .in1(N__22009),
            .in2(N__22980),
            .in3(N__35978),
            .lcout(n2125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_2_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_2_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_2_20_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1373_3_lut_LC_2_20_7 (
            .in0(N__22922),
            .in1(_gnd_net_),
            .in2(N__36016),
            .in3(N__22003),
            .lcout(n2117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_2_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_2_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_2_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_2_lut_LC_2_21_0 (
            .in0(_gnd_net_),
            .in1(N__37603),
            .in2(_gnd_net_),
            .in3(N__21976),
            .lcout(n2001),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(n12222),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_2_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_2_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_2_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_3_lut_LC_2_21_1 (
            .in0(_gnd_net_),
            .in1(N__53790),
            .in2(N__27493),
            .in3(N__21973),
            .lcout(n2000),
            .ltout(),
            .carryin(n12222),
            .carryout(n12223),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_2_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_2_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_2_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_4_lut_LC_2_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26935),
            .in3(N__22102),
            .lcout(n1999),
            .ltout(),
            .carryin(n12223),
            .carryout(n12224),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_2_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_2_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_2_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_5_lut_LC_2_21_3 (
            .in0(_gnd_net_),
            .in1(N__53791),
            .in2(N__26908),
            .in3(N__22099),
            .lcout(n1998),
            .ltout(),
            .carryin(n12224),
            .carryout(n12225),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_2_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_2_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_2_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_6_lut_LC_2_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27454),
            .in3(N__22096),
            .lcout(n1997),
            .ltout(),
            .carryin(n12225),
            .carryout(n12226),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_2_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_2_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_2_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_7_lut_LC_2_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27538),
            .in3(N__22093),
            .lcout(n1996),
            .ltout(),
            .carryin(n12226),
            .carryout(n12227),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_2_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_2_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_2_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_8_lut_LC_2_21_6 (
            .in0(_gnd_net_),
            .in1(N__54254),
            .in2(N__24693),
            .in3(N__22090),
            .lcout(n1995),
            .ltout(),
            .carryin(n12227),
            .carryout(n12228),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_2_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_2_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_2_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_9_lut_LC_2_21_7 (
            .in0(_gnd_net_),
            .in1(N__53792),
            .in2(N__24805),
            .in3(N__22087),
            .lcout(n1994),
            .ltout(),
            .carryin(n12228),
            .carryout(n12229),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_2_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_2_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_2_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_10_lut_LC_2_22_0 (
            .in0(_gnd_net_),
            .in1(N__54255),
            .in2(N__24499),
            .in3(N__22084),
            .lcout(n1993),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(n12230),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_2_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_2_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_2_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_11_lut_LC_2_22_1 (
            .in0(_gnd_net_),
            .in1(N__54926),
            .in2(N__24408),
            .in3(N__22081),
            .lcout(n1992),
            .ltout(),
            .carryin(n12230),
            .carryout(n12231),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_2_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_2_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_2_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_12_lut_LC_2_22_2 (
            .in0(_gnd_net_),
            .in1(N__54256),
            .in2(N__23112),
            .in3(N__22078),
            .lcout(n1991),
            .ltout(),
            .carryin(n12231),
            .carryout(n12232),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_2_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_2_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_2_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_13_lut_LC_2_22_3 (
            .in0(_gnd_net_),
            .in1(N__54927),
            .in2(N__24183),
            .in3(N__22075),
            .lcout(n1990),
            .ltout(),
            .carryin(n12232),
            .carryout(n12233),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_2_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_2_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_2_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_14_lut_LC_2_22_4 (
            .in0(_gnd_net_),
            .in1(N__24765),
            .in2(N__55132),
            .in3(N__22183),
            .lcout(n1989),
            .ltout(),
            .carryin(n12233),
            .carryout(n12234),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_2_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_2_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_2_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_15_lut_LC_2_22_5 (
            .in0(_gnd_net_),
            .in1(N__26973),
            .in2(N__54729),
            .in3(N__22180),
            .lcout(n1988),
            .ltout(),
            .carryin(n12234),
            .carryout(n12235),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_2_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_2_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_2_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_16_lut_LC_2_22_6 (
            .in0(_gnd_net_),
            .in1(N__24725),
            .in2(N__55133),
            .in3(N__22177),
            .lcout(n1987),
            .ltout(),
            .carryin(n12235),
            .carryout(n12236),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_2_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_2_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_2_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_17_lut_LC_2_22_7 (
            .in0(_gnd_net_),
            .in1(N__24513),
            .in2(N__54730),
            .in3(N__22174),
            .lcout(n1986),
            .ltout(),
            .carryin(n12236),
            .carryout(n12237),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_2_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_2_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_2_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_18_lut_LC_2_23_0 (
            .in0(_gnd_net_),
            .in1(N__24530),
            .in2(N__54731),
            .in3(N__22171),
            .lcout(n1985),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(n12238),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_2_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_2_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_2_23_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1302_19_lut_LC_2_23_1 (
            .in0(N__54266),
            .in1(N__35910),
            .in2(N__27379),
            .in3(N__22168),
            .lcout(n2016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_2_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_2_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_2_23_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1240_3_lut_LC_2_23_2 (
            .in0(_gnd_net_),
            .in1(N__22144),
            .in2(N__23160),
            .in3(N__35765),
            .lcout(n1920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_2_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_2_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_2_23_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1182_3_lut_LC_2_23_3 (
            .in0(_gnd_net_),
            .in1(N__24978),
            .in2(N__24964),
            .in3(N__35594),
            .lcout(n1830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_2_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_2_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_2_23_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1305_3_lut_LC_2_23_7 (
            .in0(N__35895),
            .in1(N__22138),
            .in2(N__24537),
            .in3(_gnd_net_),
            .lcout(n2017),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_2_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_2_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_2_24_0.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i1116_3_lut_LC_2_24_0 (
            .in0(N__35481),
            .in1(N__23449),
            .in2(N__22240),
            .in3(_gnd_net_),
            .lcout(n1732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_2_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_2_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_2_24_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_i1115_3_lut_LC_2_24_1 (
            .in0(N__23472),
            .in1(N__35482),
            .in2(_gnd_net_),
            .in3(N__22228),
            .lcout(n1731),
            .ltout(n1731_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9979_4_lut_LC_2_24_2.C_ON=1'b0;
    defparam i9979_4_lut_LC_2_24_2.SEQ_MODE=4'b0000;
    defparam i9979_4_lut_LC_2_24_2.LUT_INIT=16'b1111111011110000;
    LogicCell40 i9979_4_lut_LC_2_24_2 (
            .in0(N__28048),
            .in1(N__25044),
            .in2(N__22219),
            .in3(N__25004),
            .lcout(n11694),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_2_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_2_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_2_24_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1113_3_lut_LC_2_24_3 (
            .in0(_gnd_net_),
            .in1(N__35483),
            .in2(N__22267),
            .in3(N__22216),
            .lcout(n1729),
            .ltout(n1729_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_81_LC_2_24_4.C_ON=1'b0;
    defparam i1_2_lut_adj_81_LC_2_24_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_81_LC_2_24_4.LUT_INIT=16'b1100000011000000;
    LogicCell40 i1_2_lut_adj_81_LC_2_24_4 (
            .in0(_gnd_net_),
            .in1(N__24927),
            .in2(N__22207),
            .in3(_gnd_net_),
            .lcout(n14116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_2_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_2_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_2_24_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1117_3_lut_LC_2_24_5 (
            .in0(N__22204),
            .in1(N__28099),
            .in2(_gnd_net_),
            .in3(N__35480),
            .lcout(n1733),
            .ltout(n1733_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_2_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_2_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_2_24_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1184_3_lut_LC_2_24_6 (
            .in0(_gnd_net_),
            .in1(N__25033),
            .in2(N__22195),
            .in3(N__35584),
            .lcout(n1832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_2_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_2_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_2_24_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1238_3_lut_LC_2_24_7 (
            .in0(_gnd_net_),
            .in1(N__24377),
            .in2(N__22192),
            .in3(N__35766),
            .lcout(n1918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_148_LC_2_25_0.C_ON=1'b0;
    defparam i1_4_lut_adj_148_LC_2_25_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_148_LC_2_25_0.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_148_LC_2_25_0 (
            .in0(N__22334),
            .in1(N__22256),
            .in2(N__22359),
            .in3(N__23425),
            .lcout(n13343),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_2_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_2_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_2_25_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1114_3_lut_LC_2_25_1 (
            .in0(_gnd_net_),
            .in1(N__22312),
            .in2(N__35492),
            .in3(N__22335),
            .lcout(n1730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_2_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_2_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_2_25_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1112_3_lut_LC_2_25_2 (
            .in0(N__22355),
            .in1(_gnd_net_),
            .in2(N__22306),
            .in3(N__35476),
            .lcout(n1728),
            .ltout(n1728_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_79_LC_2_25_3.C_ON=1'b0;
    defparam i1_3_lut_adj_79_LC_2_25_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_79_LC_2_25_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_79_LC_2_25_3 (
            .in0(_gnd_net_),
            .in1(N__24848),
            .in2(N__22297),
            .in3(N__27872),
            .lcout(n13962),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12374_3_lut_LC_2_25_4.C_ON=1'b0;
    defparam i12374_3_lut_LC_2_25_4.SEQ_MODE=4'b0000;
    defparam i12374_3_lut_LC_2_25_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12374_3_lut_LC_2_25_4 (
            .in0(_gnd_net_),
            .in1(N__22294),
            .in2(N__23290),
            .in3(N__35469),
            .lcout(n1727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12477_1_lut_LC_2_25_5.C_ON=1'b0;
    defparam i12477_1_lut_LC_2_25_5.SEQ_MODE=4'b0000;
    defparam i12477_1_lut_LC_2_25_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12477_1_lut_LC_2_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35491),
            .in3(_gnd_net_),
            .lcout(n14949),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1110_3_lut_LC_2_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1110_3_lut_LC_2_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1110_3_lut_LC_2_25_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1110_3_lut_LC_2_25_6 (
            .in0(_gnd_net_),
            .in1(N__23663),
            .in2(N__22288),
            .in3(N__35468),
            .lcout(n1726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_2_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_2_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_2_25_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1105_3_lut_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(N__23611),
            .in2(N__35493),
            .in3(N__22279),
            .lcout(n1721),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_2_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_2_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_2_26_0.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1046_3_lut_LC_2_26_0 (
            .in0(N__25402),
            .in1(N__25416),
            .in2(N__35388),
            .in3(_gnd_net_),
            .lcout(n1630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_2_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_2_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_2_26_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1049_3_lut_LC_2_26_1 (
            .in0(_gnd_net_),
            .in1(N__25060),
            .in2(N__27574),
            .in3(N__35364),
            .lcout(n1633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_127_LC_2_26_2.C_ON=1'b0;
    defparam i1_4_lut_adj_127_LC_2_26_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_127_LC_2_26_2.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_127_LC_2_26_2 (
            .in0(N__25352),
            .in1(N__23356),
            .in2(N__25389),
            .in3(N__23752),
            .lcout(),
            .ltout(n13986_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12825_4_lut_LC_2_26_3.C_ON=1'b0;
    defparam i12825_4_lut_LC_2_26_3.SEQ_MODE=4'b0000;
    defparam i12825_4_lut_LC_2_26_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12825_4_lut_LC_2_26_3 (
            .in0(N__25725),
            .in1(N__25689),
            .in2(N__22366),
            .in3(N__25662),
            .lcout(n1554),
            .ltout(n1554_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_2_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_2_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_2_26_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1042_3_lut_LC_2_26_4 (
            .in0(N__25296),
            .in1(_gnd_net_),
            .in2(N__22363),
            .in3(N__25270),
            .lcout(n1626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_2_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_2_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_2_26_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_2_26_5 (
            .in0(_gnd_net_),
            .in1(N__25353),
            .in2(N__25339),
            .in3(N__35365),
            .lcout(n1628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_2_26_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_2_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_2_26_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1045_3_lut_LC_2_26_6 (
            .in0(N__25385),
            .in1(_gnd_net_),
            .in2(N__35389),
            .in3(N__25369),
            .lcout(n1629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_2_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_2_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_2_26_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1047_3_lut_LC_2_26_7 (
            .in0(_gnd_net_),
            .in1(N__25462),
            .in2(N__25432),
            .in3(N__35372),
            .lcout(n1631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_2_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_2_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_2_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_2_lut_LC_2_27_0 (
            .in0(_gnd_net_),
            .in1(N__23577),
            .in2(_gnd_net_),
            .in3(N__22321),
            .lcout(n1501),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(n12152),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_2_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_2_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_2_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_3_lut_LC_2_27_1 (
            .in0(_gnd_net_),
            .in1(N__54732),
            .in2(N__23706),
            .in3(N__22318),
            .lcout(n1500),
            .ltout(),
            .carryin(n12152),
            .carryout(n12153),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_2_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_2_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_2_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_4_lut_LC_2_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23742),
            .in3(N__22315),
            .lcout(n1499),
            .ltout(),
            .carryin(n12153),
            .carryout(n12154),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_2_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_2_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_2_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_5_lut_LC_2_27_3 (
            .in0(_gnd_net_),
            .in1(N__54733),
            .in2(N__25942),
            .in3(N__22396),
            .lcout(n1498),
            .ltout(),
            .carryin(n12154),
            .carryout(n12155),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_2_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_2_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_2_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_6_lut_LC_2_27_4 (
            .in0(_gnd_net_),
            .in1(N__23634),
            .in2(_gnd_net_),
            .in3(N__22393),
            .lcout(n1497),
            .ltout(),
            .carryin(n12155),
            .carryout(n12156),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_2_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_2_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_2_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_7_lut_LC_2_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26065),
            .in3(N__22390),
            .lcout(n1496),
            .ltout(),
            .carryin(n12156),
            .carryout(n12157),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_2_27_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_2_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_2_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_8_lut_LC_2_27_6 (
            .in0(_gnd_net_),
            .in1(N__54734),
            .in2(N__25522),
            .in3(N__22387),
            .lcout(n1495),
            .ltout(),
            .carryin(n12157),
            .carryout(n12158),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_2_27_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_2_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_2_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_9_lut_LC_2_27_7 (
            .in0(_gnd_net_),
            .in1(N__25614),
            .in2(N__55061),
            .in3(N__22384),
            .lcout(n1494),
            .ltout(),
            .carryin(n12158),
            .carryout(n12159),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_2_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_2_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_2_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_10_lut_LC_2_28_0 (
            .in0(_gnd_net_),
            .in1(N__54744),
            .in2(N__25972),
            .in3(N__22381),
            .lcout(n1493),
            .ltout(),
            .carryin(bfn_2_28_0_),
            .carryout(n12160),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_2_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_2_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_2_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_11_lut_LC_2_28_1 (
            .in0(_gnd_net_),
            .in1(N__25846),
            .in2(N__55062),
            .in3(N__22378),
            .lcout(n1492),
            .ltout(),
            .carryin(n12160),
            .carryout(n12161),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_2_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_2_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_2_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_12_lut_LC_2_28_2 (
            .in0(_gnd_net_),
            .in1(N__54748),
            .in2(N__26134),
            .in3(N__22375),
            .lcout(n1491),
            .ltout(),
            .carryin(n12161),
            .carryout(n12162),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_2_28_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_2_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_2_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_13_lut_LC_2_28_3 (
            .in0(_gnd_net_),
            .in1(N__54742),
            .in2(N__25900),
            .in3(N__22372),
            .lcout(n1490),
            .ltout(),
            .carryin(n12162),
            .carryout(n12163),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_2_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_2_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_2_28_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_967_14_lut_LC_2_28_4 (
            .in0(N__54743),
            .in1(N__25882),
            .in2(N__35310),
            .in3(N__22369),
            .lcout(n1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12804_1_lut_LC_2_28_6.C_ON=1'b0;
    defparam i12804_1_lut_LC_2_28_6.SEQ_MODE=4'b0000;
    defparam i12804_1_lut_LC_2_28_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12804_1_lut_LC_2_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35275),
            .lcout(n15276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i971_3_lut_LC_2_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_2_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_2_28_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i971_3_lut_LC_2_28_7 (
            .in0(_gnd_net_),
            .in1(N__26133),
            .in2(N__35286),
            .in3(N__22456),
            .lcout(n1523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i0_LC_2_29_0.C_ON=1'b1;
    defparam blink_counter_634__i0_LC_2_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i0_LC_2_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i0_LC_2_29_0 (
            .in0(_gnd_net_),
            .in1(N__22450),
            .in2(_gnd_net_),
            .in3(N__22444),
            .lcout(n26_adj_678),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(n12717),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i1_LC_2_29_1.C_ON=1'b1;
    defparam blink_counter_634__i1_LC_2_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i1_LC_2_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i1_LC_2_29_1 (
            .in0(_gnd_net_),
            .in1(N__22441),
            .in2(_gnd_net_),
            .in3(N__22435),
            .lcout(n25_adj_677),
            .ltout(),
            .carryin(n12717),
            .carryout(n12718),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i2_LC_2_29_2.C_ON=1'b1;
    defparam blink_counter_634__i2_LC_2_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i2_LC_2_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i2_LC_2_29_2 (
            .in0(_gnd_net_),
            .in1(N__22432),
            .in2(_gnd_net_),
            .in3(N__22426),
            .lcout(n24_adj_676),
            .ltout(),
            .carryin(n12718),
            .carryout(n12719),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i3_LC_2_29_3.C_ON=1'b1;
    defparam blink_counter_634__i3_LC_2_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i3_LC_2_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i3_LC_2_29_3 (
            .in0(_gnd_net_),
            .in1(N__22423),
            .in2(_gnd_net_),
            .in3(N__22417),
            .lcout(n23_adj_675),
            .ltout(),
            .carryin(n12719),
            .carryout(n12720),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i4_LC_2_29_4.C_ON=1'b1;
    defparam blink_counter_634__i4_LC_2_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i4_LC_2_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i4_LC_2_29_4 (
            .in0(_gnd_net_),
            .in1(N__22414),
            .in2(_gnd_net_),
            .in3(N__22408),
            .lcout(n22_adj_674),
            .ltout(),
            .carryin(n12720),
            .carryout(n12721),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i5_LC_2_29_5.C_ON=1'b1;
    defparam blink_counter_634__i5_LC_2_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i5_LC_2_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i5_LC_2_29_5 (
            .in0(_gnd_net_),
            .in1(N__22405),
            .in2(_gnd_net_),
            .in3(N__22399),
            .lcout(n21_adj_673),
            .ltout(),
            .carryin(n12721),
            .carryout(n12722),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i6_LC_2_29_6.C_ON=1'b1;
    defparam blink_counter_634__i6_LC_2_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i6_LC_2_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i6_LC_2_29_6 (
            .in0(_gnd_net_),
            .in1(N__22537),
            .in2(_gnd_net_),
            .in3(N__22531),
            .lcout(n20_adj_672),
            .ltout(),
            .carryin(n12722),
            .carryout(n12723),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i7_LC_2_29_7.C_ON=1'b1;
    defparam blink_counter_634__i7_LC_2_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i7_LC_2_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i7_LC_2_29_7 (
            .in0(_gnd_net_),
            .in1(N__22528),
            .in2(_gnd_net_),
            .in3(N__22522),
            .lcout(n19_adj_671),
            .ltout(),
            .carryin(n12723),
            .carryout(n12724),
            .clk(N__56045),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i8_LC_2_30_0.C_ON=1'b1;
    defparam blink_counter_634__i8_LC_2_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i8_LC_2_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i8_LC_2_30_0 (
            .in0(_gnd_net_),
            .in1(N__22519),
            .in2(_gnd_net_),
            .in3(N__22513),
            .lcout(n18_adj_670),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(n12725),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i9_LC_2_30_1.C_ON=1'b1;
    defparam blink_counter_634__i9_LC_2_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i9_LC_2_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i9_LC_2_30_1 (
            .in0(_gnd_net_),
            .in1(N__22510),
            .in2(_gnd_net_),
            .in3(N__22504),
            .lcout(n17_adj_669),
            .ltout(),
            .carryin(n12725),
            .carryout(n12726),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i10_LC_2_30_2.C_ON=1'b1;
    defparam blink_counter_634__i10_LC_2_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i10_LC_2_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i10_LC_2_30_2 (
            .in0(_gnd_net_),
            .in1(N__22501),
            .in2(_gnd_net_),
            .in3(N__22495),
            .lcout(n16_adj_668),
            .ltout(),
            .carryin(n12726),
            .carryout(n12727),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i11_LC_2_30_3.C_ON=1'b1;
    defparam blink_counter_634__i11_LC_2_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i11_LC_2_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i11_LC_2_30_3 (
            .in0(_gnd_net_),
            .in1(N__22492),
            .in2(_gnd_net_),
            .in3(N__22486),
            .lcout(n15_adj_667),
            .ltout(),
            .carryin(n12727),
            .carryout(n12728),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i12_LC_2_30_4.C_ON=1'b1;
    defparam blink_counter_634__i12_LC_2_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i12_LC_2_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i12_LC_2_30_4 (
            .in0(_gnd_net_),
            .in1(N__22483),
            .in2(_gnd_net_),
            .in3(N__22477),
            .lcout(n14_adj_666),
            .ltout(),
            .carryin(n12728),
            .carryout(n12729),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i13_LC_2_30_5.C_ON=1'b1;
    defparam blink_counter_634__i13_LC_2_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i13_LC_2_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i13_LC_2_30_5 (
            .in0(_gnd_net_),
            .in1(N__22474),
            .in2(_gnd_net_),
            .in3(N__22468),
            .lcout(n13_adj_665),
            .ltout(),
            .carryin(n12729),
            .carryout(n12730),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i14_LC_2_30_6.C_ON=1'b1;
    defparam blink_counter_634__i14_LC_2_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i14_LC_2_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i14_LC_2_30_6 (
            .in0(_gnd_net_),
            .in1(N__22465),
            .in2(_gnd_net_),
            .in3(N__22459),
            .lcout(n12_adj_664),
            .ltout(),
            .carryin(n12730),
            .carryout(n12731),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i15_LC_2_30_7.C_ON=1'b1;
    defparam blink_counter_634__i15_LC_2_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i15_LC_2_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i15_LC_2_30_7 (
            .in0(_gnd_net_),
            .in1(N__22597),
            .in2(_gnd_net_),
            .in3(N__22591),
            .lcout(n11_adj_663),
            .ltout(),
            .carryin(n12731),
            .carryout(n12732),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i16_LC_2_31_0.C_ON=1'b1;
    defparam blink_counter_634__i16_LC_2_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i16_LC_2_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i16_LC_2_31_0 (
            .in0(_gnd_net_),
            .in1(N__22588),
            .in2(_gnd_net_),
            .in3(N__22582),
            .lcout(n10_adj_662),
            .ltout(),
            .carryin(bfn_2_31_0_),
            .carryout(n12733),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i17_LC_2_31_1.C_ON=1'b1;
    defparam blink_counter_634__i17_LC_2_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i17_LC_2_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i17_LC_2_31_1 (
            .in0(_gnd_net_),
            .in1(N__22579),
            .in2(_gnd_net_),
            .in3(N__22573),
            .lcout(n9_adj_661),
            .ltout(),
            .carryin(n12733),
            .carryout(n12734),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i18_LC_2_31_2.C_ON=1'b1;
    defparam blink_counter_634__i18_LC_2_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i18_LC_2_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i18_LC_2_31_2 (
            .in0(_gnd_net_),
            .in1(N__22570),
            .in2(_gnd_net_),
            .in3(N__22564),
            .lcout(n8_adj_660),
            .ltout(),
            .carryin(n12734),
            .carryout(n12735),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i19_LC_2_31_3.C_ON=1'b1;
    defparam blink_counter_634__i19_LC_2_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i19_LC_2_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i19_LC_2_31_3 (
            .in0(_gnd_net_),
            .in1(N__22561),
            .in2(_gnd_net_),
            .in3(N__22555),
            .lcout(n7_adj_659),
            .ltout(),
            .carryin(n12735),
            .carryout(n12736),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i20_LC_2_31_4.C_ON=1'b1;
    defparam blink_counter_634__i20_LC_2_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i20_LC_2_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i20_LC_2_31_4 (
            .in0(_gnd_net_),
            .in1(N__22552),
            .in2(_gnd_net_),
            .in3(N__22546),
            .lcout(n6_adj_658),
            .ltout(),
            .carryin(n12736),
            .carryout(n12737),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i21_LC_2_31_5.C_ON=1'b1;
    defparam blink_counter_634__i21_LC_2_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i21_LC_2_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i21_LC_2_31_5 (
            .in0(_gnd_net_),
            .in1(N__36825),
            .in2(_gnd_net_),
            .in3(N__22543),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n12737),
            .carryout(n12738),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i22_LC_2_31_6.C_ON=1'b1;
    defparam blink_counter_634__i22_LC_2_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i22_LC_2_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i22_LC_2_31_6 (
            .in0(_gnd_net_),
            .in1(N__36804),
            .in2(_gnd_net_),
            .in3(N__22540),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n12738),
            .carryout(n12739),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i23_LC_2_31_7.C_ON=1'b1;
    defparam blink_counter_634__i23_LC_2_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i23_LC_2_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i23_LC_2_31_7 (
            .in0(_gnd_net_),
            .in1(N__36783),
            .in2(_gnd_net_),
            .in3(N__22696),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n12739),
            .carryout(n12740),
            .clk(N__56051),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i24_LC_2_32_0.C_ON=1'b1;
    defparam blink_counter_634__i24_LC_2_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i24_LC_2_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i24_LC_2_32_0 (
            .in0(_gnd_net_),
            .in1(N__36843),
            .in2(_gnd_net_),
            .in3(N__22693),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_2_32_0_),
            .carryout(n12741),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_634__i25_LC_2_32_1.C_ON=1'b0;
    defparam blink_counter_634__i25_LC_2_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_634__i25_LC_2_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_634__i25_LC_2_32_1 (
            .in0(_gnd_net_),
            .in1(N__36882),
            .in2(_gnd_net_),
            .in3(N__22690),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i5_4_lut_LC_2_32_5 .C_ON=1'b0;
    defparam \debounce.i5_4_lut_LC_2_32_5 .SEQ_MODE=4'b0000;
    defparam \debounce.i5_4_lut_LC_2_32_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \debounce.i5_4_lut_LC_2_32_5  (
            .in0(N__22687),
            .in1(N__22672),
            .in2(N__22657),
            .in3(N__22636),
            .lcout(\debounce.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i2_LC_2_32_6 .C_ON=1'b0;
    defparam \debounce.reg_B_i2_LC_2_32_6 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i2_LC_2_32_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \debounce.reg_B_i2_LC_2_32_6  (
            .in0(_gnd_net_),
            .in1(N__23907),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(reg_B_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_3_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_3_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_3_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_2_lut_LC_3_17_0 (
            .in0(_gnd_net_),
            .in1(N__37516),
            .in2(_gnd_net_),
            .in3(N__22615),
            .lcout(n2401),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(n12296),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_3_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_3_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_3_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_3_lut_LC_3_17_1 (
            .in0(_gnd_net_),
            .in1(N__53415),
            .in2(N__26533),
            .in3(N__22612),
            .lcout(n2400),
            .ltout(),
            .carryin(n12296),
            .carryout(n12297),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_3_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_3_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_3_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_4_lut_LC_3_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26872),
            .in3(N__22609),
            .lcout(n2399),
            .ltout(),
            .carryin(n12297),
            .carryout(n12298),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_3_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_3_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_3_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_5_lut_LC_3_17_3 (
            .in0(_gnd_net_),
            .in1(N__53416),
            .in2(N__26841),
            .in3(N__22600),
            .lcout(n2398),
            .ltout(),
            .carryin(n12298),
            .carryout(n12299),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_3_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_3_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_3_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_6_lut_LC_3_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24316),
            .in3(N__22723),
            .lcout(n2397),
            .ltout(),
            .carryin(n12299),
            .carryout(n12300),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_3_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_3_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_3_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_7_lut_LC_3_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24054),
            .in3(N__22720),
            .lcout(n2396),
            .ltout(),
            .carryin(n12300),
            .carryout(n12301),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_3_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_3_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_3_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_8_lut_LC_3_17_6 (
            .in0(_gnd_net_),
            .in1(N__53418),
            .in2(N__32394),
            .in3(N__22717),
            .lcout(n2395),
            .ltout(),
            .carryin(n12301),
            .carryout(n12302),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_3_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_3_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_3_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_9_lut_LC_3_17_7 (
            .in0(_gnd_net_),
            .in1(N__53417),
            .in2(N__32362),
            .in3(N__22714),
            .lcout(n2394),
            .ltout(),
            .carryin(n12302),
            .carryout(n12303),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_3_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_3_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_3_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_10_lut_LC_3_18_0 (
            .in0(_gnd_net_),
            .in1(N__53764),
            .in2(N__32302),
            .in3(N__22711),
            .lcout(n2393),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(n12304),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_3_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_3_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_3_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_11_lut_LC_3_18_1 (
            .in0(_gnd_net_),
            .in1(N__53767),
            .in2(N__32278),
            .in3(N__22708),
            .lcout(n2392),
            .ltout(),
            .carryin(n12304),
            .carryout(n12305),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_3_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_3_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_3_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_12_lut_LC_3_18_2 (
            .in0(_gnd_net_),
            .in1(N__53765),
            .in2(N__32425),
            .in3(N__22705),
            .lcout(n2391),
            .ltout(),
            .carryin(n12305),
            .carryout(n12306),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_3_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_3_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_3_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_13_lut_LC_3_18_3 (
            .in0(_gnd_net_),
            .in1(N__53768),
            .in2(N__32245),
            .in3(N__22702),
            .lcout(n2390),
            .ltout(),
            .carryin(n12306),
            .carryout(n12307),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_3_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_3_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_3_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_14_lut_LC_3_18_4 (
            .in0(_gnd_net_),
            .in1(N__53766),
            .in2(N__32335),
            .in3(N__22699),
            .lcout(n2389),
            .ltout(),
            .carryin(n12307),
            .carryout(n12308),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_3_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_3_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_3_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_15_lut_LC_3_18_5 (
            .in0(_gnd_net_),
            .in1(N__53769),
            .in2(N__32455),
            .in3(N__22756),
            .lcout(n2388),
            .ltout(),
            .carryin(n12308),
            .carryout(n12309),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_3_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_3_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_3_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_16_lut_LC_3_18_6 (
            .in0(_gnd_net_),
            .in1(N__32655),
            .in2(N__54248),
            .in3(N__22753),
            .lcout(n2387),
            .ltout(),
            .carryin(n12309),
            .carryout(n12310),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_3_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_3_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_3_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_17_lut_LC_3_18_7 (
            .in0(_gnd_net_),
            .in1(N__53773),
            .in2(N__32640),
            .in3(N__22744),
            .lcout(n2386),
            .ltout(),
            .carryin(n12310),
            .carryout(n12311),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_3_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_3_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_3_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_18_lut_LC_3_19_0 (
            .in0(_gnd_net_),
            .in1(N__24333),
            .in2(N__54249),
            .in3(N__22741),
            .lcout(n2385),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(n12312),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_3_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_3_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_3_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_19_lut_LC_3_19_1 (
            .in0(_gnd_net_),
            .in1(N__24108),
            .in2(N__54252),
            .in3(N__22738),
            .lcout(n2384),
            .ltout(),
            .carryin(n12312),
            .carryout(n12313),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_3_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_3_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_3_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_20_lut_LC_3_19_2 (
            .in0(_gnd_net_),
            .in1(N__39012),
            .in2(N__54250),
            .in3(N__22735),
            .lcout(n2383),
            .ltout(),
            .carryin(n12313),
            .carryout(n12314),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_3_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_3_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_3_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_21_lut_LC_3_19_3 (
            .in0(_gnd_net_),
            .in1(N__29539),
            .in2(N__54253),
            .in3(N__22732),
            .lcout(n2382),
            .ltout(),
            .carryin(n12314),
            .carryout(n12315),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_3_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_3_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_3_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_22_lut_LC_3_19_4 (
            .in0(_gnd_net_),
            .in1(N__26596),
            .in2(N__54251),
            .in3(N__22729),
            .lcout(n2381),
            .ltout(),
            .carryin(n12315),
            .carryout(n12316),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_3_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_3_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_3_19_5.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1570_23_lut_LC_3_19_5 (
            .in0(N__53789),
            .in1(N__34950),
            .in2(N__31921),
            .in3(N__22726),
            .lcout(n2412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_3_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_3_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_3_19_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1386_3_lut_LC_3_19_6 (
            .in0(_gnd_net_),
            .in1(N__22852),
            .in2(N__24453),
            .in3(N__35991),
            .lcout(n2130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_3_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_3_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_3_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1584_3_lut_LC_3_19_7 (
            .in0(_gnd_net_),
            .in1(N__32276),
            .in2(N__22840),
            .in3(N__34906),
            .lcout(n2424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_3_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_3_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_3_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1384_3_lut_LC_3_20_1 (
            .in0(_gnd_net_),
            .in1(N__22831),
            .in2(N__24261),
            .in3(N__35992),
            .lcout(n2128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_3_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_3_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_3_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1453_3_lut_LC_3_20_2 (
            .in0(_gnd_net_),
            .in1(N__26732),
            .in2(N__22822),
            .in3(N__36150),
            .lcout(n2229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_3_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_3_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_3_20_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1316_3_lut_LC_3_20_3 (
            .in0(N__27537),
            .in1(_gnd_net_),
            .in2(N__35894),
            .in3(N__22807),
            .lcout(n2028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_3_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_3_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_3_20_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1452_3_lut_LC_3_20_4 (
            .in0(_gnd_net_),
            .in1(N__26762),
            .in2(N__22801),
            .in3(N__36149),
            .lcout(n2228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_20_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1457_3_lut_LC_3_20_5 (
            .in0(_gnd_net_),
            .in1(N__27993),
            .in2(N__36191),
            .in3(N__22786),
            .lcout(n2233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_95_LC_3_20_6.C_ON=1'b0;
    defparam i1_4_lut_adj_95_LC_3_20_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_95_LC_3_20_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_95_LC_3_20_6 (
            .in0(N__29705),
            .in1(N__27635),
            .in2(N__22890),
            .in3(N__24208),
            .lcout(n14160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_3_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_3_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_3_20_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1442_3_lut_LC_3_20_7 (
            .in0(_gnd_net_),
            .in1(N__22768),
            .in2(N__36192),
            .in3(N__27053),
            .lcout(n2218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_92_LC_3_21_0.C_ON=1'b0;
    defparam i1_4_lut_adj_92_LC_3_21_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_92_LC_3_21_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_92_LC_3_21_0 (
            .in0(N__24644),
            .in1(N__29615),
            .in2(N__22976),
            .in3(N__23021),
            .lcout(n14146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_3_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_3_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_3_21_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1309_3_lut_LC_3_21_1 (
            .in0(_gnd_net_),
            .in1(N__24766),
            .in2(N__23005),
            .in3(N__35863),
            .lcout(n2021),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_3_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_3_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_3_21_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1318_3_lut_LC_3_21_2 (
            .in0(N__22996),
            .in1(_gnd_net_),
            .in2(N__35888),
            .in3(N__26904),
            .lcout(n2030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_3_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_3_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_3_21_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1314_3_lut_LC_3_21_3 (
            .in0(N__24798),
            .in1(_gnd_net_),
            .in2(N__22990),
            .in3(N__35858),
            .lcout(n2026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_3_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_3_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_3_21_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 encoder0_position_31__I_0_i1239_3_lut_LC_3_21_4 (
            .in0(N__35747),
            .in1(N__22951),
            .in2(_gnd_net_),
            .in3(N__23194),
            .lcout(n1919),
            .ltout(n1919_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_3_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_3_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_3_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1306_3_lut_LC_3_21_5 (
            .in0(_gnd_net_),
            .in1(N__22939),
            .in2(N__22933),
            .in3(N__35867),
            .lcout(n2018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_3_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_3_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_3_21_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1308_3_lut_LC_3_21_6 (
            .in0(N__26974),
            .in1(_gnd_net_),
            .in2(N__35889),
            .in3(N__22900),
            .lcout(n2020),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_3_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_3_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_3_21_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1307_3_lut_LC_3_21_7 (
            .in0(_gnd_net_),
            .in1(N__24733),
            .in2(N__22867),
            .in3(N__35862),
            .lcout(n2019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_3_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_3_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_3_22_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1311_3_lut_LC_3_22_0 (
            .in0(_gnd_net_),
            .in1(N__22858),
            .in2(N__23113),
            .in3(N__35875),
            .lcout(n2023),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_3_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_3_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_3_22_1.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i1244_3_lut_LC_3_22_1 (
            .in0(N__35727),
            .in1(N__27859),
            .in2(N__23128),
            .in3(_gnd_net_),
            .lcout(n1924),
            .ltout(n1924_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_87_LC_3_22_2.C_ON=1'b0;
    defparam i1_3_lut_adj_87_LC_3_22_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_87_LC_3_22_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_87_LC_3_22_2 (
            .in0(_gnd_net_),
            .in1(N__24794),
            .in2(N__23095),
            .in3(N__24401),
            .lcout(n13770),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_3_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_3_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_3_22_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1245_3_lut_LC_3_22_3 (
            .in0(_gnd_net_),
            .in1(N__27801),
            .in2(N__35752),
            .in3(N__23092),
            .lcout(n1925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_3_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_3_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_3_22_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1243_3_lut_LC_3_22_4 (
            .in0(N__27306),
            .in1(_gnd_net_),
            .in2(N__23080),
            .in3(N__35726),
            .lcout(n1923),
            .ltout(n1923_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_88_LC_3_22_5.C_ON=1'b0;
    defparam i1_3_lut_adj_88_LC_3_22_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_88_LC_3_22_5.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_88_LC_3_22_5 (
            .in0(_gnd_net_),
            .in1(N__24494),
            .in2(N__23065),
            .in3(N__24686),
            .lcout(n13772),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_3_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_3_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_3_22_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1248_3_lut_LC_3_22_7 (
            .in0(N__35725),
            .in1(_gnd_net_),
            .in2(N__23062),
            .in3(N__27236),
            .lcout(n1928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_3_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_3_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_3_23_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1251_3_lut_LC_3_23_0 (
            .in0(_gnd_net_),
            .in1(N__23047),
            .in2(N__27712),
            .in3(N__35721),
            .lcout(n1931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_3_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_3_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_3_23_2.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1174_3_lut_LC_3_23_2 (
            .in0(N__25189),
            .in1(N__25211),
            .in2(N__35622),
            .in3(_gnd_net_),
            .lcout(n1822),
            .ltout(n1822_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_86_LC_3_23_3.C_ON=1'b0;
    defparam i1_3_lut_adj_86_LC_3_23_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_86_LC_3_23_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_86_LC_3_23_3 (
            .in0(_gnd_net_),
            .in1(N__23150),
            .in2(N__23038),
            .in3(N__23180),
            .lcout(n14134),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_3_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_3_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_3_23_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1246_3_lut_LC_3_23_4 (
            .in0(_gnd_net_),
            .in1(N__23218),
            .in2(N__27835),
            .in3(N__35720),
            .lcout(n1926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12540_1_lut_LC_3_23_5.C_ON=1'b0;
    defparam i12540_1_lut_LC_3_23_5.SEQ_MODE=4'b0000;
    defparam i12540_1_lut_LC_3_23_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12540_1_lut_LC_3_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35890),
            .in3(_gnd_net_),
            .lcout(n15012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_3_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_3_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_3_23_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1104_3_lut_LC_3_23_6 (
            .in0(N__35487),
            .in1(_gnd_net_),
            .in2(N__23539),
            .in3(N__23209),
            .lcout(n1720),
            .ltout(n1720_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_3_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_3_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_3_23_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1171_3_lut_LC_3_23_7 (
            .in0(_gnd_net_),
            .in1(N__35600),
            .in2(N__23197),
            .in3(N__25096),
            .lcout(n1819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12497_1_lut_LC_3_24_0.C_ON=1'b0;
    defparam i12497_1_lut_LC_3_24_0.SEQ_MODE=4'b0000;
    defparam i12497_1_lut_LC_3_24_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12497_1_lut_LC_3_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35595),
            .lcout(n14969),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_3_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_3_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_3_24_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1172_3_lut_LC_3_24_1 (
            .in0(N__25134),
            .in1(_gnd_net_),
            .in2(N__35621),
            .in3(N__25120),
            .lcout(n1820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12500_4_lut_LC_3_24_2.C_ON=1'b0;
    defparam i12500_4_lut_LC_3_24_2.SEQ_MODE=4'b0000;
    defparam i12500_4_lut_LC_3_24_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12500_4_lut_LC_3_24_2 (
            .in0(N__25107),
            .in1(N__25133),
            .in2(N__23311),
            .in3(N__25080),
            .lcout(n1752),
            .ltout(n1752_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_3_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_3_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_3_24_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1176_3_lut_LC_3_24_3 (
            .in0(N__25245),
            .in1(_gnd_net_),
            .in2(N__23164),
            .in3(N__25225),
            .lcout(n1824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_3_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_3_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_3_24_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i1173_3_lut_LC_3_24_4 (
            .in0(_gnd_net_),
            .in1(N__35599),
            .in2(N__25153),
            .in3(N__25173),
            .lcout(n1821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_149_LC_3_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_149_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_149_LC_3_24_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_149_LC_3_24_5 (
            .in0(N__23266),
            .in1(N__23388),
            .in2(N__23253),
            .in3(N__23134),
            .lcout(),
            .ltout(n14110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12480_4_lut_LC_3_24_6.C_ON=1'b0;
    defparam i12480_4_lut_LC_3_24_6.SEQ_MODE=4'b0000;
    defparam i12480_4_lut_LC_3_24_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12480_4_lut_LC_3_24_6 (
            .in0(N__25638),
            .in1(N__23603),
            .in2(N__23350),
            .in3(N__23531),
            .lcout(n1653),
            .ltout(n1653_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_3_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_3_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_3_24_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1107_3_lut_LC_3_24_7 (
            .in0(N__23249),
            .in1(_gnd_net_),
            .in2(N__23347),
            .in3(N__23344),
            .lcout(n1723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_80_LC_3_25_0.C_ON=1'b0;
    defparam i1_4_lut_adj_80_LC_3_25_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_80_LC_3_25_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_80_LC_3_25_0 (
            .in0(N__25241),
            .in1(N__27341),
            .in2(N__25212),
            .in3(N__23332),
            .lcout(),
            .ltout(n13968_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_82_LC_3_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_82_LC_3_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_82_LC_3_25_1.LUT_INIT=16'b1111111011111010;
    LogicCell40 i1_4_lut_adj_82_LC_3_25_1 (
            .in0(N__25169),
            .in1(N__23326),
            .in2(N__23320),
            .in3(N__23317),
            .lcout(n13972),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_3_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_3_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_3_25_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_i1106_3_lut_LC_3_25_2 (
            .in0(N__23387),
            .in1(N__35486),
            .in2(_gnd_net_),
            .in3(N__23302),
            .lcout(n1722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_147_LC_3_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_147_LC_3_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_147_LC_3_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_147_LC_3_25_3 (
            .in0(N__23501),
            .in1(N__23282),
            .in2(N__23664),
            .in3(N__23408),
            .lcout(n14104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_3_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_3_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_3_25_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1040_3_lut_LC_3_25_4 (
            .in0(N__25555),
            .in1(_gnd_net_),
            .in2(N__25759),
            .in3(N__35382),
            .lcout(n1624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_3_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_3_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_3_25_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1108_3_lut_LC_3_25_5 (
            .in0(N__35484),
            .in1(_gnd_net_),
            .in2(N__23233),
            .in3(N__23409),
            .lcout(n1724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_3_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_3_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_3_25_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1109_3_lut_LC_3_25_6 (
            .in0(_gnd_net_),
            .in1(N__23502),
            .in2(N__23488),
            .in3(N__35485),
            .lcout(n1725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_3_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_3_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_3_25_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_3_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29897),
            .lcout(n13_adj_637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_3_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_3_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_3_26_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1048_3_lut_LC_3_26_0 (
            .in0(N__25488),
            .in1(_gnd_net_),
            .in2(N__25474),
            .in3(N__35373),
            .lcout(n1632),
            .ltout(n1632_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9920_3_lut_LC_3_26_1.C_ON=1'b0;
    defparam i9920_3_lut_LC_3_26_1.SEQ_MODE=4'b0000;
    defparam i9920_3_lut_LC_3_26_1.LUT_INIT=16'b1111000010100000;
    LogicCell40 i9920_3_lut_LC_3_26_1 (
            .in0(N__28097),
            .in1(_gnd_net_),
            .in2(N__23452),
            .in3(N__23441),
            .lcout(n11634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_3_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_3_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_3_26_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1041_3_lut_LC_3_26_2 (
            .in0(_gnd_net_),
            .in1(N__25255),
            .in2(N__25591),
            .in3(N__35378),
            .lcout(n1625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_3_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_3_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_3_26_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1039_3_lut_LC_3_26_3 (
            .in0(_gnd_net_),
            .in1(N__25810),
            .in2(N__35391),
            .in3(N__25741),
            .lcout(n1623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12820_1_lut_LC_3_26_4.C_ON=1'b0;
    defparam i12820_1_lut_LC_3_26_4.SEQ_MODE=4'b0000;
    defparam i12820_1_lut_LC_3_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12820_1_lut_LC_3_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35374),
            .lcout(n15292),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i979_3_lut_LC_3_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_3_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_3_26_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i979_3_lut_LC_3_26_5 (
            .in0(_gnd_net_),
            .in1(N__23743),
            .in2(N__23368),
            .in3(N__35282),
            .lcout(n1531),
            .ltout(n1531_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9983_4_lut_LC_3_26_6.C_ON=1'b0;
    defparam i9983_4_lut_LC_3_26_6.SEQ_MODE=4'b0000;
    defparam i9983_4_lut_LC_3_26_6.LUT_INIT=16'b1111111011110000;
    LogicCell40 i9983_4_lut_LC_3_26_6 (
            .in0(N__25487),
            .in1(N__27570),
            .in2(N__23359),
            .in3(N__25454),
            .lcout(n11698),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_3_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_3_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1043_3_lut_LC_3_26_7.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1043_3_lut_LC_3_26_7 (
            .in0(N__25306),
            .in1(N__25323),
            .in2(N__35390),
            .in3(_gnd_net_),
            .lcout(n1627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i977_3_lut_LC_3_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_3_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_3_27_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i977_3_lut_LC_3_27_0 (
            .in0(N__23641),
            .in1(N__23623),
            .in2(N__35279),
            .in3(_gnd_net_),
            .lcout(n1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_3_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_3_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_3_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_3_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29928),
            .lcout(n14_adj_638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i978_3_lut_LC_3_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_3_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_3_27_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i978_3_lut_LC_3_27_2 (
            .in0(_gnd_net_),
            .in1(N__23617),
            .in2(N__35280),
            .in3(N__25934),
            .lcout(n1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_3_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_3_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_3_27_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1038_3_lut_LC_3_27_3 (
            .in0(_gnd_net_),
            .in1(N__25724),
            .in2(N__25702),
            .in3(N__35384),
            .lcout(n1622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_3_27_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_3_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_3_27_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i20_3_lut_LC_3_27_4 (
            .in0(N__29929),
            .in1(N__33271),
            .in2(_gnd_net_),
            .in3(N__39546),
            .lcout(n300),
            .ltout(n300_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i981_3_lut_LC_3_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_3_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_3_27_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i981_3_lut_LC_3_27_5 (
            .in0(_gnd_net_),
            .in1(N__23560),
            .in2(N__23554),
            .in3(N__35258),
            .lcout(n1533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i970_3_lut_LC_3_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_3_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_3_27_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i970_3_lut_LC_3_27_6 (
            .in0(_gnd_net_),
            .in1(N__25896),
            .in2(N__35281),
            .in3(N__23551),
            .lcout(n1522),
            .ltout(n1522_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_3_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_3_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_3_27_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1037_3_lut_LC_3_27_7 (
            .in0(_gnd_net_),
            .in1(N__25678),
            .in2(N__23542),
            .in3(N__35383),
            .lcout(n1621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i975_3_lut_LC_3_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_3_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_3_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i975_3_lut_LC_3_28_0 (
            .in0(_gnd_net_),
            .in1(N__25514),
            .in2(N__23773),
            .in3(N__35246),
            .lcout(n1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i976_3_lut_LC_3_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i976_3_lut_LC_3_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i976_3_lut_LC_3_28_1.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i976_3_lut_LC_3_28_1 (
            .in0(N__26054),
            .in1(N__23764),
            .in2(N__35274),
            .in3(_gnd_net_),
            .lcout(n1528),
            .ltout(n1528_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_78_LC_3_28_2.C_ON=1'b0;
    defparam i1_2_lut_adj_78_LC_3_28_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_78_LC_3_28_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_78_LC_3_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23758),
            .in3(N__25286),
            .lcout(),
            .ltout(n13978_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_126_LC_3_28_3.C_ON=1'b0;
    defparam i1_4_lut_adj_126_LC_3_28_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_126_LC_3_28_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_126_LC_3_28_3 (
            .in0(N__25544),
            .in1(N__25802),
            .in2(N__23755),
            .in3(N__25583),
            .lcout(n13984),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i912_3_lut_LC_3_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_3_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_3_28_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i912_3_lut_LC_3_28_4 (
            .in0(N__25776),
            .in1(_gnd_net_),
            .in2(N__23833),
            .in3(N__36720),
            .lcout(n1432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_75_LC_3_28_5.C_ON=1'b0;
    defparam i1_4_lut_adj_75_LC_3_28_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_75_LC_3_28_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_75_LC_3_28_5 (
            .in0(N__26121),
            .in1(N__25964),
            .in2(N__25845),
            .in3(N__23716),
            .lcout(n14094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i913_3_lut_LC_3_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_3_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_3_28_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i913_3_lut_LC_3_28_6 (
            .in0(N__23677),
            .in1(N__26110),
            .in2(_gnd_net_),
            .in3(N__36721),
            .lcout(n1433),
            .ltout(n1433_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i980_3_lut_LC_3_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_3_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_3_28_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i980_3_lut_LC_3_28_7 (
            .in0(N__35247),
            .in1(_gnd_net_),
            .in2(N__23686),
            .in3(N__23683),
            .lcout(n1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_3_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_3_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_3_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_2_lut_LC_3_29_0 (
            .in0(_gnd_net_),
            .in1(N__26109),
            .in2(_gnd_net_),
            .in3(N__23671),
            .lcout(n1401),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(n12141),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_3_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_3_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_3_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_3_lut_LC_3_29_1 (
            .in0(_gnd_net_),
            .in1(N__54738),
            .in2(N__25777),
            .in3(N__23824),
            .lcout(n1400),
            .ltout(),
            .carryin(n12141),
            .carryout(n12142),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_3_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_3_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_3_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_4_lut_LC_3_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26307),
            .in3(N__23821),
            .lcout(n1399),
            .ltout(),
            .carryin(n12142),
            .carryout(n12143),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_3_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_3_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_3_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_5_lut_LC_3_29_3 (
            .in0(_gnd_net_),
            .in1(N__54739),
            .in2(N__26187),
            .in3(N__23806),
            .lcout(n1398),
            .ltout(),
            .carryin(n12143),
            .carryout(n12144),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_3_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_3_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_3_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_6_lut_LC_3_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26092),
            .in3(N__23803),
            .lcout(n1397),
            .ltout(),
            .carryin(n12144),
            .carryout(n12145),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_3_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_3_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_3_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_7_lut_LC_3_29_5 (
            .in0(_gnd_net_),
            .in1(N__26019),
            .in2(_gnd_net_),
            .in3(N__23800),
            .lcout(n1396),
            .ltout(),
            .carryin(n12145),
            .carryout(n12146),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_3_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_3_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_3_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_8_lut_LC_3_29_6 (
            .in0(_gnd_net_),
            .in1(N__54741),
            .in2(N__28329),
            .in3(N__23785),
            .lcout(n1395),
            .ltout(),
            .carryin(n12146),
            .carryout(n12147),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_3_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_3_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_3_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_9_lut_LC_3_29_7 (
            .in0(_gnd_net_),
            .in1(N__54740),
            .in2(N__28362),
            .in3(N__23782),
            .lcout(n1394),
            .ltout(),
            .carryin(n12147),
            .carryout(n12148),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_3_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_3_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_3_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_10_lut_LC_3_30_0 (
            .in0(_gnd_net_),
            .in1(N__55070),
            .in2(N__28389),
            .in3(N__23779),
            .lcout(n1393),
            .ltout(),
            .carryin(bfn_3_30_0_),
            .carryout(n12149),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_3_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_3_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_3_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_11_lut_LC_3_30_1 (
            .in0(_gnd_net_),
            .in1(N__55072),
            .in2(N__28408),
            .in3(N__23776),
            .lcout(n1392),
            .ltout(),
            .carryin(n12149),
            .carryout(n12150),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_3_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_3_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_12_lut_LC_3_30_2 (
            .in0(_gnd_net_),
            .in1(N__26216),
            .in2(N__55209),
            .in3(N__23866),
            .lcout(n1391),
            .ltout(),
            .carryin(n12150),
            .carryout(n12151),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_3_30_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_3_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_3_30_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_900_13_lut_LC_3_30_3 (
            .in0(N__55071),
            .in1(N__36756),
            .in2(N__26164),
            .in3(N__23863),
            .lcout(n1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i842_3_lut_LC_3_30_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_3_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_3_30_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i842_3_lut_LC_3_30_5 (
            .in0(_gnd_net_),
            .in1(N__23842),
            .in2(N__28516),
            .in3(N__36629),
            .lcout(n1330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i2_4_lut_adj_26_LC_3_30_6 .C_ON=1'b0;
    defparam \debounce.i2_4_lut_adj_26_LC_3_30_6 .SEQ_MODE=4'b0000;
    defparam \debounce.i2_4_lut_adj_26_LC_3_30_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \debounce.i2_4_lut_adj_26_LC_3_30_6  (
            .in0(N__28143),
            .in1(N__28119),
            .in2(N__28450),
            .in3(N__28473),
            .lcout(\debounce.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i843_3_lut_LC_3_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_3_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_3_30_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i843_3_lut_LC_3_30_7 (
            .in0(_gnd_net_),
            .in1(N__28263),
            .in2(N__23854),
            .in3(N__36628),
            .lcout(n1331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_3_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_3_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_3_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_2_lut_LC_3_31_0 (
            .in0(_gnd_net_),
            .in1(N__28300),
            .in2(_gnd_net_),
            .in3(N__23860),
            .lcout(n1301),
            .ltout(),
            .carryin(bfn_3_31_0_),
            .carryout(n12131),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_3_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_3_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_3_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_3_lut_LC_3_31_1 (
            .in0(_gnd_net_),
            .in1(N__55063),
            .in2(N__28282),
            .in3(N__23857),
            .lcout(n1300),
            .ltout(),
            .carryin(n12131),
            .carryout(n12132),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_3_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_3_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_3_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_4_lut_LC_3_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28264),
            .in3(N__23845),
            .lcout(n1299),
            .ltout(),
            .carryin(n12132),
            .carryout(n12133),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_3_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_3_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_3_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_5_lut_LC_3_31_3 (
            .in0(_gnd_net_),
            .in1(N__55064),
            .in2(N__28515),
            .in3(N__23836),
            .lcout(n1298),
            .ltout(),
            .carryin(n12133),
            .carryout(n12134),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_3_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_3_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_3_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_6_lut_LC_3_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28558),
            .in3(N__23947),
            .lcout(n1297),
            .ltout(),
            .carryin(n12134),
            .carryout(n12135),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_3_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_3_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_3_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_7_lut_LC_3_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28537),
            .in3(N__23944),
            .lcout(n1296),
            .ltout(),
            .carryin(n12135),
            .carryout(n12136),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_3_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_3_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_3_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_8_lut_LC_3_31_6 (
            .in0(_gnd_net_),
            .in1(N__55066),
            .in2(N__28231),
            .in3(N__23941),
            .lcout(n1295),
            .ltout(),
            .carryin(n12136),
            .carryout(n12137),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_3_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_3_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_3_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_9_lut_LC_3_31_7 (
            .in0(_gnd_net_),
            .in1(N__55065),
            .in2(N__28594),
            .in3(N__23938),
            .lcout(n1294),
            .ltout(),
            .carryin(n12137),
            .carryout(n12138),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_3_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_3_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_3_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_10_lut_LC_3_32_0 (
            .in0(_gnd_net_),
            .in1(N__55067),
            .in2(N__28714),
            .in3(N__23935),
            .lcout(n1293),
            .ltout(),
            .carryin(bfn_3_32_0_),
            .carryout(n12139),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_3_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_3_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_3_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_11_lut_LC_3_32_1 (
            .in0(_gnd_net_),
            .in1(N__55068),
            .in2(N__26256),
            .in3(N__23932),
            .lcout(n1292),
            .ltout(),
            .carryin(n12139),
            .carryout(n12140),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_3_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_3_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_3_32_2.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_833_12_lut_LC_3_32_2 (
            .in0(N__55069),
            .in1(N__36663),
            .in2(N__26353),
            .in3(N__23929),
            .lcout(n1323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i2_LC_3_32_3 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i2_LC_3_32_3 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i2_LC_3_32_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \debounce.reg_out_i0_i2_LC_3_32_3  (
            .in0(N__27944),
            .in1(N__23926),
            .in2(_gnd_net_),
            .in3(N__38070),
            .lcout(h1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56057),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i3_4_lut_LC_3_32_4 .C_ON=1'b0;
    defparam \debounce.i3_4_lut_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \debounce.i3_4_lut_LC_3_32_4 .LUT_INIT=16'b1101111011111111;
    LogicCell40 \debounce.i3_4_lut_LC_3_32_4  (
            .in0(N__23925),
            .in1(N__23917),
            .in2(N__23908),
            .in3(N__27943),
            .lcout(\debounce.cnt_next_9__N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i769_3_lut_LC_3_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_3_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_3_32_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i769_3_lut_LC_3_32_7 (
            .in0(_gnd_net_),
            .in1(N__36541),
            .in2(N__28789),
            .in3(N__24010),
            .lcout(n1225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_104_LC_4_17_0.C_ON=1'b0;
    defparam i1_2_lut_adj_104_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_104_LC_4_17_0.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_104_LC_4_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31395),
            .in3(N__31358),
            .lcout(n14410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_4_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_4_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_4_17_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1454_3_lut_LC_4_17_1 (
            .in0(_gnd_net_),
            .in1(N__24001),
            .in2(N__36207),
            .in3(N__26709),
            .lcout(n2230),
            .ltout(n2230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_4_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_4_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_4_17_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1521_3_lut_LC_4_17_2 (
            .in0(N__39133),
            .in1(_gnd_net_),
            .in2(N__23992),
            .in3(N__31378),
            .lcout(n2329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_4_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_4_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_4_17_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1656_3_lut_LC_4_17_3 (
            .in0(_gnd_net_),
            .in1(N__28960),
            .in2(N__28980),
            .in3(N__35046),
            .lcout(n2528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_17_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1445_3_lut_LC_4_17_4 (
            .in0(_gnd_net_),
            .in1(N__24588),
            .in2(N__23989),
            .in3(N__36194),
            .lcout(n2221),
            .ltout(n2221_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_4_17_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1512_3_lut_LC_4_17_5 (
            .in0(_gnd_net_),
            .in1(N__31678),
            .in2(N__23974),
            .in3(N__39132),
            .lcout(n2320),
            .ltout(n2320_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_17_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1579_3_lut_LC_4_17_6 (
            .in0(N__34925),
            .in1(_gnd_net_),
            .in2(N__23971),
            .in3(N__23968),
            .lcout(n2419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_4_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_4_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_4_17_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1591_3_lut_LC_4_17_7 (
            .in0(_gnd_net_),
            .in1(N__26871),
            .in2(N__23962),
            .in3(N__34924),
            .lcout(n2431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_4_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_4_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_4_18_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1589_3_lut_LC_4_18_0 (
            .in0(_gnd_net_),
            .in1(N__23953),
            .in2(N__34927),
            .in3(N__24312),
            .lcout(n2429),
            .ltout(n2429_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_114_LC_4_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_114_LC_4_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_114_LC_4_18_1.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_114_LC_4_18_1 (
            .in0(N__29411),
            .in1(N__29018),
            .in2(N__24076),
            .in3(N__26461),
            .lcout(n13423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_112_LC_4_18_2.C_ON=1'b0;
    defparam i1_4_lut_adj_112_LC_4_18_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_112_LC_4_18_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_112_LC_4_18_2 (
            .in0(N__28937),
            .in1(N__30884),
            .in2(N__31239),
            .in3(N__31292),
            .lcout(),
            .ltout(n14210_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_113_LC_4_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_113_LC_4_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_113_LC_4_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_113_LC_4_18_3 (
            .in0(N__30681),
            .in1(N__28895),
            .in2(N__24073),
            .in3(N__29207),
            .lcout(),
            .ltout(n14214_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_115_LC_4_18_4.C_ON=1'b0;
    defparam i1_4_lut_adj_115_LC_4_18_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_115_LC_4_18_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_115_LC_4_18_4 (
            .in0(N__31138),
            .in1(N__31019),
            .in2(N__24070),
            .in3(N__24067),
            .lcout(n14220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_18_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1588_3_lut_LC_4_18_5 (
            .in0(_gnd_net_),
            .in1(N__24061),
            .in2(N__24055),
            .in3(N__34896),
            .lcout(n2428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_110_LC_4_19_0.C_ON=1'b0;
    defparam i1_4_lut_adj_110_LC_4_19_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_110_LC_4_19_0.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_110_LC_4_19_0 (
            .in0(N__24308),
            .in1(N__24053),
            .in2(N__26821),
            .in3(N__32605),
            .lcout(),
            .ltout(n14016_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_111_LC_4_19_1.C_ON=1'b0;
    defparam i1_4_lut_adj_111_LC_4_19_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_111_LC_4_19_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_111_LC_4_19_1 (
            .in0(N__24329),
            .in1(N__24104),
            .in2(N__24028),
            .in3(N__39011),
            .lcout(),
            .ltout(n14022_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12879_4_lut_LC_4_19_2.C_ON=1'b0;
    defparam i12879_4_lut_LC_4_19_2.SEQ_MODE=4'b0000;
    defparam i12879_4_lut_LC_4_19_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12879_4_lut_LC_4_19_2 (
            .in0(N__26592),
            .in1(N__29538),
            .in2(N__24025),
            .in3(N__31917),
            .lcout(n2346),
            .ltout(n2346_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_19_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1587_3_lut_LC_4_19_3 (
            .in0(_gnd_net_),
            .in1(N__24022),
            .in2(N__24013),
            .in3(N__32384),
            .lcout(n2427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_4_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_4_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_4_19_4.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1576_3_lut_LC_4_19_4 (
            .in0(N__34905),
            .in1(N__24127),
            .in2(N__24109),
            .in3(_gnd_net_),
            .lcout(n2416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_4_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_4_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_4_19_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1577_3_lut_LC_4_19_5 (
            .in0(N__24121),
            .in1(_gnd_net_),
            .in2(N__24334),
            .in3(N__34904),
            .lcout(n2417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_4_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_4_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_4_19_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1581_3_lut_LC_4_19_6 (
            .in0(_gnd_net_),
            .in1(N__24115),
            .in2(N__34928),
            .in3(N__32334),
            .lcout(n2421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12876_1_lut_LC_4_19_7.C_ON=1'b0;
    defparam i12876_1_lut_LC_4_19_7.SEQ_MODE=4'b0000;
    defparam i12876_1_lut_LC_4_19_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12876_1_lut_LC_4_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34900),
            .lcout(n15348),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_20_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1509_3_lut_LC_4_20_0 (
            .in0(_gnd_net_),
            .in1(N__32088),
            .in2(N__32074),
            .in3(N__39072),
            .lcout(n2317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10059_4_lut_LC_4_20_1.C_ON=1'b0;
    defparam i10059_4_lut_LC_4_20_1.SEQ_MODE=4'b0000;
    defparam i10059_4_lut_LC_4_20_1.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10059_4_lut_LC_4_20_1 (
            .in0(N__31517),
            .in1(N__32160),
            .in2(N__31437),
            .in3(N__31476),
            .lcout(),
            .ltout(n11774_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_105_LC_4_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_105_LC_4_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_105_LC_4_20_2.LUT_INIT=16'b1111111111101010;
    LogicCell40 i1_4_lut_adj_105_LC_4_20_2 (
            .in0(N__31659),
            .in1(N__24091),
            .in2(N__24082),
            .in3(N__29464),
            .lcout(),
            .ltout(n14188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_106_LC_4_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_106_LC_4_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_106_LC_4_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_106_LC_4_20_3 (
            .in0(N__32087),
            .in1(N__32121),
            .in2(N__24079),
            .in3(N__39179),
            .lcout(n14194),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_4_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_4_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_4_20_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1520_3_lut_LC_4_20_4 (
            .in0(N__31333),
            .in1(_gnd_net_),
            .in2(N__31362),
            .in3(N__39067),
            .lcout(n2328),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_4_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_4_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_4_20_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1443_3_lut_LC_4_20_5 (
            .in0(_gnd_net_),
            .in1(N__24349),
            .in2(N__36206),
            .in3(N__27606),
            .lcout(n2219),
            .ltout(n2219_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_4_20_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1510_3_lut_LC_4_20_6 (
            .in0(N__32110),
            .in1(_gnd_net_),
            .in2(N__24337),
            .in3(N__39071),
            .lcout(n2318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_4_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_4_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_4_20_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1522_3_lut_LC_4_20_7 (
            .in0(N__31433),
            .in1(_gnd_net_),
            .in2(N__39105),
            .in3(N__31414),
            .lcout(n2330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_4_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_4_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_4_21_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1387_3_lut_LC_4_21_0 (
            .in0(N__24289),
            .in1(_gnd_net_),
            .in2(N__27180),
            .in3(N__36031),
            .lcout(n2131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_4_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_4_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_4_21_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i1317_3_lut_LC_4_21_1 (
            .in0(_gnd_net_),
            .in1(N__35870),
            .in2(N__24277),
            .in3(N__27453),
            .lcout(n2029),
            .ltout(n2029_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_94_LC_4_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_94_LC_4_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_94_LC_4_21_2.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_94_LC_4_21_2 (
            .in0(N__24224),
            .in1(N__24424),
            .in2(N__24211),
            .in3(N__24133),
            .lcout(n14154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_4_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_4_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_4_21_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i1310_3_lut_LC_4_21_3 (
            .in0(_gnd_net_),
            .in1(N__35869),
            .in2(N__24202),
            .in3(N__24187),
            .lcout(n2022),
            .ltout(n2022_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_93_LC_4_21_4.C_ON=1'b0;
    defparam i1_4_lut_adj_93_LC_4_21_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_93_LC_4_21_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_93_LC_4_21_4 (
            .in0(N__27128),
            .in1(N__24620),
            .in2(N__24142),
            .in3(N__24139),
            .lcout(n14152),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_4_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_4_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_4_21_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1315_3_lut_LC_4_21_5 (
            .in0(_gnd_net_),
            .in1(N__35868),
            .in2(N__24694),
            .in3(N__24670),
            .lcout(n2027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_4_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_4_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_4_21_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1378_3_lut_LC_4_21_6 (
            .in0(N__24624),
            .in1(_gnd_net_),
            .in2(N__24604),
            .in3(N__36032),
            .lcout(n2122),
            .ltout(n2122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_97_LC_4_21_7.C_ON=1'b0;
    defparam i1_3_lut_adj_97_LC_4_21_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_97_LC_4_21_7.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_97_LC_4_21_7 (
            .in0(N__24557),
            .in1(_gnd_net_),
            .in2(N__24541),
            .in3(N__29505),
            .lcout(n13748),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12543_4_lut_LC_4_22_0.C_ON=1'b0;
    defparam i12543_4_lut_LC_4_22_0.SEQ_MODE=4'b0000;
    defparam i12543_4_lut_LC_4_22_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12543_4_lut_LC_4_22_0 (
            .in0(N__24538),
            .in1(N__27372),
            .in2(N__24514),
            .in3(N__24703),
            .lcout(n1950),
            .ltout(n1950_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_4_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_4_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_4_22_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1313_3_lut_LC_4_22_1 (
            .in0(N__24498),
            .in1(_gnd_net_),
            .in2(N__24478),
            .in3(N__24475),
            .lcout(n2025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_4_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_4_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_4_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1319_3_lut_LC_4_22_2 (
            .in0(_gnd_net_),
            .in1(N__24466),
            .in2(N__26931),
            .in3(N__35874),
            .lcout(n2031),
            .ltout(n2031_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9965_4_lut_LC_4_22_3.C_ON=1'b0;
    defparam i9965_4_lut_LC_4_22_3.SEQ_MODE=4'b0000;
    defparam i9965_4_lut_LC_4_22_3.LUT_INIT=16'b1111101011111000;
    LogicCell40 i9965_4_lut_LC_4_22_3 (
            .in0(N__27164),
            .in1(N__26661),
            .in2(N__24427),
            .in3(N__27914),
            .lcout(n11680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_4_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_4_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_4_22_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1312_3_lut_LC_4_22_4 (
            .in0(_gnd_net_),
            .in1(N__24418),
            .in2(N__24409),
            .in3(N__35873),
            .lcout(n2024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12521_4_lut_LC_4_22_6.C_ON=1'b0;
    defparam i12521_4_lut_LC_4_22_6.SEQ_MODE=4'b0000;
    defparam i12521_4_lut_LC_4_22_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12521_4_lut_LC_4_22_6 (
            .in0(N__24378),
            .in1(N__24355),
            .in2(N__27211),
            .in3(N__27413),
            .lcout(n1851),
            .ltout(n1851_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_4_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_4_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_4_22_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1247_3_lut_LC_4_22_7 (
            .in0(N__27741),
            .in1(_gnd_net_),
            .in2(N__24820),
            .in3(N__24817),
            .lcout(n1927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_4_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_4_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_4_23_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1181_3_lut_LC_4_23_0 (
            .in0(_gnd_net_),
            .in1(N__24916),
            .in2(N__24946),
            .in3(N__35620),
            .lcout(n1829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_4_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_4_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_4_23_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1242_3_lut_LC_4_23_2 (
            .in0(N__27324),
            .in1(_gnd_net_),
            .in2(N__35761),
            .in3(N__24778),
            .lcout(n1922),
            .ltout(n1922_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_89_LC_4_23_3.C_ON=1'b0;
    defparam i1_4_lut_adj_89_LC_4_23_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_89_LC_4_23_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_89_LC_4_23_3 (
            .in0(N__26960),
            .in1(N__24748),
            .in2(N__24742),
            .in3(N__24739),
            .lcout(),
            .ltout(n13778_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_91_LC_4_23_4.C_ON=1'b0;
    defparam i1_4_lut_adj_91_LC_4_23_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_91_LC_4_23_4.LUT_INIT=16'b1111111011111100;
    LogicCell40 i1_4_lut_adj_91_LC_4_23_4 (
            .in0(N__27508),
            .in1(N__24729),
            .in2(N__24706),
            .in3(N__26878),
            .lcout(n13782),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_4_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_4_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_4_23_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1183_3_lut_LC_4_23_5 (
            .in0(N__35619),
            .in1(N__24991),
            .in2(N__25021),
            .in3(_gnd_net_),
            .lcout(n1831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_4_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_4_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_4_23_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1179_3_lut_LC_4_23_6 (
            .in0(_gnd_net_),
            .in1(N__24874),
            .in2(N__24904),
            .in3(N__35615),
            .lcout(n1827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12375_3_lut_LC_4_23_7.C_ON=1'b0;
    defparam i12375_3_lut_LC_4_23_7.SEQ_MODE=4'b0000;
    defparam i12375_3_lut_LC_4_23_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 i12375_3_lut_LC_4_23_7 (
            .in0(_gnd_net_),
            .in1(N__24832),
            .in2(N__35628),
            .in3(N__24864),
            .lcout(n1826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_4_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_4_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_2_lut_LC_4_24_0 (
            .in0(_gnd_net_),
            .in1(N__28043),
            .in2(_gnd_net_),
            .in3(N__24697),
            .lcout(n1801),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(n12191),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_4_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_4_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_4_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_3_lut_LC_4_24_1 (
            .in0(_gnd_net_),
            .in1(N__25048),
            .in2(N__54589),
            .in3(N__25024),
            .lcout(n1800),
            .ltout(),
            .carryin(n12191),
            .carryout(n12192),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_4_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_4_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_4_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_4_lut_LC_4_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25017),
            .in3(N__24985),
            .lcout(n1799),
            .ltout(),
            .carryin(n12192),
            .carryout(n12193),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_4_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_4_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_4_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_5_lut_LC_4_24_3 (
            .in0(_gnd_net_),
            .in1(N__54083),
            .in2(N__24982),
            .in3(N__24949),
            .lcout(n1798),
            .ltout(),
            .carryin(n12193),
            .carryout(n12194),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_4_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_4_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_4_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_6_lut_LC_4_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24945),
            .in3(N__24910),
            .lcout(n1797),
            .ltout(),
            .carryin(n12194),
            .carryout(n12195),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_4_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_4_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_4_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_7_lut_LC_4_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27771),
            .in3(N__24907),
            .lcout(n1796),
            .ltout(),
            .carryin(n12195),
            .carryout(n12196),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_4_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_4_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_4_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_8_lut_LC_4_24_6 (
            .in0(_gnd_net_),
            .in1(N__54082),
            .in2(N__24903),
            .in3(N__24868),
            .lcout(n1795),
            .ltout(),
            .carryin(n12196),
            .carryout(n12197),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_4_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_4_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_4_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_9_lut_LC_4_24_7 (
            .in0(_gnd_net_),
            .in1(N__54084),
            .in2(N__24865),
            .in3(N__24826),
            .lcout(n1794),
            .ltout(),
            .carryin(n12197),
            .carryout(n12198),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_4_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_4_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_4_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_10_lut_LC_4_25_0 (
            .in0(_gnd_net_),
            .in1(N__55162),
            .in2(N__27885),
            .in3(N__24823),
            .lcout(n1793),
            .ltout(),
            .carryin(bfn_4_25_0_),
            .carryout(n12199),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_4_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_4_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_4_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_11_lut_LC_4_25_1 (
            .in0(_gnd_net_),
            .in1(N__55166),
            .in2(N__25246),
            .in3(N__25219),
            .lcout(n1792),
            .ltout(),
            .carryin(n12199),
            .carryout(n12200),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_4_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_4_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_4_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_12_lut_LC_4_25_2 (
            .in0(_gnd_net_),
            .in1(N__55163),
            .in2(N__27348),
            .in3(N__25216),
            .lcout(n1791),
            .ltout(),
            .carryin(n12200),
            .carryout(n12201),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_4_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_4_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_4_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_13_lut_LC_4_25_3 (
            .in0(_gnd_net_),
            .in1(N__55167),
            .in2(N__25213),
            .in3(N__25177),
            .lcout(n1790),
            .ltout(),
            .carryin(n12201),
            .carryout(n12202),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_4_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_4_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_4_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_14_lut_LC_4_25_4 (
            .in0(_gnd_net_),
            .in1(N__55164),
            .in2(N__25174),
            .in3(N__25144),
            .lcout(n1789),
            .ltout(),
            .carryin(n12202),
            .carryout(n12203),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_4_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_4_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_4_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_15_lut_LC_4_25_5 (
            .in0(_gnd_net_),
            .in1(N__55168),
            .in2(N__25141),
            .in3(N__25114),
            .lcout(n1788),
            .ltout(),
            .carryin(n12203),
            .carryout(n12204),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_4_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_4_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_4_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_16_lut_LC_4_25_6 (
            .in0(_gnd_net_),
            .in1(N__25111),
            .in2(N__55226),
            .in3(N__25087),
            .lcout(n1787),
            .ltout(),
            .carryin(n12204),
            .carryout(n12205),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_4_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_4_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_4_25_7.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1168_17_lut_LC_4_25_7 (
            .in0(N__55165),
            .in1(N__25084),
            .in2(N__35646),
            .in3(N__25063),
            .lcout(n1818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_4_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_4_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_4_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_2_lut_LC_4_26_0 (
            .in0(_gnd_net_),
            .in1(N__27563),
            .in2(_gnd_net_),
            .in3(N__25051),
            .lcout(n1601),
            .ltout(),
            .carryin(bfn_4_26_0_),
            .carryout(n12164),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_4_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_4_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_4_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_3_lut_LC_4_26_1 (
            .in0(_gnd_net_),
            .in1(N__54057),
            .in2(N__25492),
            .in3(N__25465),
            .lcout(n1600),
            .ltout(),
            .carryin(n12164),
            .carryout(n12165),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_4_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_4_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_4_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_4_lut_LC_4_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25461),
            .in3(N__25420),
            .lcout(n1599),
            .ltout(),
            .carryin(n12165),
            .carryout(n12166),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_4_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_4_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_4_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_5_lut_LC_4_26_3 (
            .in0(_gnd_net_),
            .in1(N__54058),
            .in2(N__25417),
            .in3(N__25393),
            .lcout(n1598),
            .ltout(),
            .carryin(n12166),
            .carryout(n12167),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_4_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_4_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_4_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_6_lut_LC_4_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25390),
            .in3(N__25360),
            .lcout(n1597),
            .ltout(),
            .carryin(n12167),
            .carryout(n12168),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_4_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_4_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_4_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_7_lut_LC_4_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25357),
            .in3(N__25327),
            .lcout(n1596),
            .ltout(),
            .carryin(n12168),
            .carryout(n12169),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_4_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_4_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_4_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_8_lut_LC_4_26_6 (
            .in0(_gnd_net_),
            .in1(N__54580),
            .in2(N__25324),
            .in3(N__25300),
            .lcout(n1595),
            .ltout(),
            .carryin(n12169),
            .carryout(n12170),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_4_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_4_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_4_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_9_lut_LC_4_26_7 (
            .in0(_gnd_net_),
            .in1(N__54059),
            .in2(N__25297),
            .in3(N__25258),
            .lcout(n1594),
            .ltout(),
            .carryin(n12170),
            .carryout(n12171),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_4_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_4_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_4_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_10_lut_LC_4_27_0 (
            .in0(_gnd_net_),
            .in1(N__54771),
            .in2(N__25590),
            .in3(N__25249),
            .lcout(n1593),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(n12172),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_4_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_4_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_4_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_11_lut_LC_4_27_1 (
            .in0(_gnd_net_),
            .in1(N__54584),
            .in2(N__25551),
            .in3(N__25744),
            .lcout(n1592),
            .ltout(),
            .carryin(n12172),
            .carryout(n12173),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_4_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_4_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_4_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_12_lut_LC_4_27_2 (
            .in0(_gnd_net_),
            .in1(N__54772),
            .in2(N__25809),
            .in3(N__25735),
            .lcout(n1591),
            .ltout(),
            .carryin(n12173),
            .carryout(n12174),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_4_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_4_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_4_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_13_lut_LC_4_27_3 (
            .in0(_gnd_net_),
            .in1(N__54585),
            .in2(N__25732),
            .in3(N__25693),
            .lcout(n1590),
            .ltout(),
            .carryin(n12174),
            .carryout(n12175),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_4_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_4_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_4_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_14_lut_LC_4_27_4 (
            .in0(_gnd_net_),
            .in1(N__25690),
            .in2(N__54975),
            .in3(N__25672),
            .lcout(n1589),
            .ltout(),
            .carryin(n12175),
            .carryout(n12176),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_4_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_4_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_4_27_5.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1034_15_lut_LC_4_27_5 (
            .in0(N__54773),
            .in1(N__35409),
            .in2(N__25669),
            .in3(N__25645),
            .lcout(n1620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i974_3_lut_LC_4_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_4_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_4_27_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i974_3_lut_LC_4_27_7 (
            .in0(_gnd_net_),
            .in1(N__25621),
            .in2(N__25603),
            .in3(N__35257),
            .lcout(n1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i973_3_lut_LC_4_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_4_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_4_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i973_3_lut_LC_4_28_0 (
            .in0(_gnd_net_),
            .in1(N__25968),
            .in2(N__25567),
            .in3(N__35256),
            .lcout(n1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i908_3_lut_LC_4_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_4_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_4_28_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i908_3_lut_LC_4_28_1 (
            .in0(_gnd_net_),
            .in1(N__25528),
            .in2(N__26026),
            .in3(N__36711),
            .lcout(n1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i905_3_lut_LC_4_28_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_4_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_4_28_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i905_3_lut_LC_4_28_2 (
            .in0(_gnd_net_),
            .in1(N__25990),
            .in2(N__36733),
            .in3(N__28390),
            .lcout(n1425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i906_3_lut_LC_4_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_4_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_4_28_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i906_3_lut_LC_4_28_3 (
            .in0(_gnd_net_),
            .in1(N__36715),
            .in2(N__28366),
            .in3(N__25981),
            .lcout(n1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i911_3_lut_LC_4_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_4_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_4_28_4.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i911_3_lut_LC_4_28_4 (
            .in0(N__26308),
            .in1(N__25948),
            .in2(N__36732),
            .in3(_gnd_net_),
            .lcout(n1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i903_3_lut_LC_4_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_4_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_4_28_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i903_3_lut_LC_4_28_5 (
            .in0(_gnd_net_),
            .in1(N__26221),
            .in2(N__25912),
            .in3(N__36719),
            .lcout(n1423),
            .ltout(n1423_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12807_4_lut_LC_4_28_6.C_ON=1'b0;
    defparam i12807_4_lut_LC_4_28_6.SEQ_MODE=4'b0000;
    defparam i12807_4_lut_LC_4_28_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12807_4_lut_LC_4_28_6 (
            .in0(N__25881),
            .in1(N__25864),
            .in2(N__25855),
            .in3(N__25852),
            .lcout(n1455),
            .ltout(n1455_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i972_3_lut_LC_4_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_4_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_4_28_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i972_3_lut_LC_4_28_7 (
            .in0(_gnd_net_),
            .in1(N__25844),
            .in2(N__25822),
            .in3(N__25819),
            .lcout(n1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i845_3_lut_LC_4_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_4_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_4_29_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i845_3_lut_LC_4_29_0 (
            .in0(N__25786),
            .in1(N__28296),
            .in2(_gnd_net_),
            .in3(N__36627),
            .lcout(n1333),
            .ltout(n1333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9926_3_lut_LC_4_29_1.C_ON=1'b0;
    defparam i9926_3_lut_LC_4_29_1.SEQ_MODE=4'b0000;
    defparam i9926_3_lut_LC_4_29_1.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9926_3_lut_LC_4_29_1 (
            .in0(_gnd_net_),
            .in1(N__26108),
            .in2(N__25762),
            .in3(N__26300),
            .lcout(),
            .ltout(n11640_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_72_LC_4_29_2.C_ON=1'b0;
    defparam i1_4_lut_adj_72_LC_4_29_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_72_LC_4_29_2.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_72_LC_4_29_2 (
            .in0(N__26090),
            .in1(N__26018),
            .in2(N__26197),
            .in3(N__26183),
            .lcout(),
            .ltout(n13315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12790_4_lut_LC_4_29_3.C_ON=1'b0;
    defparam i12790_4_lut_LC_4_29_3.SEQ_MODE=4'b0000;
    defparam i12790_4_lut_LC_4_29_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12790_4_lut_LC_4_29_3 (
            .in0(N__26220),
            .in1(N__26160),
            .in2(N__26146),
            .in3(N__28306),
            .lcout(n1356),
            .ltout(n1356_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i904_3_lut_LC_4_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_4_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_4_29_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i904_3_lut_LC_4_29_4 (
            .in0(_gnd_net_),
            .in1(N__28404),
            .in2(N__26143),
            .in3(N__26140),
            .lcout(n1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_4_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_4_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_4_29_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i21_3_lut_LC_4_29_5 (
            .in0(N__39535),
            .in1(N__33244),
            .in2(_gnd_net_),
            .in3(N__29905),
            .lcout(n299),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12787_1_lut_LC_4_29_6.C_ON=1'b0;
    defparam i12787_1_lut_LC_4_29_6.SEQ_MODE=4'b0000;
    defparam i12787_1_lut_LC_4_29_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12787_1_lut_LC_4_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36739),
            .in3(_gnd_net_),
            .lcout(n15259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i909_3_lut_LC_4_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_4_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_4_29_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i909_3_lut_LC_4_29_7 (
            .in0(_gnd_net_),
            .in1(N__26091),
            .in2(N__26074),
            .in3(N__36725),
            .lcout(n1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i841_3_lut_LC_4_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_4_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_4_30_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i841_3_lut_LC_4_30_0 (
            .in0(_gnd_net_),
            .in1(N__26032),
            .in2(N__28557),
            .in3(N__36626),
            .lcout(n1329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i839_3_lut_LC_4_30_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_4_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_4_30_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i839_3_lut_LC_4_30_1 (
            .in0(_gnd_net_),
            .in1(N__28227),
            .in2(N__36635),
            .in3(N__26002),
            .lcout(n1327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i838_3_lut_LC_4_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_4_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_4_30_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i838_3_lut_LC_4_30_2 (
            .in0(_gnd_net_),
            .in1(N__25996),
            .in2(N__28593),
            .in3(N__36618),
            .lcout(n1326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12774_4_lut_LC_4_30_3.C_ON=1'b0;
    defparam i12774_4_lut_LC_4_30_3.SEQ_MODE=4'b0000;
    defparam i12774_4_lut_LC_4_30_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12774_4_lut_LC_4_30_3 (
            .in0(N__28483),
            .in1(N__26352),
            .in2(N__26260),
            .in3(N__28693),
            .lcout(n1257),
            .ltout(n1257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12771_1_lut_LC_4_30_4.C_ON=1'b0;
    defparam i12771_1_lut_LC_4_30_4.SEQ_MODE=4'b0000;
    defparam i12771_1_lut_LC_4_30_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12771_1_lut_LC_4_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26332),
            .in3(_gnd_net_),
            .lcout(n15243),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i777_3_lut_LC_4_30_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_4_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_4_30_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i777_3_lut_LC_4_30_5 (
            .in0(N__28169),
            .in1(N__26329),
            .in2(_gnd_net_),
            .in3(N__36537),
            .lcout(n1233),
            .ltout(n1233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i844_3_lut_LC_4_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_4_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_4_30_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i844_3_lut_LC_4_30_6 (
            .in0(_gnd_net_),
            .in1(N__26317),
            .in2(N__26311),
            .in3(N__36625),
            .lcout(n1332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i840_3_lut_LC_4_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_4_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_4_30_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i840_3_lut_LC_4_30_7 (
            .in0(N__26284),
            .in1(_gnd_net_),
            .in2(N__36636),
            .in3(N__28536),
            .lcout(n1328),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i770_3_lut_LC_4_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_4_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_4_31_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i770_3_lut_LC_4_31_0 (
            .in0(_gnd_net_),
            .in1(N__28758),
            .in2(N__36546),
            .in3(N__26278),
            .lcout(n1226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i776_3_lut_LC_4_31_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_4_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_4_31_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i776_3_lut_LC_4_31_1 (
            .in0(_gnd_net_),
            .in1(N__26269),
            .in2(N__28629),
            .in3(N__36529),
            .lcout(n1232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i836_3_lut_LC_4_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_4_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_4_31_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i836_3_lut_LC_4_31_2 (
            .in0(_gnd_net_),
            .in1(N__26252),
            .in2(N__26230),
            .in3(N__36630),
            .lcout(n1324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12755_4_lut_LC_4_31_3.C_ON=1'b0;
    defparam i12755_4_lut_LC_4_31_3.SEQ_MODE=4'b0000;
    defparam i12755_4_lut_LC_4_31_3.LUT_INIT=16'b0000000000010101;
    LogicCell40 i12755_4_lut_LC_4_31_3 (
            .in0(N__28800),
            .in1(N__26359),
            .in2(N__26368),
            .in3(N__28738),
            .lcout(n1158),
            .ltout(n1158_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12752_1_lut_LC_4_31_4.C_ON=1'b0;
    defparam i12752_1_lut_LC_4_31_4.SEQ_MODE=4'b0000;
    defparam i12752_1_lut_LC_4_31_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12752_1_lut_LC_4_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26416),
            .in3(_gnd_net_),
            .lcout(n15224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i775_3_lut_LC_4_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_4_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_4_31_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i775_3_lut_LC_4_31_6 (
            .in0(_gnd_net_),
            .in1(N__28683),
            .in2(N__36545),
            .in3(N__26413),
            .lcout(n1231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i773_3_lut_LC_4_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_4_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_4_31_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i773_3_lut_LC_4_31_7 (
            .in0(_gnd_net_),
            .in1(N__26404),
            .in2(N__26391),
            .in3(N__36536),
            .lcout(n1229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i706_3_lut_LC_4_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_4_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_4_32_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i706_3_lut_LC_4_32_0 (
            .in0(_gnd_net_),
            .in1(N__30343),
            .in2(N__33904),
            .in3(N__36957),
            .lcout(n1130),
            .ltout(n1130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_68_LC_4_32_1.C_ON=1'b0;
    defparam i1_2_lut_adj_68_LC_4_32_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_68_LC_4_32_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_68_LC_4_32_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26371),
            .in3(N__28649),
            .lcout(n14068),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9991_4_lut_LC_4_32_3.C_ON=1'b0;
    defparam i9991_4_lut_LC_4_32_3.SEQ_MODE=4'b0000;
    defparam i9991_4_lut_LC_4_32_3.LUT_INIT=16'b1111110011111000;
    LogicCell40 i9991_4_lut_LC_4_32_3 (
            .in0(N__28177),
            .in1(N__28682),
            .in2(N__30453),
            .in3(N__28622),
            .lcout(n11706),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i1_LC_4_32_4 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i1_LC_4_32_4 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i1_LC_4_32_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i1_LC_4_32_4  (
            .in0(N__38171),
            .in1(N__28120),
            .in2(_gnd_net_),
            .in3(N__27945),
            .lcout(h2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_118_LC_5_17_0.C_ON=1'b0;
    defparam i1_4_lut_adj_118_LC_5_17_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_118_LC_5_17_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_118_LC_5_17_0 (
            .in0(N__37391),
            .in1(N__30728),
            .in2(N__34511),
            .in3(N__30800),
            .lcout(n13798),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_5_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_5_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_5_17_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1709_3_lut_LC_5_17_1 (
            .in0(_gnd_net_),
            .in1(N__30972),
            .in2(N__38943),
            .in3(N__28849),
            .lcout(n2613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_5_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1653_3_lut_LC_5_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1653_3_lut_LC_5_17_2 (
            .in0(_gnd_net_),
            .in1(N__29134),
            .in2(N__31240),
            .in3(N__35048),
            .lcout(n2525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_5_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_5_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_5_17_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1655_3_lut_LC_5_17_3 (
            .in0(N__28921),
            .in1(_gnd_net_),
            .in2(N__35092),
            .in3(N__28941),
            .lcout(n2527),
            .ltout(n2527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_119_LC_5_17_4.C_ON=1'b0;
    defparam i1_4_lut_adj_119_LC_5_17_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_119_LC_5_17_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_119_LC_5_17_4 (
            .in0(N__34346),
            .in1(N__30665),
            .in2(N__26443),
            .in3(N__30852),
            .lcout(),
            .ltout(n13796_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_120_LC_5_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_120_LC_5_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_120_LC_5_17_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_120_LC_5_17_5 (
            .in0(N__26440),
            .in1(N__34598),
            .in2(N__26434),
            .in3(N__31107),
            .lcout(n13804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_5_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_5_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_5_17_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1654_3_lut_LC_5_17_6 (
            .in0(N__28876),
            .in1(_gnd_net_),
            .in2(N__28912),
            .in3(N__35047),
            .lcout(n2526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_116_LC_5_18_0.C_ON=1'b0;
    defparam i1_3_lut_adj_116_LC_5_18_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_116_LC_5_18_0.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_116_LC_5_18_0 (
            .in0(_gnd_net_),
            .in1(N__29105),
            .in2(N__29073),
            .in3(N__29322),
            .lcout(),
            .ltout(n14354_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_117_LC_5_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_117_LC_5_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_117_LC_5_18_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_117_LC_5_18_1 (
            .in0(N__31571),
            .in1(N__29279),
            .in2(N__26431),
            .in3(N__26428),
            .lcout(),
            .ltout(n14224_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12906_4_lut_LC_5_18_2.C_ON=1'b0;
    defparam i12906_4_lut_LC_5_18_2.SEQ_MODE=4'b0000;
    defparam i12906_4_lut_LC_5_18_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12906_4_lut_LC_5_18_2 (
            .in0(N__31193),
            .in1(N__29782),
            .in2(N__26422),
            .in3(N__29248),
            .lcout(n2445),
            .ltout(n2445_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_5_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_5_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_5_18_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1649_3_lut_LC_5_18_3 (
            .in0(N__29106),
            .in1(_gnd_net_),
            .in2(N__26419),
            .in3(N__29092),
            .lcout(n2521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_5_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_5_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_5_18_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1650_3_lut_LC_5_18_4 (
            .in0(_gnd_net_),
            .in1(N__29119),
            .in2(N__31297),
            .in3(N__35085),
            .lcout(n2522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_5_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_5_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_5_18_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1645_3_lut_LC_5_18_5 (
            .in0(N__29323),
            .in1(_gnd_net_),
            .in2(N__35108),
            .in3(N__29299),
            .lcout(n2517),
            .ltout(n2517_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_122_LC_5_18_6.C_ON=1'b0;
    defparam i1_4_lut_adj_122_LC_5_18_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_122_LC_5_18_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_122_LC_5_18_6 (
            .in0(N__29734),
            .in1(N__31049),
            .in2(N__26509),
            .in3(N__26506),
            .lcout(n13810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_5_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_5_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_5_18_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1646_3_lut_LC_5_18_7 (
            .in0(_gnd_net_),
            .in1(N__29069),
            .in2(N__35107),
            .in3(N__29053),
            .lcout(n2518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_19_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1642_3_lut_LC_5_19_0 (
            .in0(_gnd_net_),
            .in1(N__29263),
            .in2(N__29284),
            .in3(N__35053),
            .lcout(n2514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1 (
            .in0(N__29691),
            .in1(_gnd_net_),
            .in2(N__26500),
            .in3(N__36205),
            .lcout(n2217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_19_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1582_3_lut_LC_5_19_2 (
            .in0(N__26488),
            .in1(_gnd_net_),
            .in2(N__34926),
            .in3(N__32241),
            .lcout(n2422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_19_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1593_3_lut_LC_5_19_3 (
            .in0(N__37505),
            .in1(N__26476),
            .in2(_gnd_net_),
            .in3(N__34890),
            .lcout(n2433),
            .ltout(n2433_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9955_3_lut_LC_5_19_4.C_ON=1'b0;
    defparam i9955_3_lut_LC_5_19_4.SEQ_MODE=4'b0000;
    defparam i9955_3_lut_LC_5_19_4.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9955_3_lut_LC_5_19_4 (
            .in0(_gnd_net_),
            .in1(N__37679),
            .in2(N__26464),
            .in3(N__29657),
            .lcout(n11670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_5_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_5_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_5_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1575_3_lut_LC_5_19_5 (
            .in0(_gnd_net_),
            .in1(N__39013),
            .in2(N__26455),
            .in3(N__34894),
            .lcout(n2415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_5_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_5_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_5_19_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1506_3_lut_LC_5_19_6 (
            .in0(_gnd_net_),
            .in1(N__31969),
            .in2(N__32008),
            .in3(N__39104),
            .lcout(n2314),
            .ltout(n2314_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_5_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_5_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_5_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1573_3_lut_LC_5_19_7 (
            .in0(_gnd_net_),
            .in1(N__26581),
            .in2(N__26572),
            .in3(N__34895),
            .lcout(n2413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_5_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_5_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_5_20_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1518_3_lut_LC_5_20_0 (
            .in0(N__31839),
            .in1(_gnd_net_),
            .in2(N__31816),
            .in3(N__39095),
            .lcout(n2326),
            .ltout(n2326_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1585_3_lut_LC_5_20_1 (
            .in0(N__34865),
            .in1(_gnd_net_),
            .in2(N__26569),
            .in3(N__26566),
            .lcout(n2425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_5_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_5_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_5_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1524_3_lut_LC_5_20_2 (
            .in0(_gnd_net_),
            .in1(N__31521),
            .in2(N__31498),
            .in3(N__39096),
            .lcout(n2332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_20_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1657_3_lut_LC_5_20_3 (
            .in0(_gnd_net_),
            .in1(N__28996),
            .in2(N__35103),
            .in3(N__29025),
            .lcout(n2529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_20_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1592_3_lut_LC_5_20_4 (
            .in0(_gnd_net_),
            .in1(N__26554),
            .in2(N__26529),
            .in3(N__34864),
            .lcout(n2432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12853_4_lut_LC_5_20_5.C_ON=1'b0;
    defparam i12853_4_lut_LC_5_20_5.SEQ_MODE=4'b0000;
    defparam i12853_4_lut_LC_5_20_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12853_4_lut_LC_5_20_5 (
            .in0(N__32039),
            .in1(N__31991),
            .in2(N__31953),
            .in3(N__26542),
            .lcout(n2247),
            .ltout(n2247_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_5_20_6.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1525_3_lut_LC_5_20_6 (
            .in0(N__32161),
            .in1(N__31534),
            .in2(N__26536),
            .in3(_gnd_net_),
            .lcout(n2333),
            .ltout(n2333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10051_4_lut_LC_5_20_7.C_ON=1'b0;
    defparam i10051_4_lut_LC_5_20_7.SEQ_MODE=4'b0000;
    defparam i10051_4_lut_LC_5_20_7.LUT_INIT=16'b1111111110101000;
    LogicCell40 i10051_4_lut_LC_5_20_7 (
            .in0(N__26861),
            .in1(N__37512),
            .in2(N__26845),
            .in3(N__26842),
            .lcout(n11766),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_5_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_5_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_5_21_0.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i1446_3_lut_LC_5_21_0 (
            .in0(N__36201),
            .in1(N__27105),
            .in2(N__26812),
            .in3(_gnd_net_),
            .lcout(n2222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9902_3_lut_LC_5_21_1.C_ON=1'b0;
    defparam i9902_3_lut_LC_5_21_1.SEQ_MODE=4'b0000;
    defparam i9902_3_lut_LC_5_21_1.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9902_3_lut_LC_5_21_1 (
            .in0(_gnd_net_),
            .in1(N__27977),
            .in2(N__26797),
            .in3(N__26622),
            .lcout(),
            .ltout(n11616_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_99_LC_5_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_99_LC_5_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_99_LC_5_21_2.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_99_LC_5_21_2 (
            .in0(N__26769),
            .in1(N__26739),
            .in2(N__26713),
            .in3(N__26693),
            .lcout(n13382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12518_1_lut_LC_5_21_3.C_ON=1'b0;
    defparam i12518_1_lut_LC_5_21_3.SEQ_MODE=4'b0000;
    defparam i12518_1_lut_LC_5_21_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12518_1_lut_LC_5_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35751),
            .lcout(n14990),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_5_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_5_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_5_21_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1321_3_lut_LC_5_21_5 (
            .in0(N__37599),
            .in1(N__26680),
            .in2(_gnd_net_),
            .in3(N__35871),
            .lcout(n2033),
            .ltout(n2033_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_5_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_5_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_5_21_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1388_3_lut_LC_5_21_6 (
            .in0(_gnd_net_),
            .in1(N__26650),
            .in2(N__26638),
            .in3(N__36018),
            .lcout(n2132),
            .ltout(n2132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_5_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_5_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_5_21_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1455_3_lut_LC_5_21_7 (
            .in0(_gnd_net_),
            .in1(N__26611),
            .in2(N__26599),
            .in3(N__36200),
            .lcout(n2231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_5_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_5_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_5_22_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1320_3_lut_LC_5_22_0 (
            .in0(_gnd_net_),
            .in1(N__27193),
            .in2(N__27489),
            .in3(N__35872),
            .lcout(n2032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_5_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_5_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_5_22_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1379_3_lut_LC_5_22_1 (
            .in0(_gnd_net_),
            .in1(N__27151),
            .in2(N__36045),
            .in3(N__27132),
            .lcout(n2123),
            .ltout(n2123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_96_LC_5_22_2.C_ON=1'b0;
    defparam i1_4_lut_adj_96_LC_5_22_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_96_LC_5_22_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_96_LC_5_22_2 (
            .in0(N__29370),
            .in1(N__29181),
            .in2(N__27091),
            .in3(N__29571),
            .lcout(),
            .ltout(n13746_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_98_LC_5_22_3.C_ON=1'b0;
    defparam i1_4_lut_adj_98_LC_5_22_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_98_LC_5_22_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_98_LC_5_22_3 (
            .in0(N__27088),
            .in1(N__27596),
            .in2(N__27067),
            .in3(N__27064),
            .lcout(),
            .ltout(n13754_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_100_LC_5_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_100_LC_5_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_100_LC_5_22_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_100_LC_5_22_4 (
            .in0(N__27058),
            .in1(N__29676),
            .in2(N__27031),
            .in3(N__27028),
            .lcout(n13760),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_5_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_5_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_5_23_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1241_3_lut_LC_5_23_0 (
            .in0(N__27006),
            .in1(_gnd_net_),
            .in2(N__35754),
            .in3(N__26986),
            .lcout(n1921),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_5_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_5_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_5_23_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1252_3_lut_LC_5_23_1 (
            .in0(_gnd_net_),
            .in1(N__28020),
            .in2(N__26947),
            .in3(N__35729),
            .lcout(n1932),
            .ltout(n1932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9971_4_lut_LC_5_23_2.C_ON=1'b0;
    defparam i9971_4_lut_LC_5_23_2.SEQ_MODE=4'b0000;
    defparam i9971_4_lut_LC_5_23_2.LUT_INIT=16'b1111111111100000;
    LogicCell40 i9971_4_lut_LC_5_23_2 (
            .in0(N__27482),
            .in1(N__37598),
            .in2(N__26911),
            .in3(N__26900),
            .lcout(n11686),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_5_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_5_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_5_23_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1249_3_lut_LC_5_23_3 (
            .in0(_gnd_net_),
            .in1(N__27547),
            .in2(N__27277),
            .in3(N__35733),
            .lcout(n1929),
            .ltout(n1929_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_90_LC_5_23_4.C_ON=1'b0;
    defparam i1_2_lut_adj_90_LC_5_23_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_90_LC_5_23_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_90_LC_5_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27511),
            .in3(N__27438),
            .lcout(n14136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_5_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_5_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_5_23_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1253_3_lut_LC_5_23_5 (
            .in0(N__27502),
            .in1(N__32695),
            .in2(_gnd_net_),
            .in3(N__35728),
            .lcout(n1933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_5_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_5_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_5_23_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1250_3_lut_LC_5_23_6 (
            .in0(_gnd_net_),
            .in1(N__27680),
            .in2(N__35753),
            .in3(N__27463),
            .lcout(n1930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_5_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_5_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_5_23_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1237_3_lut_LC_5_23_7 (
            .in0(_gnd_net_),
            .in1(N__27427),
            .in2(N__27415),
            .in3(N__35737),
            .lcout(n1917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_5_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_5_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_5_24_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1175_3_lut_LC_5_24_0 (
            .in0(_gnd_net_),
            .in1(N__27361),
            .in2(N__27355),
            .in3(N__35611),
            .lcout(n1823),
            .ltout(n1823_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_84_LC_5_24_1.C_ON=1'b0;
    defparam i1_3_lut_adj_84_LC_5_24_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_84_LC_5_24_1.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_84_LC_5_24_1 (
            .in0(N__27302),
            .in1(_gnd_net_),
            .in2(N__27280),
            .in3(N__27778),
            .lcout(),
            .ltout(n14126_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_85_LC_5_24_2.C_ON=1'b0;
    defparam i1_4_lut_adj_85_LC_5_24_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_85_LC_5_24_2.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_85_LC_5_24_2 (
            .in0(N__27276),
            .in1(N__27240),
            .in2(N__27214),
            .in3(N__27658),
            .lcout(n14128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_5_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_5_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_5_24_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1177_3_lut_LC_5_24_3 (
            .in0(N__27199),
            .in1(_gnd_net_),
            .in2(N__35624),
            .in3(N__27886),
            .lcout(n1825),
            .ltout(n1825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_83_LC_5_24_4.C_ON=1'b0;
    defparam i1_4_lut_adj_83_LC_5_24_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_83_LC_5_24_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_83_LC_5_24_4 (
            .in0(N__27821),
            .in1(N__27797),
            .in2(N__27781),
            .in3(N__27725),
            .lcout(n14122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_5_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_5_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_5_24_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1180_3_lut_LC_5_24_6 (
            .in0(_gnd_net_),
            .in1(N__27772),
            .in2(N__27751),
            .in3(N__35607),
            .lcout(n1828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9973_4_lut_LC_5_24_7.C_ON=1'b0;
    defparam i9973_4_lut_LC_5_24_7.SEQ_MODE=4'b0000;
    defparam i9973_4_lut_LC_5_24_7.LUT_INIT=16'b1111110011111000;
    LogicCell40 i9973_4_lut_LC_5_24_7 (
            .in0(N__32690),
            .in1(N__27710),
            .in2(N__27681),
            .in3(N__28019),
            .lcout(n11688),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_5_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_5_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_5_25_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1376_3_lut_LC_5_25_0 (
            .in0(_gnd_net_),
            .in1(N__27651),
            .in2(N__27622),
            .in3(N__36036),
            .lcout(n2120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_5_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_5_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_5_25_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i19_3_lut_LC_5_25_1 (
            .in0(N__33301),
            .in1(N__39465),
            .in2(_gnd_net_),
            .in3(N__29951),
            .lcout(n301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_5_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_5_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_5_25_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_5_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29819),
            .lcout(n21_adj_645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_5_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_5_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_5_25_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_5_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39309),
            .in3(_gnd_net_),
            .lcout(n29_adj_653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_5_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_5_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_5_25_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_5_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30064),
            .lcout(n4_adj_628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_5_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_5_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_5_25_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i17_3_lut_LC_5_25_7 (
            .in0(N__32971),
            .in1(N__39466),
            .in2(_gnd_net_),
            .in3(N__30140),
            .lcout(n303),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_5_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_5_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_5_26_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1185_3_lut_LC_5_26_0 (
            .in0(N__28060),
            .in1(N__28044),
            .in2(_gnd_net_),
            .in3(N__35623),
            .lcout(n1833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_5_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_5_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_5_26_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_5_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36287),
            .lcout(n8_adj_632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_5_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_5_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_5_26_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i13_3_lut_LC_5_26_2 (
            .in0(N__33034),
            .in1(N__39396),
            .in2(_gnd_net_),
            .in3(N__29826),
            .lcout(n307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i0_LC_5_26_3 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i0_LC_5_26_3 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i0_LC_5_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i0_LC_5_26_3  (
            .in0(N__38132),
            .in1(N__28446),
            .in2(_gnd_net_),
            .in3(N__27952),
            .lcout(h3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_5_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_5_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_5_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_5_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39394),
            .lcout(n2_adj_626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_5_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_5_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_5_26_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i14_3_lut_LC_5_26_5 (
            .in0(N__39395),
            .in1(N__33022),
            .in2(_gnd_net_),
            .in3(N__38305),
            .lcout(n306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_5_26_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_5_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_5_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_5_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30106),
            .lcout(n6_adj_630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_5_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_5_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_5_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_5_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32182),
            .lcout(n22_adj_646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_5_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_5_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_5_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_5_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29976),
            .lcout(n16_adj_640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10846_3_lut_LC_5_27_2.C_ON=1'b0;
    defparam i10846_3_lut_LC_5_27_2.SEQ_MODE=4'b0000;
    defparam i10846_3_lut_LC_5_27_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 i10846_3_lut_LC_5_27_2 (
            .in0(_gnd_net_),
            .in1(N__33427),
            .in2(N__30318),
            .in3(N__28210),
            .lcout(),
            .ltout(n13257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10847_3_lut_LC_5_27_3.C_ON=1'b0;
    defparam i10847_3_lut_LC_5_27_3.SEQ_MODE=4'b0000;
    defparam i10847_3_lut_LC_5_27_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 i10847_3_lut_LC_5_27_3 (
            .in0(N__39444),
            .in1(_gnd_net_),
            .in2(N__28102),
            .in3(N__30068),
            .lcout(n830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2139_2_lut_LC_5_27_4.C_ON=1'b0;
    defparam i2139_2_lut_LC_5_27_4.SEQ_MODE=4'b0000;
    defparam i2139_2_lut_LC_5_27_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2139_2_lut_LC_5_27_4 (
            .in0(_gnd_net_),
            .in1(N__39443),
            .in2(_gnd_net_),
            .in3(N__33367),
            .lcout(n402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_5_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_5_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_5_27_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_5_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30390),
            .in3(_gnd_net_),
            .lcout(n9_adj_633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_5_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_5_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_5_27_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i18_3_lut_LC_5_27_6 (
            .in0(N__29977),
            .in1(N__33325),
            .in2(_gnd_net_),
            .in3(N__39445),
            .lcout(n302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_5_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_5_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_5_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_5_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29955),
            .lcout(n15_adj_639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_2_lut_LC_5_28_0.C_ON=1'b1;
    defparam add_709_2_lut_LC_5_28_0.SEQ_MODE=4'b0000;
    defparam add_709_2_lut_LC_5_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_2_lut_LC_5_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30199),
            .in3(N__28069),
            .lcout(n2290),
            .ltout(),
            .carryin(bfn_5_28_0_),
            .carryout(n12096),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_3_lut_LC_5_28_1.C_ON=1'b1;
    defparam add_709_3_lut_LC_5_28_1.SEQ_MODE=4'b0000;
    defparam add_709_3_lut_LC_5_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_3_lut_LC_5_28_1 (
            .in0(_gnd_net_),
            .in1(N__54599),
            .in2(N__30085),
            .in3(N__28066),
            .lcout(n2289),
            .ltout(),
            .carryin(n12096),
            .carryout(n12097),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_4_lut_LC_5_28_2.C_ON=1'b1;
    defparam add_709_4_lut_LC_5_28_2.SEQ_MODE=4'b0000;
    defparam add_709_4_lut_LC_5_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_4_lut_LC_5_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30157),
            .in3(N__28063),
            .lcout(n2288),
            .ltout(),
            .carryin(n12097),
            .carryout(n12098),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_5_lut_LC_5_28_3.C_ON=1'b1;
    defparam add_709_5_lut_LC_5_28_3.SEQ_MODE=4'b0000;
    defparam add_709_5_lut_LC_5_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_5_lut_LC_5_28_3 (
            .in0(_gnd_net_),
            .in1(N__30043),
            .in2(N__54977),
            .in3(N__28204),
            .lcout(n2287),
            .ltout(),
            .carryin(n12098),
            .carryout(n12099),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_6_lut_LC_5_28_4.C_ON=1'b1;
    defparam add_709_6_lut_LC_5_28_4.SEQ_MODE=4'b0000;
    defparam add_709_6_lut_LC_5_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_6_lut_LC_5_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30223),
            .in3(N__28201),
            .lcout(n2286),
            .ltout(),
            .carryin(n12099),
            .carryout(n12100),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_709_7_lut_LC_5_28_5.C_ON=1'b0;
    defparam add_709_7_lut_LC_5_28_5.SEQ_MODE=4'b0000;
    defparam add_709_7_lut_LC_5_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_709_7_lut_LC_5_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28198),
            .in3(N__28189),
            .lcout(n2285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10850_3_lut_LC_5_28_6.C_ON=1'b0;
    defparam i10850_3_lut_LC_5_28_6.SEQ_MODE=4'b0000;
    defparam i10850_3_lut_LC_5_28_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 i10850_3_lut_LC_5_28_6 (
            .in0(_gnd_net_),
            .in1(N__33496),
            .in2(N__30317),
            .in3(N__28186),
            .lcout(),
            .ltout(n13261_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10851_3_lut_LC_5_28_7.C_ON=1'b0;
    defparam i10851_3_lut_LC_5_28_7.SEQ_MODE=4'b0000;
    defparam i10851_3_lut_LC_5_28_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 i10851_3_lut_LC_5_28_7 (
            .in0(N__39486),
            .in1(_gnd_net_),
            .in2(N__28180),
            .in3(N__30121),
            .lcout(n832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_5_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_5_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_5_29_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i3_3_lut_LC_5_29_0 (
            .in0(N__32929),
            .in1(N__39497),
            .in2(_gnd_net_),
            .in3(N__32479),
            .lcout(n317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_5_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_5_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_5_29_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i23_3_lut_LC_5_29_1 (
            .in0(N__39496),
            .in1(N__33184),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(n297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i1_LC_5_29_2 .C_ON=1'b0;
    defparam \debounce.reg_B_i1_LC_5_29_2 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i1_LC_5_29_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i1_LC_5_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28147),
            .lcout(reg_B_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56054),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_5_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_5_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_5_29_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_5_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32209),
            .lcout(n30_adj_654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i0_LC_5_29_4 .C_ON=1'b0;
    defparam \debounce.reg_B_i0_LC_5_29_4 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i0_LC_5_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i0_LC_5_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28477),
            .lcout(reg_B_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56054),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_5_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_5_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_5_29_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_5_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30036),
            .lcout(n11_adj_635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10848_3_lut_LC_5_29_6.C_ON=1'b0;
    defparam i10848_3_lut_LC_5_29_6.SEQ_MODE=4'b0000;
    defparam i10848_3_lut_LC_5_29_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10848_3_lut_LC_5_29_6 (
            .in0(_gnd_net_),
            .in1(N__30307),
            .in2(N__33472),
            .in3(N__28426),
            .lcout(n13259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_5_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_5_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_5_30_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29871),
            .lcout(n12_adj_636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i837_3_lut_LC_5_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_5_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_5_30_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i837_3_lut_LC_5_30_2 (
            .in0(_gnd_net_),
            .in1(N__36631),
            .in2(N__28713),
            .in3(N__28420),
            .lcout(n1325),
            .ltout(n1325_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_71_LC_5_30_3.C_ON=1'b0;
    defparam i1_4_lut_adj_71_LC_5_30_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_71_LC_5_30_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_71_LC_5_30_3 (
            .in0(N__28382),
            .in1(N__28355),
            .in2(N__28339),
            .in3(N__28322),
            .lcout(n13734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_5_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_5_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_5_30_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i22_3_lut_LC_5_30_4 (
            .in0(N__33214),
            .in1(N__39534),
            .in2(_gnd_net_),
            .in3(N__29872),
            .lcout(n298),
            .ltout(n298_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9928_3_lut_LC_5_30_5.C_ON=1'b0;
    defparam i9928_3_lut_LC_5_30_5.SEQ_MODE=4'b0000;
    defparam i9928_3_lut_LC_5_30_5.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9928_3_lut_LC_5_30_5 (
            .in0(_gnd_net_),
            .in1(N__28278),
            .in2(N__28267),
            .in3(N__28259),
            .lcout(n11642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i772_3_lut_LC_5_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_5_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_5_30_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i772_3_lut_LC_5_30_6 (
            .in0(_gnd_net_),
            .in1(N__36540),
            .in2(N__28659),
            .in3(N__28243),
            .lcout(n1228),
            .ltout(n1228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_69_LC_5_30_7.C_ON=1'b0;
    defparam i1_3_lut_adj_69_LC_5_30_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_69_LC_5_30_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_69_LC_5_30_7 (
            .in0(_gnd_net_),
            .in1(N__28583),
            .in2(N__28717),
            .in3(N__28706),
            .lcout(n14078),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i708_3_lut_LC_5_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_5_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_5_31_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i708_3_lut_LC_5_31_0 (
            .in0(N__33928),
            .in1(N__30355),
            .in2(N__36958),
            .in3(_gnd_net_),
            .lcout(n1132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i705_3_lut_LC_5_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_5_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_5_31_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i705_3_lut_LC_5_31_2 (
            .in0(_gnd_net_),
            .in1(N__30328),
            .in2(N__36959),
            .in3(N__33850),
            .lcout(n1129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i709_3_lut_LC_5_31_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_5_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_5_31_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i709_3_lut_LC_5_31_3 (
            .in0(_gnd_net_),
            .in1(N__33948),
            .in2(N__30367),
            .in3(N__36941),
            .lcout(n1133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i771_3_lut_LC_5_31_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_5_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_5_31_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i771_3_lut_LC_5_31_4 (
            .in0(N__36539),
            .in1(_gnd_net_),
            .in2(N__30543),
            .in3(N__28603),
            .lcout(n1227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i774_3_lut_LC_5_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_5_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_5_31_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i774_3_lut_LC_5_31_5 (
            .in0(_gnd_net_),
            .in1(N__36538),
            .in2(N__30449),
            .in3(N__28567),
            .lcout(n1230),
            .ltout(n1230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_70_LC_5_31_6.C_ON=1'b0;
    defparam i1_4_lut_adj_70_LC_5_31_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_70_LC_5_31_6.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_70_LC_5_31_6 (
            .in0(N__28532),
            .in1(N__28511),
            .in2(N__28492),
            .in3(N__28489),
            .lcout(n13318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_5_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_5_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_5_31_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_5_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30418),
            .in3(_gnd_net_),
            .lcout(n10_adj_634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i703_3_lut_LC_5_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_5_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_5_32_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i703_3_lut_LC_5_32_2 (
            .in0(_gnd_net_),
            .in1(N__30586),
            .in2(N__30517),
            .in3(N__36948),
            .lcout(n1127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i701_3_lut_LC_5_32_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_5_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_5_32_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i701_3_lut_LC_5_32_4 (
            .in0(_gnd_net_),
            .in1(N__30565),
            .in2(N__33778),
            .in3(N__36950),
            .lcout(n1125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i702_3_lut_LC_5_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_5_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_5_32_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i702_3_lut_LC_5_32_6 (
            .in0(_gnd_net_),
            .in1(N__30577),
            .in2(N__30493),
            .in3(N__36949),
            .lcout(n1126),
            .ltout(n1126_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_63_LC_5_32_7.C_ON=1'b0;
    defparam i1_3_lut_adj_63_LC_5_32_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_63_LC_5_32_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_63_LC_5_32_7 (
            .in0(_gnd_net_),
            .in1(N__30536),
            .in2(N__28768),
            .in3(N__28754),
            .lcout(n13994),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_14_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_14_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_2_lut_LC_6_14_0 (
            .in0(_gnd_net_),
            .in1(N__32776),
            .in2(_gnd_net_),
            .in3(N__28732),
            .lcout(n2601),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(n12339),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_14_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_14_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_3_lut_LC_6_14_1 (
            .in0(_gnd_net_),
            .in1(N__38985),
            .in2(N__53063),
            .in3(N__28729),
            .lcout(n2600),
            .ltout(),
            .carryin(n12339),
            .carryout(n12340),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_14_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_14_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_4_lut_LC_6_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31627),
            .in3(N__28726),
            .lcout(n2599),
            .ltout(),
            .carryin(n12340),
            .carryout(n12341),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_14_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_14_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_5_lut_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(N__53064),
            .in2(N__34461),
            .in3(N__28723),
            .lcout(n2598),
            .ltout(),
            .carryin(n12341),
            .carryout(n12342),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_14_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_14_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_6_lut_LC_6_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34297),
            .in3(N__28720),
            .lcout(n2597),
            .ltout(),
            .carryin(n12342),
            .carryout(n12343),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_14_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_14_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_7_lut_LC_6_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30619),
            .in3(N__28834),
            .lcout(n2596),
            .ltout(),
            .carryin(n12343),
            .carryout(n12344),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_14_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_14_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_8_lut_LC_6_14_6 (
            .in0(_gnd_net_),
            .in1(N__52985),
            .in2(N__30745),
            .in3(N__28831),
            .lcout(n2595),
            .ltout(),
            .carryin(n12344),
            .carryout(n12345),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_14_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_14_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_9_lut_LC_6_14_7 (
            .in0(_gnd_net_),
            .in1(N__53065),
            .in2(N__34414),
            .in3(N__28828),
            .lcout(n2594),
            .ltout(),
            .carryin(n12345),
            .carryout(n12346),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_15_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_15_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_10_lut_LC_6_15_0 (
            .in0(_gnd_net_),
            .in1(N__53007),
            .in2(N__34518),
            .in3(N__28825),
            .lcout(n2593),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(n12347),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_15_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_15_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_11_lut_LC_6_15_1 (
            .in0(_gnd_net_),
            .in1(N__53014),
            .in2(N__30813),
            .in3(N__28822),
            .lcout(n2592),
            .ltout(),
            .carryin(n12347),
            .carryout(n12348),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_15_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_15_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_15_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_12_lut_LC_6_15_2 (
            .in0(_gnd_net_),
            .in1(N__53008),
            .in2(N__30853),
            .in3(N__28819),
            .lcout(n2591),
            .ltout(),
            .carryin(n12348),
            .carryout(n12349),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_15_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_15_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_15_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_13_lut_LC_6_15_3 (
            .in0(_gnd_net_),
            .in1(N__53015),
            .in2(N__30670),
            .in3(N__28816),
            .lcout(n2590),
            .ltout(),
            .carryin(n12349),
            .carryout(n12350),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_15_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_15_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_15_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_14_lut_LC_6_15_4 (
            .in0(_gnd_net_),
            .in1(N__53009),
            .in2(N__34353),
            .in3(N__28813),
            .lcout(n2589),
            .ltout(),
            .carryin(n12350),
            .carryout(n12351),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_15_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_15_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_15_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_15_lut_LC_6_15_5 (
            .in0(_gnd_net_),
            .in1(N__53016),
            .in2(N__37404),
            .in3(N__28810),
            .lcout(n2588),
            .ltout(),
            .carryin(n12351),
            .carryout(n12352),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_15_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_15_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_15_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_16_lut_LC_6_15_6 (
            .in0(_gnd_net_),
            .in1(N__53010),
            .in2(N__34609),
            .in3(N__28867),
            .lcout(n2587),
            .ltout(),
            .carryin(n12352),
            .carryout(n12353),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_15_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_15_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_15_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_17_lut_LC_6_15_7 (
            .in0(_gnd_net_),
            .in1(N__31108),
            .in2(N__53108),
            .in3(N__28864),
            .lcout(n2586),
            .ltout(),
            .carryin(n12353),
            .carryout(n12354),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_16_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_18_lut_LC_6_16_0 (
            .in0(_gnd_net_),
            .in1(N__31056),
            .in2(N__53662),
            .in3(N__28861),
            .lcout(n2585),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(n12355),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_16_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_19_lut_LC_6_16_1 (
            .in0(_gnd_net_),
            .in1(N__53340),
            .in2(N__30783),
            .in3(N__28858),
            .lcout(n2584),
            .ltout(),
            .carryin(n12355),
            .carryout(n12356),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_16_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_16_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_20_lut_LC_6_16_2 (
            .in0(_gnd_net_),
            .in1(N__30993),
            .in2(N__53663),
            .in3(N__28855),
            .lcout(n2583),
            .ltout(),
            .carryin(n12356),
            .carryout(n12357),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_16_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_16_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_21_lut_LC_6_16_3 (
            .in0(_gnd_net_),
            .in1(N__31555),
            .in2(N__53347),
            .in3(N__28852),
            .lcout(n2582),
            .ltout(),
            .carryin(n12357),
            .carryout(n12358),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_16_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_16_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_22_lut_LC_6_16_4 (
            .in0(_gnd_net_),
            .in1(N__30971),
            .in2(N__53664),
            .in3(N__28843),
            .lcout(n2581),
            .ltout(),
            .carryin(n12358),
            .carryout(n12359),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_16_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_23_lut_LC_6_16_5 (
            .in0(_gnd_net_),
            .in1(N__34547),
            .in2(N__53348),
            .in3(N__28840),
            .lcout(n2580),
            .ltout(),
            .carryin(n12359),
            .carryout(n12360),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_16_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_16_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_24_lut_LC_6_16_6 (
            .in0(_gnd_net_),
            .in1(N__53124),
            .in2(N__31177),
            .in3(N__28837),
            .lcout(n2579),
            .ltout(),
            .carryin(n12360),
            .carryout(n12361),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_16_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_16_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_16_7.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1704_25_lut_LC_6_16_7 (
            .in0(N__53125),
            .in1(N__30931),
            .in2(N__35157),
            .in3(N__29044),
            .lcout(n2610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_2_lut_LC_6_17_0 (
            .in0(_gnd_net_),
            .in1(N__37686),
            .in2(_gnd_net_),
            .in3(N__29041),
            .lcout(n2501),
            .ltout(),
            .carryin(bfn_6_17_0_),
            .carryout(n12317),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_3_lut_LC_6_17_1 (
            .in0(_gnd_net_),
            .in1(N__53177),
            .in2(N__29446),
            .in3(N__29038),
            .lcout(n2500),
            .ltout(),
            .carryin(n12317),
            .carryout(n12318),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_4_lut_LC_6_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29665),
            .in3(N__29035),
            .lcout(n2499),
            .ltout(),
            .carryin(n12318),
            .carryout(n12319),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_5_lut_LC_6_17_3 (
            .in0(_gnd_net_),
            .in1(N__53178),
            .in2(N__29424),
            .in3(N__29032),
            .lcout(n2498),
            .ltout(),
            .carryin(n12319),
            .carryout(n12320),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_6_lut_LC_6_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29029),
            .in3(N__28987),
            .lcout(n2497),
            .ltout(),
            .carryin(n12320),
            .carryout(n12321),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_7_lut_LC_6_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28984),
            .in3(N__28951),
            .lcout(n2496),
            .ltout(),
            .carryin(n12321),
            .carryout(n12322),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_8_lut_LC_6_17_6 (
            .in0(_gnd_net_),
            .in1(N__53736),
            .in2(N__28948),
            .in3(N__28915),
            .lcout(n2495),
            .ltout(),
            .carryin(n12322),
            .carryout(n12323),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_9_lut_LC_6_17_7 (
            .in0(_gnd_net_),
            .in1(N__53179),
            .in2(N__28911),
            .in3(N__28870),
            .lcout(n2494),
            .ltout(),
            .carryin(n12323),
            .carryout(n12324),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_10_lut_LC_6_18_0 (
            .in0(_gnd_net_),
            .in1(N__53349),
            .in2(N__31232),
            .in3(N__29128),
            .lcout(n2493),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(n12325),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_11_lut_LC_6_18_1 (
            .in0(_gnd_net_),
            .in1(N__53356),
            .in2(N__30891),
            .in3(N__29125),
            .lcout(n2492),
            .ltout(),
            .carryin(n12325),
            .carryout(n12326),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_12_lut_LC_6_18_2 (
            .in0(_gnd_net_),
            .in1(N__53350),
            .in2(N__30699),
            .in3(N__29122),
            .lcout(n2491),
            .ltout(),
            .carryin(n12326),
            .carryout(n12327),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_13_lut_LC_6_18_3 (
            .in0(_gnd_net_),
            .in1(N__53357),
            .in2(N__31296),
            .in3(N__29113),
            .lcout(n2490),
            .ltout(),
            .carryin(n12327),
            .carryout(n12328),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_14_lut_LC_6_18_4 (
            .in0(_gnd_net_),
            .in1(N__53351),
            .in2(N__29110),
            .in3(N__29086),
            .lcout(n2489),
            .ltout(),
            .carryin(n12328),
            .carryout(n12329),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_15_lut_LC_6_18_5 (
            .in0(_gnd_net_),
            .in1(N__53358),
            .in2(N__29224),
            .in3(N__29083),
            .lcout(n2488),
            .ltout(),
            .carryin(n12329),
            .carryout(n12330),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_16_lut_LC_6_18_6 (
            .in0(_gnd_net_),
            .in1(N__53352),
            .in2(N__31137),
            .in3(N__29080),
            .lcout(n2487),
            .ltout(),
            .carryin(n12330),
            .carryout(n12331),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_17_lut_LC_6_18_7 (
            .in0(_gnd_net_),
            .in1(N__29077),
            .in2(N__53665),
            .in3(N__29047),
            .lcout(n2486),
            .ltout(),
            .carryin(n12331),
            .carryout(n12332),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_18_lut_LC_6_19_0 (
            .in0(_gnd_net_),
            .in1(N__29321),
            .in2(N__53666),
            .in3(N__29293),
            .lcout(n2485),
            .ltout(),
            .carryin(bfn_6_19_0_),
            .carryout(n12333),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_19_lut_LC_6_19_1 (
            .in0(_gnd_net_),
            .in1(N__53366),
            .in2(N__31032),
            .in3(N__29290),
            .lcout(n2484),
            .ltout(),
            .carryin(n12333),
            .carryout(n12334),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_20_lut_LC_6_19_2 (
            .in0(_gnd_net_),
            .in1(N__31578),
            .in2(N__53667),
            .in3(N__29287),
            .lcout(n2483),
            .ltout(),
            .carryin(n12334),
            .carryout(n12335),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_21_lut_LC_6_19_3 (
            .in0(_gnd_net_),
            .in1(N__29280),
            .in2(N__54676),
            .in3(N__29257),
            .lcout(n2482),
            .ltout(),
            .carryin(n12335),
            .carryout(n12336),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_22_lut_LC_6_19_4 (
            .in0(_gnd_net_),
            .in1(N__29781),
            .in2(N__53668),
            .in3(N__29254),
            .lcout(n2481),
            .ltout(),
            .carryin(n12336),
            .carryout(n12337),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_23_lut_LC_6_19_5 (
            .in0(_gnd_net_),
            .in1(N__31194),
            .in2(N__54677),
            .in3(N__29251),
            .lcout(n2480),
            .ltout(),
            .carryin(n12337),
            .carryout(n12338),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_19_6.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1637_24_lut_LC_6_19_6 (
            .in0(N__53373),
            .in1(N__29247),
            .in2(N__35133),
            .in3(N__29227),
            .lcout(n2511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_6_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_6_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_6_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1648_3_lut_LC_6_19_7 (
            .in0(_gnd_net_),
            .in1(N__29223),
            .in2(N__29191),
            .in3(N__35052),
            .lcout(n2520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1449_rep_27_3_lut_LC_6_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1449_rep_27_3_lut_LC_6_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1449_rep_27_3_lut_LC_6_20_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1449_rep_27_3_lut_LC_6_20_0 (
            .in0(_gnd_net_),
            .in1(N__29182),
            .in2(N__36198),
            .in3(N__29149),
            .lcout(n2225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_6_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1448_3_lut_LC_6_20_1 (
            .in0(_gnd_net_),
            .in1(N__29521),
            .in2(N__29506),
            .in3(N__36173),
            .lcout(n2224),
            .ltout(n2224_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_101_LC_6_20_2.C_ON=1'b0;
    defparam i1_2_lut_adj_101_LC_6_20_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_101_LC_6_20_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_101_LC_6_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29473),
            .in3(N__31835),
            .lcout(),
            .ltout(n14174_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_102_LC_6_20_3.C_ON=1'b0;
    defparam i1_4_lut_adj_102_LC_6_20_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_102_LC_6_20_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_102_LC_6_20_3 (
            .in0(N__31892),
            .in1(N__31793),
            .in2(N__29470),
            .in3(N__32498),
            .lcout(),
            .ltout(n14178_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_103_LC_6_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_103_LC_6_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_103_LC_6_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_103_LC_6_20_4 (
            .in0(N__31730),
            .in1(N__31761),
            .in2(N__29467),
            .in3(N__31701),
            .lcout(n14184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_20_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1660_3_lut_LC_6_20_5 (
            .in0(N__29455),
            .in1(_gnd_net_),
            .in2(N__29445),
            .in3(N__35067),
            .lcout(n2532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_6_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_6_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_6_20_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1658_3_lut_LC_6_20_6 (
            .in0(N__29425),
            .in1(_gnd_net_),
            .in2(N__35102),
            .in3(N__29398),
            .lcout(n2530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_6_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_6_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_6_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1450_3_lut_LC_6_20_7 (
            .in0(_gnd_net_),
            .in1(N__29389),
            .in2(N__29374),
            .in3(N__36169),
            .lcout(n2226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_6_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_6_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_6_21_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1661_3_lut_LC_6_21_0 (
            .in0(N__29338),
            .in1(N__37690),
            .in2(_gnd_net_),
            .in3(N__35075),
            .lcout(n2533),
            .ltout(n2533_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9967_3_lut_LC_6_21_1.C_ON=1'b0;
    defparam i9967_3_lut_LC_6_21_1.SEQ_MODE=4'b0000;
    defparam i9967_3_lut_LC_6_21_1.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9967_3_lut_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__32771),
            .in2(N__29326),
            .in3(N__31619),
            .lcout(),
            .ltout(n11682_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_121_LC_6_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_121_LC_6_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_121_LC_6_21_2.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_121_LC_6_21_2 (
            .in0(N__30602),
            .in1(N__34280),
            .in2(N__29737),
            .in3(N__34443),
            .lcout(n13397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_6_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_6_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_6_21_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1517_3_lut_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__31777),
            .in2(N__31801),
            .in3(N__39098),
            .lcout(n2325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_6_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_6_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_6_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1374_3_lut_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(N__29725),
            .in2(N__29716),
            .in3(N__36044),
            .lcout(n2118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_6_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_6_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_6_21_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1659_3_lut_LC_6_21_6 (
            .in0(N__29661),
            .in1(_gnd_net_),
            .in2(N__29641),
            .in3(N__35074),
            .lcout(n2531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_6_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_6_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_6_21_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1513_3_lut_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__31734),
            .in2(N__31714),
            .in3(N__39097),
            .lcout(n2321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_6_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_6_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_6_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1380_3_lut_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__29625),
            .in2(N__29599),
            .in3(N__36037),
            .lcout(n2124),
            .ltout(n2124_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_6_22_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1447_3_lut_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(N__29560),
            .in2(N__29545),
            .in3(N__36199),
            .lcout(n2223),
            .ltout(n2223_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_6_22_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1514_3_lut_LC_6_22_2 (
            .in0(N__31744),
            .in1(_gnd_net_),
            .in2(N__29542),
            .in3(N__39119),
            .lcout(n2322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_22_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1507_3_lut_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(N__32046),
            .in2(N__39144),
            .in3(N__32017),
            .lcout(n2315),
            .ltout(n2315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_6_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_6_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_6_22_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1574_3_lut_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(N__29797),
            .in2(N__29785),
            .in3(N__34931),
            .lcout(n2414),
            .ltout(n2414_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_6_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_6_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_6_22_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1641_3_lut_LC_6_22_5 (
            .in0(N__35105),
            .in1(_gnd_net_),
            .in2(N__29764),
            .in3(N__29761),
            .lcout(n2513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12903_1_lut_LC_6_22_6.C_ON=1'b0;
    defparam i12903_1_lut_LC_6_22_6.SEQ_MODE=4'b0000;
    defparam i12903_1_lut_LC_6_22_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12903_1_lut_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35104),
            .lcout(n15375),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12850_1_lut_LC_6_22_7.C_ON=1'b0;
    defparam i12850_1_lut_LC_6_22_7.SEQ_MODE=4'b0000;
    defparam i12850_1_lut_LC_6_22_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12850_1_lut_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39143),
            .in3(_gnd_net_),
            .lcout(n15322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i0_LC_6_23_0 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i0_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i0_LC_6_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i0_LC_6_23_0  (
            .in0(_gnd_net_),
            .in1(N__32568),
            .in2(_gnd_net_),
            .in3(N__29752),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(\quad_counter0.n12623 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i1_LC_6_23_1 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i1_LC_6_23_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i1_LC_6_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i1_LC_6_23_1  (
            .in0(_gnd_net_),
            .in1(N__49765),
            .in2(N__32590),
            .in3(N__29749),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(\quad_counter0.n12623 ),
            .carryout(\quad_counter0.n12624 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i2_LC_6_23_2 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i2_LC_6_23_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i2_LC_6_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i2_LC_6_23_2  (
            .in0(_gnd_net_),
            .in1(N__32475),
            .in2(N__49829),
            .in3(N__29746),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(\quad_counter0.n12624 ),
            .carryout(\quad_counter0.n12625 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i3_LC_6_23_3 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i3_LC_6_23_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i3_LC_6_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i3_LC_6_23_3  (
            .in0(_gnd_net_),
            .in1(N__49769),
            .in2(N__32208),
            .in3(N__29743),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(\quad_counter0.n12625 ),
            .carryout(\quad_counter0.n12626 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i4_LC_6_23_4 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i4_LC_6_23_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i4_LC_6_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i4_LC_6_23_4  (
            .in0(_gnd_net_),
            .in1(N__39302),
            .in2(N__49830),
            .in3(N__29740),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(\quad_counter0.n12626 ),
            .carryout(\quad_counter0.n12627 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i5_LC_6_23_5 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i5_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i5_LC_6_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i5_LC_6_23_5  (
            .in0(_gnd_net_),
            .in1(N__49773),
            .in2(N__32737),
            .in3(N__29848),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(\quad_counter0.n12627 ),
            .carryout(\quad_counter0.n12628 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i6_LC_6_23_6 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i6_LC_6_23_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i6_LC_6_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i6_LC_6_23_6  (
            .in0(_gnd_net_),
            .in1(N__37772),
            .in2(N__49831),
            .in3(N__29845),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(\quad_counter0.n12628 ),
            .carryout(\quad_counter0.n12629 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i7_LC_6_23_7 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i7_LC_6_23_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i7_LC_6_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i7_LC_6_23_7  (
            .in0(_gnd_net_),
            .in1(N__49777),
            .in2(N__37986),
            .in3(N__29842),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(\quad_counter0.n12629 ),
            .carryout(\quad_counter0.n12630 ),
            .clk(N__56040),
            .ce(N__50436),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i8_LC_6_24_0 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i8_LC_6_24_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i8_LC_6_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i8_LC_6_24_0  (
            .in0(_gnd_net_),
            .in1(N__49832),
            .in2(N__32800),
            .in3(N__29839),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(\quad_counter0.n12631 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i9_LC_6_24_1 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i9_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i9_LC_6_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i9_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__37712),
            .in2(N__49880),
            .in3(N__29836),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(\quad_counter0.n12631 ),
            .carryout(\quad_counter0.n12632 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i10_LC_6_24_2 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i10_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i10_LC_6_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i10_LC_6_24_2  (
            .in0(_gnd_net_),
            .in1(N__49836),
            .in2(N__37547),
            .in3(N__29833),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(\quad_counter0.n12632 ),
            .carryout(\quad_counter0.n12633 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i11_LC_6_24_3 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i11_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i11_LC_6_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i11_LC_6_24_3  (
            .in0(_gnd_net_),
            .in1(N__32181),
            .in2(N__49881),
            .in3(N__29830),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(\quad_counter0.n12633 ),
            .carryout(\quad_counter0.n12634 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i12_LC_6_24_4 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i12_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i12_LC_6_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i12_LC_6_24_4  (
            .in0(_gnd_net_),
            .in1(N__49840),
            .in2(N__29827),
            .in3(N__29803),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(\quad_counter0.n12634 ),
            .carryout(\quad_counter0.n12635 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i13_LC_6_24_5 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i13_LC_6_24_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i13_LC_6_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i13_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(N__38297),
            .in2(N__49882),
            .in3(N__29800),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(\quad_counter0.n12635 ),
            .carryout(\quad_counter0.n12636 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i14_LC_6_24_6 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i14_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i14_LC_6_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i14_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(N__49844),
            .in2(N__37632),
            .in3(N__29986),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(\quad_counter0.n12636 ),
            .carryout(\quad_counter0.n12637 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i15_LC_6_24_7 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i15_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i15_LC_6_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i15_LC_6_24_7  (
            .in0(_gnd_net_),
            .in1(N__32715),
            .in2(N__49883),
            .in3(N__29983),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(\quad_counter0.n12637 ),
            .carryout(\quad_counter0.n12638 ),
            .clk(N__56043),
            .ce(N__50437),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i16_LC_6_25_0 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i16_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i16_LC_6_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i16_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__49848),
            .in2(N__30145),
            .in3(N__29980),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(bfn_6_25_0_),
            .carryout(\quad_counter0.n12639 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i17_LC_6_25_1 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i17_LC_6_25_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i17_LC_6_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i17_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__29975),
            .in2(N__49884),
            .in3(N__29959),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(\quad_counter0.n12639 ),
            .carryout(\quad_counter0.n12640 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i18_LC_6_25_2 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i18_LC_6_25_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i18_LC_6_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i18_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__49852),
            .in2(N__29956),
            .in3(N__29932),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(\quad_counter0.n12640 ),
            .carryout(\quad_counter0.n12641 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i19_LC_6_25_3 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i19_LC_6_25_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i19_LC_6_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i19_LC_6_25_3  (
            .in0(_gnd_net_),
            .in1(N__29922),
            .in2(N__49885),
            .in3(N__29908),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(\quad_counter0.n12641 ),
            .carryout(\quad_counter0.n12642 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i20_LC_6_25_4 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i20_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i20_LC_6_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i20_LC_6_25_4  (
            .in0(_gnd_net_),
            .in1(N__49856),
            .in2(N__29901),
            .in3(N__29875),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(\quad_counter0.n12642 ),
            .carryout(\quad_counter0.n12643 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i21_LC_6_25_5 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i21_LC_6_25_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i21_LC_6_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i21_LC_6_25_5  (
            .in0(_gnd_net_),
            .in1(N__29865),
            .in2(N__49886),
            .in3(N__29851),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(\quad_counter0.n12643 ),
            .carryout(\quad_counter0.n12644 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i22_LC_6_25_6 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i22_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i22_LC_6_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i22_LC_6_25_6  (
            .in0(_gnd_net_),
            .in1(N__49860),
            .in2(N__30035),
            .in3(N__30013),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(\quad_counter0.n12644 ),
            .carryout(\quad_counter0.n12645 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i23_LC_6_25_7 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i23_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i23_LC_6_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i23_LC_6_25_7  (
            .in0(_gnd_net_),
            .in1(N__30407),
            .in2(N__49887),
            .in3(N__30010),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(\quad_counter0.n12645 ),
            .carryout(\quad_counter0.n12646 ),
            .clk(N__56047),
            .ce(N__50432),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i24_LC_6_26_0 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i24_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i24_LC_6_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i24_LC_6_26_0  (
            .in0(_gnd_net_),
            .in1(N__30389),
            .in2(N__49888),
            .in3(N__30007),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(bfn_6_26_0_),
            .carryout(\quad_counter0.n12647 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i25_LC_6_26_1 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i25_LC_6_26_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i25_LC_6_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i25_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__49867),
            .in2(N__36297),
            .in3(N__30004),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(\quad_counter0.n12647 ),
            .carryout(\quad_counter0.n12648 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i26_LC_6_26_2 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i26_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i26_LC_6_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i26_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(N__30271),
            .in2(N__49889),
            .in3(N__30001),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(\quad_counter0.n12648 ),
            .carryout(\quad_counter0.n12649 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i27_LC_6_26_3 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i27_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i27_LC_6_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i27_LC_6_26_3  (
            .in0(_gnd_net_),
            .in1(N__49871),
            .in2(N__30120),
            .in3(N__29998),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(\quad_counter0.n12649 ),
            .carryout(\quad_counter0.n12650 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i28_LC_6_26_4 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i28_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i28_LC_6_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i28_LC_6_26_4  (
            .in0(_gnd_net_),
            .in1(N__38257),
            .in2(N__49890),
            .in3(N__29995),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(\quad_counter0.n12650 ),
            .carryout(\quad_counter0.n12651 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i29_LC_6_26_5 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i29_LC_6_26_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i29_LC_6_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i29_LC_6_26_5  (
            .in0(_gnd_net_),
            .in1(N__49875),
            .in2(N__30075),
            .in3(N__29992),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(\quad_counter0.n12651 ),
            .carryout(\quad_counter0.n12652 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i30_LC_6_26_6 .C_ON=1'b1;
    defparam \quad_counter0.position_637__i30_LC_6_26_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i30_LC_6_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_637__i30_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(N__30245),
            .in2(N__49891),
            .in3(N__29989),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(\quad_counter0.n12652 ),
            .carryout(\quad_counter0.n12653 ),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_637__i31_LC_6_26_7 .C_ON=1'b0;
    defparam \quad_counter0.position_637__i31_LC_6_26_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_637__i31_LC_6_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.position_637__i31_LC_6_26_7  (
            .in0(N__39467),
            .in1(N__49879),
            .in2(_gnd_net_),
            .in3(N__30148),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56049),
            .ce(N__50431),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_27_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30144),
            .lcout(n17_adj_641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37628),
            .lcout(n19_adj_643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_6_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_6_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_6_27_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_6_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30239),
            .lcout(n3_adj_627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_6_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_6_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_6_27_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_6_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32716),
            .lcout(n18_adj_642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_6_27_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_6_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_6_27_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_6_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32799),
            .lcout(n25_adj_649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_6_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_6_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_6_27_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_6_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37713),
            .lcout(n24_adj_648),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_6_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_6_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_6_27_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i28_3_lut_LC_6_27_7 (
            .in0(_gnd_net_),
            .in1(N__39442),
            .in2(N__30116),
            .in3(N__33491),
            .lcout(n175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_6_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_6_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_6_28_0.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i1_3_lut_LC_6_28_0 (
            .in0(N__39476),
            .in1(_gnd_net_),
            .in2(N__32539),
            .in3(N__32572),
            .lcout(n319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_6_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_6_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_6_28_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i30_3_lut_LC_6_28_1 (
            .in0(_gnd_net_),
            .in1(N__39471),
            .in2(N__30076),
            .in3(N__33419),
            .lcout(n404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_124_LC_6_28_2.C_ON=1'b0;
    defparam i1_3_lut_adj_124_LC_6_28_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_124_LC_6_28_2.LUT_INIT=16'b1100000000000000;
    LogicCell40 i1_3_lut_adj_124_LC_6_28_2 (
            .in0(_gnd_net_),
            .in1(N__30187),
            .in2(N__39529),
            .in3(N__33393),
            .lcout(),
            .ltout(n14170_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i500_4_lut_LC_6_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_6_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_6_28_3.LUT_INIT=16'b1010100000001000;
    LogicCell40 encoder0_position_31__I_0_i500_4_lut_LC_6_28_3 (
            .in0(N__33363),
            .in1(N__39475),
            .in2(N__30208),
            .in3(N__30205),
            .lcout(n828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_6_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_6_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_6_28_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i27_3_lut_LC_6_28_4 (
            .in0(_gnd_net_),
            .in1(N__30276),
            .in2(N__39528),
            .in3(N__33522),
            .lcout(n293),
            .ltout(n293_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_65_LC_6_28_5.C_ON=1'b0;
    defparam i1_4_lut_adj_65_LC_6_28_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_65_LC_6_28_5.LUT_INIT=16'b1111111011001100;
    LogicCell40 i1_4_lut_adj_65_LC_6_28_5 (
            .in0(N__33492),
            .in1(N__33420),
            .in2(N__30190),
            .in3(N__33462),
            .lcout(n5_adj_697),
            .ltout(n5_adj_697_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_66_LC_6_28_6.C_ON=1'b0;
    defparam i1_3_lut_adj_66_LC_6_28_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_66_LC_6_28_6.LUT_INIT=16'b1100000000000000;
    LogicCell40 i1_3_lut_adj_66_LC_6_28_6 (
            .in0(_gnd_net_),
            .in1(N__33392),
            .in2(N__30181),
            .in3(N__33362),
            .lcout(n13254),
            .ltout(n13254_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10852_3_lut_LC_6_28_7.C_ON=1'b0;
    defparam i10852_3_lut_LC_6_28_7.SEQ_MODE=4'b0000;
    defparam i10852_3_lut_LC_6_28_7.LUT_INIT=16'b1100101011001010;
    LogicCell40 i10852_3_lut_LC_6_28_7 (
            .in0(N__33523),
            .in1(N__30178),
            .in2(N__30172),
            .in3(_gnd_net_),
            .lcout(n13263),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10849_3_lut_LC_6_29_0.C_ON=1'b0;
    defparam i10849_3_lut_LC_6_29_0.SEQ_MODE=4'b0000;
    defparam i10849_3_lut_LC_6_29_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 i10849_3_lut_LC_6_29_0 (
            .in0(_gnd_net_),
            .in1(N__38262),
            .in2(N__39531),
            .in3(N__30169),
            .lcout(n831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12294_3_lut_LC_6_29_1.C_ON=1'b0;
    defparam i12294_3_lut_LC_6_29_1.SEQ_MODE=4'b0000;
    defparam i12294_3_lut_LC_6_29_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 i12294_3_lut_LC_6_29_1 (
            .in0(_gnd_net_),
            .in1(N__39481),
            .in2(N__30277),
            .in3(N__30163),
            .lcout(n833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_6_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_6_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_6_29_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i29_3_lut_LC_6_29_2 (
            .in0(_gnd_net_),
            .in1(N__38261),
            .in2(N__39530),
            .in3(N__33461),
            .lcout(n174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_6_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_6_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i635_rep_55_3_lut_LC_6_29_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i635_rep_55_3_lut_LC_6_29_3 (
            .in0(_gnd_net_),
            .in1(N__34129),
            .in2(N__33793),
            .in3(N__34018),
            .lcout(n1027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10844_3_lut_LC_6_29_4.C_ON=1'b0;
    defparam i10844_3_lut_LC_6_29_4.SEQ_MODE=4'b0000;
    defparam i10844_3_lut_LC_6_29_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10844_3_lut_LC_6_29_4 (
            .in0(_gnd_net_),
            .in1(N__30319),
            .in2(N__33394),
            .in3(N__30286),
            .lcout(),
            .ltout(n13255_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10845_3_lut_LC_6_29_5.C_ON=1'b0;
    defparam i10845_3_lut_LC_6_29_5.SEQ_MODE=4'b0000;
    defparam i10845_3_lut_LC_6_29_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 i10845_3_lut_LC_6_29_5 (
            .in0(N__30249),
            .in1(_gnd_net_),
            .in2(N__30280),
            .in3(N__39485),
            .lcout(n829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_6_29_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_6_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_6_29_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_6_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30272),
            .lcout(n7_adj_631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_6_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_6_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_6_29_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i31_3_lut_LC_6_29_7 (
            .in0(_gnd_net_),
            .in1(N__39480),
            .in2(N__30250),
            .in3(N__33388),
            .lcout(n403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9995_4_lut_LC_6_30_0.C_ON=1'b0;
    defparam i9995_4_lut_LC_6_30_0.SEQ_MODE=4'b0000;
    defparam i9995_4_lut_LC_6_30_0.LUT_INIT=16'b1111111111100000;
    LogicCell40 i9995_4_lut_LC_6_30_0 (
            .in0(N__34082),
            .in1(N__34064),
            .in2(N__33737),
            .in3(N__34034),
            .lcout(n11710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9997_4_lut_LC_6_30_1.C_ON=1'b0;
    defparam i9997_4_lut_LC_6_30_1.SEQ_MODE=4'b0000;
    defparam i9997_4_lut_LC_6_30_1.LUT_INIT=16'b1111111011110000;
    LogicCell40 i9997_4_lut_LC_6_30_1 (
            .in0(N__36261),
            .in1(N__33572),
            .in2(N__34250),
            .in3(N__33707),
            .lcout(),
            .ltout(n11712_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10107_4_lut_LC_6_30_2.C_ON=1'b0;
    defparam i10107_4_lut_LC_6_30_2.SEQ_MODE=4'b0000;
    defparam i10107_4_lut_LC_6_30_2.LUT_INIT=16'b1111111110000000;
    LogicCell40 i10107_4_lut_LC_6_30_2 (
            .in0(N__33656),
            .in1(N__33620),
            .in2(N__30214),
            .in3(N__33598),
            .lcout(n861),
            .ltout(n861_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i573_3_lut_LC_6_30_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_6_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_6_30_3.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i573_3_lut_LC_6_30_3 (
            .in0(N__36262),
            .in1(N__33346),
            .in2(N__30211),
            .in3(_gnd_net_),
            .lcout(n933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_6_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_6_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_6_30_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i25_3_lut_LC_6_30_4 (
            .in0(_gnd_net_),
            .in1(N__39532),
            .in2(N__33118),
            .in3(N__30391),
            .lcout(n295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i569_3_lut_LC_6_30_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_6_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_6_30_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i569_3_lut_LC_6_30_5 (
            .in0(_gnd_net_),
            .in1(N__33657),
            .in2(N__33637),
            .in3(N__34215),
            .lcout(n929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i568_3_lut_LC_6_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_6_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_6_30_6.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i568_3_lut_LC_6_30_6 (
            .in0(N__33607),
            .in1(N__33621),
            .in2(N__34224),
            .in3(_gnd_net_),
            .lcout(n928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i571_3_lut_LC_6_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_6_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_6_30_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i571_3_lut_LC_6_30_7 (
            .in0(_gnd_net_),
            .in1(N__33708),
            .in2(N__33679),
            .in3(N__34214),
            .lcout(n931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_6_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_6_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_6_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_2_lut_LC_6_31_0 (
            .in0(_gnd_net_),
            .in1(N__33947),
            .in2(_gnd_net_),
            .in3(N__30358),
            .lcout(n1101),
            .ltout(),
            .carryin(bfn_6_31_0_),
            .carryout(n12114),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_6_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_6_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_6_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_3_lut_LC_6_31_1 (
            .in0(_gnd_net_),
            .in1(N__55227),
            .in2(N__33927),
            .in3(N__30349),
            .lcout(n1100),
            .ltout(),
            .carryin(n12114),
            .carryout(n12115),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_6_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_6_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_6_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_4_lut_LC_6_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33970),
            .in3(N__30346),
            .lcout(n1099),
            .ltout(),
            .carryin(n12115),
            .carryout(n12116),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_6_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_6_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_6_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_5_lut_LC_6_31_3 (
            .in0(_gnd_net_),
            .in1(N__55228),
            .in2(N__33897),
            .in3(N__30331),
            .lcout(n1098),
            .ltout(),
            .carryin(n12116),
            .carryout(n12117),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_6_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_6_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_6_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_6_lut_LC_6_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33849),
            .in3(N__30322),
            .lcout(n1097),
            .ltout(),
            .carryin(n12117),
            .carryout(n12118),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_6_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_6_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_6_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_7_lut_LC_6_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33874),
            .in3(N__30589),
            .lcout(n1096),
            .ltout(),
            .carryin(n12118),
            .carryout(n12119),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_6_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_6_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_6_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_8_lut_LC_6_31_6 (
            .in0(_gnd_net_),
            .in1(N__55229),
            .in2(N__30516),
            .in3(N__30580),
            .lcout(n1095),
            .ltout(),
            .carryin(n12119),
            .carryout(n12120),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_6_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_6_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_6_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_9_lut_LC_6_31_7 (
            .in0(_gnd_net_),
            .in1(N__30488),
            .in2(N__55246),
            .in3(N__30571),
            .lcout(n1094),
            .ltout(),
            .carryin(n12120),
            .carryout(n12121),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_6_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_6_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_6_32_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_31__I_0_add_699_10_lut_LC_6_32_0 (
            .in0(N__54598),
            .in1(N__33771),
            .in2(_gnd_net_),
            .in3(N__30568),
            .lcout(n1093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i636_3_lut_LC_6_32_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_6_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_6_32_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i636_3_lut_LC_6_32_1 (
            .in0(_gnd_net_),
            .in1(N__34171),
            .in2(N__33808),
            .in3(N__34015),
            .lcout(n1028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i704_3_lut_LC_6_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_6_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_6_32_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i704_3_lut_LC_6_32_2 (
            .in0(_gnd_net_),
            .in1(N__33873),
            .in2(N__30559),
            .in3(N__36951),
            .lcout(n1128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12741_4_lut_LC_6_32_4.C_ON=1'b0;
    defparam i12741_4_lut_LC_6_32_4.SEQ_MODE=4'b0000;
    defparam i12741_4_lut_LC_6_32_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12741_4_lut_LC_6_32_4 (
            .in0(N__30509),
            .in1(N__33770),
            .in2(N__30492),
            .in3(N__33826),
            .lcout(n1059),
            .ltout(n1059_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i707_3_lut_LC_6_32_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_6_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_6_32_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i707_3_lut_LC_6_32_5 (
            .in0(N__33969),
            .in1(_gnd_net_),
            .in2(N__30466),
            .in3(N__30463),
            .lcout(n1131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_6_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_6_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_6_32_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i24_3_lut_LC_6_32_6 (
            .in0(_gnd_net_),
            .in1(N__39533),
            .in2(N__33151),
            .in3(N__30417),
            .lcout(n296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_14_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_14_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_7_16_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_7_16_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_7_16_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1718_3_lut_LC_7_16_4 (
            .in0(_gnd_net_),
            .in1(N__30829),
            .in2(N__30669),
            .in3(N__38900),
            .lcout(n2622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12929_1_lut_LC_7_16_5.C_ON=1'b0;
    defparam i12929_1_lut_LC_7_16_5.SEQ_MODE=4'b0000;
    defparam i12929_1_lut_LC_7_16_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12929_1_lut_LC_7_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38930),
            .in3(_gnd_net_),
            .lcout(n15401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1720_rep_19_3_lut_LC_7_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1720_rep_19_3_lut_LC_7_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1720_rep_19_3_lut_LC_7_17_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1720_rep_19_3_lut_LC_7_17_0 (
            .in0(_gnd_net_),
            .in1(N__30823),
            .in2(N__30814),
            .in3(N__38849),
            .lcout(n2624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_7_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_7_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_7_17_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1712_3_lut_LC_7_17_1 (
            .in0(N__30784),
            .in1(_gnd_net_),
            .in2(N__38898),
            .in3(N__30760),
            .lcout(n2616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1723_rep_21_3_lut_LC_7_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1723_rep_21_3_lut_LC_7_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1723_rep_21_3_lut_LC_7_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1723_rep_21_3_lut_LC_7_17_2 (
            .in0(_gnd_net_),
            .in1(N__30754),
            .in2(N__30744),
            .in3(N__38850),
            .lcout(n2627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_7_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_7_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_7_17_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1651_3_lut_LC_7_17_3 (
            .in0(_gnd_net_),
            .in1(N__30712),
            .in2(N__30706),
            .in3(N__35101),
            .lcout(n2523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_7_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_7_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_7_17_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1711_3_lut_LC_7_17_4 (
            .in0(_gnd_net_),
            .in1(N__30640),
            .in2(N__31000),
            .in3(N__38860),
            .lcout(n2615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_7_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_7_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_7_17_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1724_3_lut_LC_7_17_5 (
            .in0(_gnd_net_),
            .in1(N__30628),
            .in2(N__38897),
            .in3(N__30618),
            .lcout(n2628),
            .ltout(n2628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_57_LC_7_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_57_LC_7_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_57_LC_7_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_57_LC_7_17_6 (
            .in0(N__38624),
            .in1(N__37425),
            .in2(N__31069),
            .in3(N__39254),
            .lcout(n14278),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_7_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_7_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_7_17_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1713_3_lut_LC_7_17_7 (
            .in0(_gnd_net_),
            .in1(N__31066),
            .in2(N__38899),
            .in3(N__31060),
            .lcout(n2617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_7_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_7_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_7_18_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_i1644_3_lut_LC_7_18_0 (
            .in0(N__31033),
            .in1(N__35084),
            .in2(_gnd_net_),
            .in3(N__31006),
            .lcout(n2516),
            .ltout(n2516_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_123_LC_7_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_123_LC_7_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_123_LC_7_18_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_123_LC_7_18_1 (
            .in0(N__30973),
            .in1(N__31547),
            .in2(N__30946),
            .in3(N__30943),
            .lcout(),
            .ltout(n13816_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12937_4_lut_LC_7_18_2.C_ON=1'b0;
    defparam i12937_4_lut_LC_7_18_2.SEQ_MODE=4'b0000;
    defparam i12937_4_lut_LC_7_18_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12937_4_lut_LC_7_18_2 (
            .in0(N__31169),
            .in1(N__34548),
            .in2(N__30934),
            .in3(N__30927),
            .lcout(n2544),
            .ltout(n2544_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_7_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_7_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_7_18_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1710_3_lut_LC_7_18_3 (
            .in0(N__30916),
            .in1(_gnd_net_),
            .in2(N__30907),
            .in3(N__31548),
            .lcout(n2614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_7_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_7_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_7_18_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1707_3_lut_LC_7_18_4 (
            .in0(N__31170),
            .in1(_gnd_net_),
            .in2(N__30904),
            .in3(N__38862),
            .lcout(n2611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1652_rep_61_3_lut_LC_7_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1652_rep_61_3_lut_LC_7_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1652_rep_61_3_lut_LC_7_18_5.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1652_rep_61_3_lut_LC_7_18_5 (
            .in0(N__30892),
            .in1(N__30859),
            .in2(N__35106),
            .in3(_gnd_net_),
            .lcout(n2524),
            .ltout(n2524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12344_3_lut_LC_7_18_6.C_ON=1'b0;
    defparam i12344_3_lut_LC_7_18_6.SEQ_MODE=4'b0000;
    defparam i12344_3_lut_LC_7_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12344_3_lut_LC_7_18_6 (
            .in0(_gnd_net_),
            .in1(N__31321),
            .in2(N__31312),
            .in3(N__38861),
            .lcout(n2623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12377_3_lut_LC_7_18_7.C_ON=1'b0;
    defparam i12377_3_lut_LC_7_18_7.SEQ_MODE=4'b0000;
    defparam i12377_3_lut_LC_7_18_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12377_3_lut_LC_7_18_7 (
            .in0(_gnd_net_),
            .in1(N__32421),
            .in2(N__31309),
            .in3(N__34930),
            .lcout(n2423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_7_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_7_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_7_19_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1729_3_lut_LC_7_19_0 (
            .in0(N__31270),
            .in1(N__32775),
            .in2(_gnd_net_),
            .in3(N__38869),
            .lcout(n2633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_7_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_7_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1586_3_lut_LC_7_19_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1586_3_lut_LC_7_19_1 (
            .in0(_gnd_net_),
            .in1(N__32358),
            .in2(N__31258),
            .in3(N__34919),
            .lcout(n2426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_7_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_7_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_7_19_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1640_3_lut_LC_7_19_2 (
            .in0(_gnd_net_),
            .in1(N__31207),
            .in2(N__31201),
            .in3(N__35097),
            .lcout(n2512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_7_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_7_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_7_19_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1580_3_lut_LC_7_19_3 (
            .in0(_gnd_net_),
            .in1(N__32451),
            .in2(N__31156),
            .in3(N__34920),
            .lcout(n2420),
            .ltout(n2420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_7_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_7_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_7_19_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1647_3_lut_LC_7_19_4 (
            .in0(_gnd_net_),
            .in1(N__31117),
            .in2(N__31111),
            .in3(N__35093),
            .lcout(n2519),
            .ltout(n2519_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_7_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_7_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_7_19_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1714_3_lut_LC_7_19_5 (
            .in0(N__38870),
            .in1(_gnd_net_),
            .in2(N__31084),
            .in3(N__31081),
            .lcout(n2618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_7_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_7_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_7_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1727_3_lut_LC_7_19_6 (
            .in0(_gnd_net_),
            .in1(N__31623),
            .in2(N__31603),
            .in3(N__38868),
            .lcout(n2631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_7_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_7_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_7_19_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1643_3_lut_LC_7_19_7 (
            .in0(_gnd_net_),
            .in1(N__31588),
            .in2(N__35109),
            .in3(N__31582),
            .lcout(n2515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_7_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_7_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_2_lut_LC_7_20_0 (
            .in0(_gnd_net_),
            .in1(N__32148),
            .in2(_gnd_net_),
            .in3(N__31525),
            .lcout(n2301),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(n12276),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_7_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_7_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_7_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_3_lut_LC_7_20_1 (
            .in0(_gnd_net_),
            .in1(N__53359),
            .in2(N__31522),
            .in3(N__31483),
            .lcout(n2300),
            .ltout(),
            .carryin(n12276),
            .carryout(n12277),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_7_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_7_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_7_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_4_lut_LC_7_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31480),
            .in3(N__31444),
            .lcout(n2299),
            .ltout(),
            .carryin(n12277),
            .carryout(n12278),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_7_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_7_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_7_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_5_lut_LC_7_20_3 (
            .in0(_gnd_net_),
            .in1(N__53360),
            .in2(N__31441),
            .in3(N__31405),
            .lcout(n2298),
            .ltout(),
            .carryin(n12278),
            .carryout(n12279),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_7_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_7_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_7_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_6_lut_LC_7_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31402),
            .in3(N__31366),
            .lcout(n2297),
            .ltout(),
            .carryin(n12279),
            .carryout(n12280),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_7_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_7_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_7_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_7_lut_LC_7_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31363),
            .in3(N__31324),
            .lcout(n2296),
            .ltout(),
            .carryin(n12280),
            .carryout(n12281),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_7_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_7_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_7_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_8_lut_LC_7_20_6 (
            .in0(_gnd_net_),
            .in1(N__53362),
            .in2(N__32511),
            .in3(N__31843),
            .lcout(n2295),
            .ltout(),
            .carryin(n12281),
            .carryout(n12282),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_7_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_7_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_7_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_9_lut_LC_7_20_7 (
            .in0(_gnd_net_),
            .in1(N__53361),
            .in2(N__31840),
            .in3(N__31804),
            .lcout(n2294),
            .ltout(),
            .carryin(n12282),
            .carryout(n12283),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_7_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_7_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_7_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_10_lut_LC_7_21_0 (
            .in0(_gnd_net_),
            .in1(N__54678),
            .in2(N__31800),
            .in3(N__31771),
            .lcout(n2293),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(n12284),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_7_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_7_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_7_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_11_lut_LC_7_21_1 (
            .in0(_gnd_net_),
            .in1(N__54240),
            .in2(N__31899),
            .in3(N__31768),
            .lcout(n2292),
            .ltout(),
            .carryin(n12284),
            .carryout(n12285),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_7_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_7_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_7_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_12_lut_LC_7_21_2 (
            .in0(_gnd_net_),
            .in1(N__54679),
            .in2(N__31866),
            .in3(N__31765),
            .lcout(n2291),
            .ltout(),
            .carryin(n12285),
            .carryout(n12286),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_7_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_7_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_7_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_13_lut_LC_7_21_3 (
            .in0(_gnd_net_),
            .in1(N__54241),
            .in2(N__31762),
            .in3(N__31738),
            .lcout(n2290_adj_604),
            .ltout(),
            .carryin(n12286),
            .carryout(n12287),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_7_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_7_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_7_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_14_lut_LC_7_21_4 (
            .in0(_gnd_net_),
            .in1(N__31735),
            .in2(N__54727),
            .in3(N__31705),
            .lcout(n2289_adj_603),
            .ltout(),
            .carryin(n12287),
            .carryout(n12288),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_7_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_7_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_7_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_15_lut_LC_7_21_5 (
            .in0(_gnd_net_),
            .in1(N__31702),
            .in2(N__54996),
            .in3(N__31666),
            .lcout(n2288_adj_602),
            .ltout(),
            .carryin(n12288),
            .carryout(n12289),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_7_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_7_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_7_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_16_lut_LC_7_21_6 (
            .in0(_gnd_net_),
            .in1(N__31663),
            .in2(N__54728),
            .in3(N__32131),
            .lcout(n2287_adj_601),
            .ltout(),
            .carryin(n12289),
            .carryout(n12290),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_7_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_7_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_7_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_17_lut_LC_7_21_7 (
            .in0(_gnd_net_),
            .in1(N__32128),
            .in2(N__54997),
            .in3(N__32098),
            .lcout(n2286_adj_600),
            .ltout(),
            .carryin(n12290),
            .carryout(n12291),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_7_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_7_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_7_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_18_lut_LC_7_22_0 (
            .in0(_gnd_net_),
            .in1(N__32095),
            .in2(N__54077),
            .in3(N__32056),
            .lcout(n2285_adj_599),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(n12292),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_7_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_7_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_7_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_19_lut_LC_7_22_1 (
            .in0(_gnd_net_),
            .in1(N__53672),
            .in2(N__39196),
            .in3(N__32053),
            .lcout(n2284),
            .ltout(),
            .carryin(n12292),
            .carryout(n12293),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_7_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_7_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_7_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_20_lut_LC_7_22_2 (
            .in0(_gnd_net_),
            .in1(N__32050),
            .in2(N__54078),
            .in3(N__32011),
            .lcout(n2283),
            .ltout(),
            .carryin(n12293),
            .carryout(n12294),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_7_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_7_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_7_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_21_lut_LC_7_22_3 (
            .in0(_gnd_net_),
            .in1(N__32007),
            .in2(N__55161),
            .in3(N__31957),
            .lcout(n2282),
            .ltout(),
            .carryin(n12294),
            .carryout(n12295),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_7_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_7_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_7_22_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1503_22_lut_LC_7_22_4 (
            .in0(N__53676),
            .in1(N__31954),
            .in2(N__34794),
            .in3(N__31924),
            .lcout(n2313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12376_3_lut_LC_7_22_5.C_ON=1'b0;
    defparam i12376_3_lut_LC_7_22_5.SEQ_MODE=4'b0000;
    defparam i12376_3_lut_LC_7_22_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12376_3_lut_LC_7_22_5 (
            .in0(_gnd_net_),
            .in1(N__31900),
            .in2(N__31876),
            .in3(N__39139),
            .lcout(n2324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_7_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_7_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_7_22_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1515_3_lut_LC_7_22_6 (
            .in0(_gnd_net_),
            .in1(N__31867),
            .in2(N__39150),
            .in3(N__31849),
            .lcout(n2323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_7_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_7_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1519_3_lut_LC_7_22_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1519_3_lut_LC_7_22_7 (
            .in0(_gnd_net_),
            .in1(N__32521),
            .in2(N__32512),
            .in3(N__39138),
            .lcout(n2327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_7_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_7_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_7_23_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_7_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32471),
            .lcout(n31_adj_655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_23_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_23_1 (
            .in0(N__37776),
            .in1(N__32845),
            .in2(_gnd_net_),
            .in3(N__39548),
            .lcout(n313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_108_LC_7_23_2.C_ON=1'b0;
    defparam i1_4_lut_adj_108_LC_7_23_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_108_LC_7_23_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_108_LC_7_23_2 (
            .in0(N__32447),
            .in1(N__32411),
            .in2(N__32395),
            .in3(N__32348),
            .lcout(n14008),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_23_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_23_3 (
            .in0(N__32860),
            .in1(N__39549),
            .in2(_gnd_net_),
            .in3(N__32733),
            .lcout(n314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_107_LC_7_23_5.C_ON=1'b0;
    defparam i1_4_lut_adj_107_LC_7_23_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_107_LC_7_23_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_107_LC_7_23_5 (
            .in0(N__32318),
            .in1(N__32298),
            .in2(N__32277),
            .in3(N__32225),
            .lcout(n14006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_7_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_7_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_7_23_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i4_3_lut_LC_7_23_6 (
            .in0(N__39550),
            .in1(N__32896),
            .in2(_gnd_net_),
            .in3(N__32201),
            .lcout(n316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_23_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_23_7 (
            .in0(N__33061),
            .in1(N__39547),
            .in2(_gnd_net_),
            .in3(N__32180),
            .lcout(n308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_24_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_24_0 (
            .in0(N__39518),
            .in1(N__32947),
            .in2(_gnd_net_),
            .in3(N__32586),
            .lcout(n318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_1 (
            .in0(N__32812),
            .in1(N__32795),
            .in2(_gnd_net_),
            .in3(N__39517),
            .lcout(n311),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_7_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_7_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_7_24_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_7_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32732),
            .lcout(n28_adj_652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_7_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_7_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_7_24_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i16_3_lut_LC_7_24_3 (
            .in0(N__32992),
            .in1(N__39516),
            .in2(_gnd_net_),
            .in3(N__32714),
            .lcout(n304),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_7_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_7_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_7_24_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_7_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37976),
            .lcout(n26_adj_650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_109_LC_7_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_109_LC_7_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_109_LC_7_24_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_109_LC_7_24_5 (
            .in0(N__32662),
            .in1(N__32641),
            .in2(N__32620),
            .in3(N__32611),
            .lcout(n14014),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_7_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_7_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_7_24_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_7_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32585),
            .lcout(n32_adj_656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_7_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_7_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_7_24_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_7_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32564),
            .lcout(n33_adj_657),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_7_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_7_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_7_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_7_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32548),
            .in3(N__32524),
            .lcout(n33),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(n12575),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_7_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_7_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_7_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_7_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32956),
            .in3(N__32941),
            .lcout(n32),
            .ltout(),
            .carryin(n12575),
            .carryout(n12576),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_7_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_7_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_7_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_7_25_2 (
            .in0(_gnd_net_),
            .in1(N__32938),
            .in2(_gnd_net_),
            .in3(N__32914),
            .lcout(n31),
            .ltout(),
            .carryin(n12576),
            .carryout(n12577),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_7_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_7_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_7_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_7_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32911),
            .in3(N__32887),
            .lcout(n30),
            .ltout(),
            .carryin(n12577),
            .carryout(n12578),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_7_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_7_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_7_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_7_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32884),
            .in3(N__32872),
            .lcout(n29),
            .ltout(),
            .carryin(n12578),
            .carryout(n12579),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_7_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_7_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_7_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_7_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32869),
            .in3(N__32848),
            .lcout(n28),
            .ltout(),
            .carryin(n12579),
            .carryout(n12580),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_7_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_7_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_7_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_7_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37753),
            .in3(N__32836),
            .lcout(n27),
            .ltout(),
            .carryin(n12580),
            .carryout(n12581),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_7_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_7_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_7_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_7_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32833),
            .in3(N__32824),
            .lcout(n26),
            .ltout(),
            .carryin(n12581),
            .carryout(n12582),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_7_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_7_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_7_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_7_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32821),
            .in3(N__32803),
            .lcout(n25),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(n12583),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_7_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_7_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_7_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_7_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33103),
            .in3(N__33094),
            .lcout(n24),
            .ltout(),
            .carryin(n12583),
            .carryout(n12584),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_7_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_7_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_7_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_7_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33091),
            .in3(N__33076),
            .lcout(n23),
            .ltout(),
            .carryin(n12584),
            .carryout(n12585),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_7_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_7_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_7_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_7_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33073),
            .in3(N__33052),
            .lcout(n22),
            .ltout(),
            .carryin(n12585),
            .carryout(n12586),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_7_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_7_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_7_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_7_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33049),
            .in3(N__33025),
            .lcout(n21),
            .ltout(),
            .carryin(n12586),
            .carryout(n12587),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_7_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_7_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_7_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_7_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38278),
            .in3(N__33013),
            .lcout(n20),
            .ltout(),
            .carryin(n12587),
            .carryout(n12588),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_7_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_7_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_7_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_7_26_6 (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(_gnd_net_),
            .in3(N__33004),
            .lcout(n19),
            .ltout(),
            .carryin(n12588),
            .carryout(n12589),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_7_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_7_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_7_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_7_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33001),
            .in3(N__32983),
            .lcout(n18),
            .ltout(),
            .carryin(n12589),
            .carryout(n12590),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_7_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_7_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_7_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_7_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32980),
            .in3(N__32959),
            .lcout(n17),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(n12591),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_7_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_7_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_7_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_7_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33337),
            .in3(N__33316),
            .lcout(n16),
            .ltout(),
            .carryin(n12591),
            .carryout(n12592),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_7_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_7_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_7_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_7_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33313),
            .in3(N__33286),
            .lcout(n15),
            .ltout(),
            .carryin(n12592),
            .carryout(n12593),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_7_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_7_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_7_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_7_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33283),
            .in3(N__33262),
            .lcout(n14),
            .ltout(),
            .carryin(n12593),
            .carryout(n12594),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_7_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_7_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_7_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_7_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33259),
            .in3(N__33232),
            .lcout(n13),
            .ltout(),
            .carryin(n12594),
            .carryout(n12595),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_7_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_7_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_7_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_7_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33229),
            .in3(N__33202),
            .lcout(n12),
            .ltout(),
            .carryin(n12595),
            .carryout(n12596),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_7_27_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_7_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_7_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_7_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33199),
            .in3(N__33172),
            .lcout(n11),
            .ltout(),
            .carryin(n12596),
            .carryout(n12597),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_7_27_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_7_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_7_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_7_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33169),
            .in3(N__33136),
            .lcout(n10),
            .ltout(),
            .carryin(n12597),
            .carryout(n12598),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_7_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_7_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_7_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_7_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33133),
            .in3(N__33106),
            .lcout(n9),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(n12599),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_7_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_7_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_7_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_7_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33550),
            .in3(N__33535),
            .lcout(n8),
            .ltout(),
            .carryin(n12599),
            .carryout(n12600),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_7_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_7_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_7_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_7_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33532),
            .in3(N__33514),
            .lcout(n7),
            .ltout(),
            .carryin(n12600),
            .carryout(n12601),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_7_28_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_7_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_7_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_7_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33511),
            .in3(N__33475),
            .lcout(n6),
            .ltout(),
            .carryin(n12601),
            .carryout(n12602),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_7_28_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_7_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_7_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_7_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38233),
            .in3(N__33445),
            .lcout(n5),
            .ltout(),
            .carryin(n12602),
            .carryout(n12603),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_7_28_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_7_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_7_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_7_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33442),
            .in3(N__33406),
            .lcout(n4),
            .ltout(),
            .carryin(n12603),
            .carryout(n12604),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_7_28_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_7_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_7_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_7_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33403),
            .in3(N__33373),
            .lcout(n3_adj_567),
            .ltout(),
            .carryin(n12604),
            .carryout(n12605),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_7_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_7_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_7_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_7_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36438),
            .in3(N__33370),
            .lcout(n2_adj_568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_7_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_7_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_7_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_2_lut_LC_7_29_0 (
            .in0(_gnd_net_),
            .in1(N__36260),
            .in2(_gnd_net_),
            .in3(N__33340),
            .lcout(n901),
            .ltout(),
            .carryin(bfn_7_29_0_),
            .carryout(n12101),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_7_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_7_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_7_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_3_lut_LC_7_29_1 (
            .in0(_gnd_net_),
            .in1(N__55172),
            .in2(N__33573),
            .in3(N__33712),
            .lcout(n900),
            .ltout(),
            .carryin(n12101),
            .carryout(n12102),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_7_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_7_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_7_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_4_lut_LC_7_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33709),
            .in3(N__33670),
            .lcout(n899),
            .ltout(),
            .carryin(n12102),
            .carryout(n12103),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_7_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_7_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_7_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_5_lut_LC_7_29_3 (
            .in0(_gnd_net_),
            .in1(N__55173),
            .in2(N__34251),
            .in3(N__33667),
            .lcout(n898),
            .ltout(),
            .carryin(n12103),
            .carryout(n12104),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_7_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_7_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_7_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_6_lut_LC_7_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33664),
            .in3(N__33628),
            .lcout(n897),
            .ltout(),
            .carryin(n12104),
            .carryout(n12105),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_7_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_7_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_7_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_7_lut_LC_7_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33625),
            .in3(N__33601),
            .lcout(n896),
            .ltout(),
            .carryin(n12105),
            .carryout(n12106),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_7_29_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_7_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_7_29_6.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_565_8_lut_LC_7_29_6 (
            .in0(N__55174),
            .in1(N__33597),
            .in2(N__34225),
            .in3(N__33583),
            .lcout(n927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i572_3_lut_LC_7_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_7_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_7_29_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i572_3_lut_LC_7_29_7 (
            .in0(_gnd_net_),
            .in1(N__33580),
            .in2(N__33574),
            .in3(N__34219),
            .lcout(n932),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_7_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_7_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_7_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_2_lut_LC_7_30_0 (
            .in0(_gnd_net_),
            .in1(N__34065),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(n1001),
            .ltout(),
            .carryin(bfn_7_30_0_),
            .carryout(n12107),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_7_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_7_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_7_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_3_lut_LC_7_30_1 (
            .in0(_gnd_net_),
            .in1(N__54594),
            .in2(N__34087),
            .in3(N__33820),
            .lcout(n1000),
            .ltout(),
            .carryin(n12107),
            .carryout(n12108),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_7_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_7_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_7_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_4_lut_LC_7_30_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33738),
            .in3(N__33817),
            .lcout(n999),
            .ltout(),
            .carryin(n12108),
            .carryout(n12109),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_7_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_7_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_7_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_5_lut_LC_7_30_3 (
            .in0(_gnd_net_),
            .in1(N__54595),
            .in2(N__34039),
            .in3(N__33814),
            .lcout(n998),
            .ltout(),
            .carryin(n12109),
            .carryout(n12110),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_7_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_7_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_7_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_6_lut_LC_7_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34191),
            .in3(N__33811),
            .lcout(n997),
            .ltout(),
            .carryin(n12110),
            .carryout(n12111),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_7_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_7_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_7_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_7_lut_LC_7_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34170),
            .in3(N__33796),
            .lcout(n996),
            .ltout(),
            .carryin(n12111),
            .carryout(n12112),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_7_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_7_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_7_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_8_lut_LC_7_30_6 (
            .in0(_gnd_net_),
            .in1(N__54596),
            .in2(N__34128),
            .in3(N__33784),
            .lcout(n995),
            .ltout(),
            .carryin(n12112),
            .carryout(n12113),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_7_30_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_7_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_7_30_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_632_9_lut_LC_7_30_7 (
            .in0(N__54597),
            .in1(N__34014),
            .in2(N__34147),
            .in3(N__33781),
            .lcout(n1026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i637_3_lut_LC_7_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_7_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_7_31_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i637_3_lut_LC_7_31_0 (
            .in0(_gnd_net_),
            .in1(N__33751),
            .in2(N__34192),
            .in3(N__34004),
            .lcout(n1029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i639_3_lut_LC_7_31_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_7_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_7_31_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i639_3_lut_LC_7_31_1 (
            .in0(_gnd_net_),
            .in1(N__33745),
            .in2(N__34016),
            .in3(N__33739),
            .lcout(n1031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i570_3_lut_LC_7_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_7_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_7_31_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i570_3_lut_LC_7_31_2 (
            .in0(_gnd_net_),
            .in1(N__34264),
            .in2(N__34255),
            .in3(N__34223),
            .lcout(n930),
            .ltout(n930_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_7_31_3.C_ON=1'b0;
    defparam i1_2_lut_LC_7_31_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_7_31_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_LC_7_31_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34174),
            .in3(N__34163),
            .lcout(),
            .ltout(n13726_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_7_31_4.C_ON=1'b0;
    defparam i1_4_lut_LC_7_31_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_7_31_4.LUT_INIT=16'b1111111011101110;
    LogicCell40 i1_4_lut_LC_7_31_4 (
            .in0(N__34146),
            .in1(N__34121),
            .in2(N__34105),
            .in3(N__34102),
            .lcout(n960),
            .ltout(n960_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i640_3_lut_LC_7_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_7_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_7_31_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i640_3_lut_LC_7_31_5 (
            .in0(N__34096),
            .in1(_gnd_net_),
            .in2(N__34090),
            .in3(N__34086),
            .lcout(n1032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i641_3_lut_LC_7_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_7_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_7_31_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i641_3_lut_LC_7_31_6 (
            .in0(N__34066),
            .in1(_gnd_net_),
            .in2(N__34048),
            .in3(N__34003),
            .lcout(n1033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i638_3_lut_LC_7_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_7_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_7_31_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i638_3_lut_LC_7_31_7 (
            .in0(_gnd_net_),
            .in1(N__34038),
            .in2(N__34017),
            .in3(N__33976),
            .lcout(n1030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9932_3_lut_LC_7_32_4.C_ON=1'b0;
    defparam i9932_3_lut_LC_7_32_4.SEQ_MODE=4'b0000;
    defparam i9932_3_lut_LC_7_32_4.LUT_INIT=16'b1100110011000000;
    LogicCell40 i9932_3_lut_LC_7_32_4 (
            .in0(_gnd_net_),
            .in1(N__33965),
            .in2(N__33949),
            .in3(N__33920),
            .lcout(),
            .ltout(n11646_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_27_LC_7_32_5.C_ON=1'b0;
    defparam i1_4_lut_adj_27_LC_7_32_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_27_LC_7_32_5.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_27_LC_7_32_5 (
            .in0(N__33890),
            .in1(N__33869),
            .in2(N__33853),
            .in3(N__33842),
            .lcout(n13323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i1_LC_7_32_7.C_ON=1'b0;
    defparam commutation_state_i1_LC_7_32_7.SEQ_MODE=4'b1000;
    defparam commutation_state_i1_LC_7_32_7.LUT_INIT=16'b1011001100010000;
    LogicCell40 commutation_state_i1_LC_7_32_7 (
            .in0(N__38088),
            .in1(N__38155),
            .in2(N__56353),
            .in3(N__38191),
            .lcout(commutation_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56068),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_9_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_9_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1726_3_lut_LC_9_17_0 (
            .in0(N__34462),
            .in1(N__34432),
            .in2(_gnd_net_),
            .in3(N__38936),
            .lcout(n2630),
            .ltout(n2630_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_60_LC_9_17_1.C_ON=1'b0;
    defparam i1_4_lut_adj_60_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_60_LC_9_17_1.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_60_LC_9_17_1 (
            .in0(N__37118),
            .in1(N__38674),
            .in2(N__34420),
            .in3(N__34363),
            .lcout(),
            .ltout(n14288_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_61_LC_9_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_61_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_61_LC_9_17_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_61_LC_9_17_2 (
            .in0(N__37472),
            .in1(N__38603),
            .in2(N__34417),
            .in3(N__37190),
            .lcout(n14294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_9_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_9_17_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1722_3_lut_LC_9_17_4 (
            .in0(N__34413),
            .in1(_gnd_net_),
            .in2(N__34393),
            .in3(N__38935),
            .lcout(n2626),
            .ltout(n2626_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_58_LC_9_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_58_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_58_LC_9_17_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_58_LC_9_17_5 (
            .in0(N__34638),
            .in1(N__34715),
            .in2(N__34378),
            .in3(N__34375),
            .lcout(),
            .ltout(n14280_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_59_LC_9_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_59_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_59_LC_9_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_59_LC_9_17_6 (
            .in0(N__37292),
            .in1(N__37019),
            .in2(N__34366),
            .in3(N__37353),
            .lcout(n14286),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_9_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_9_18_0.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1717_3_lut_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(N__38908),
            .in2(N__34357),
            .in3(N__34321),
            .lcout(n2621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_9_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_9_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_9_18_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1725_3_lut_LC_9_18_1 (
            .in0(_gnd_net_),
            .in1(N__34309),
            .in2(N__38932),
            .in3(N__34296),
            .lcout(n2629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_9_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_9_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_9_18_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1715_3_lut_LC_9_18_2 (
            .in0(_gnd_net_),
            .in1(N__34608),
            .in2(N__34576),
            .in3(N__38909),
            .lcout(n2619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_9_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_9_18_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1708_3_lut_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(N__34561),
            .in2(N__38933),
            .in3(N__34549),
            .lcout(n2612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12373_3_lut_LC_9_18_4.C_ON=1'b0;
    defparam i12373_3_lut_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam i12373_3_lut_LC_9_18_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 i12373_3_lut_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(N__34693),
            .in2(N__42429),
            .in3(N__34717),
            .lcout(n2721),
            .ltout(n2721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12303_3_lut_LC_9_18_5.C_ON=1'b0;
    defparam i12303_3_lut_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam i12303_3_lut_LC_9_18_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12303_3_lut_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(N__40243),
            .in2(N__34522),
            .in3(N__47630),
            .lcout(n2820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1721_rep_13_3_lut_LC_9_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1721_rep_13_3_lut_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1721_rep_13_3_lut_LC_9_18_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1721_rep_13_3_lut_LC_9_18_6 (
            .in0(_gnd_net_),
            .in1(N__34519),
            .in2(N__34489),
            .in3(N__38907),
            .lcout(n2625),
            .ltout(n2625_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12348_3_lut_LC_9_18_7.C_ON=1'b0;
    defparam i12348_3_lut_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam i12348_3_lut_LC_9_18_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12348_3_lut_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(N__34627),
            .in2(N__34474),
            .in3(N__42391),
            .lcout(n2724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_9_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_9_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_9_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_2_lut_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(N__38775),
            .in2(_gnd_net_),
            .in3(N__34471),
            .lcout(n2701),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(n12362),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_9_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_9_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_9_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_3_lut_LC_9_19_1 (
            .in0(_gnd_net_),
            .in1(N__53482),
            .in2(N__38736),
            .in3(N__34468),
            .lcout(n2700),
            .ltout(),
            .carryin(n12362),
            .carryout(n12363),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_9_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_9_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_9_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_4_lut_LC_9_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38794),
            .in3(N__34465),
            .lcout(n2699),
            .ltout(),
            .carryin(n12363),
            .carryout(n12364),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_9_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_9_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_5_lut_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(N__53483),
            .in2(N__38703),
            .in3(N__34660),
            .lcout(n2698),
            .ltout(),
            .carryin(n12364),
            .carryout(n12365),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_9_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_9_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_9_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_6_lut_LC_9_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37090),
            .in3(N__34657),
            .lcout(n2697),
            .ltout(),
            .carryin(n12365),
            .carryout(n12366),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_9_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_9_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_9_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_7_lut_LC_9_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37123),
            .in3(N__34654),
            .lcout(n2696),
            .ltout(),
            .carryin(n12366),
            .carryout(n12367),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_9_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_9_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_8_lut_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(N__53485),
            .in2(N__37054),
            .in3(N__34651),
            .lcout(n2695),
            .ltout(),
            .carryin(n12367),
            .carryout(n12368),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_9_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_9_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_9_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_9_lut_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(N__53484),
            .in2(N__37441),
            .in3(N__34648),
            .lcout(n2694),
            .ltout(),
            .carryin(n12368),
            .carryout(n12369),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_9_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_9_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_10_lut_LC_9_20_0 (
            .in0(_gnd_net_),
            .in1(N__37144),
            .in2(N__53831),
            .in3(N__34645),
            .lcout(n2693),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(n12370),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_9_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_9_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_9_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_11_lut_LC_9_20_1 (
            .in0(_gnd_net_),
            .in1(N__34642),
            .in2(N__53833),
            .in3(N__34618),
            .lcout(n2692),
            .ltout(),
            .carryin(n12370),
            .carryout(n12371),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_9_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_9_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_9_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_12_lut_LC_9_20_2 (
            .in0(_gnd_net_),
            .in1(N__53496),
            .in2(N__38643),
            .in3(N__34615),
            .lcout(n2691),
            .ltout(),
            .carryin(n12371),
            .carryout(n12372),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_9_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_9_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_9_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_13_lut_LC_9_20_3 (
            .in0(_gnd_net_),
            .in1(N__53489),
            .in2(N__39268),
            .in3(N__34612),
            .lcout(n2690),
            .ltout(),
            .carryin(n12372),
            .carryout(n12373),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_9_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_9_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_9_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_14_lut_LC_9_20_4 (
            .in0(_gnd_net_),
            .in1(N__34716),
            .in2(N__53832),
            .in3(N__34684),
            .lcout(n2689),
            .ltout(),
            .carryin(n12373),
            .carryout(n12374),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_9_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_9_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_9_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_15_lut_LC_9_20_5 (
            .in0(_gnd_net_),
            .in1(N__37297),
            .in2(N__53834),
            .in3(N__34681),
            .lcout(n2688),
            .ltout(),
            .carryin(n12374),
            .carryout(n12375),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_9_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_9_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_9_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_16_lut_LC_9_20_6 (
            .in0(_gnd_net_),
            .in1(N__53500),
            .in2(N__37360),
            .in3(N__34678),
            .lcout(n2687),
            .ltout(),
            .carryin(n12375),
            .carryout(n12376),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_9_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_9_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_9_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_17_lut_LC_9_20_7 (
            .in0(_gnd_net_),
            .in1(N__37026),
            .in2(N__53835),
            .in3(N__34675),
            .lcout(n2686),
            .ltout(),
            .carryin(n12376),
            .carryout(n12377),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_9_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_9_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_9_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_18_lut_LC_9_21_0 (
            .in0(_gnd_net_),
            .in1(N__37191),
            .in2(N__53836),
            .in3(N__34672),
            .lcout(n2685),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(n12378),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_9_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_9_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_9_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_19_lut_LC_9_21_1 (
            .in0(_gnd_net_),
            .in1(N__38610),
            .in2(N__53869),
            .in3(N__34669),
            .lcout(n2684),
            .ltout(),
            .carryin(n12378),
            .carryout(n12379),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_9_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_9_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_9_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_20_lut_LC_9_21_2 (
            .in0(_gnd_net_),
            .in1(N__53550),
            .in2(N__37483),
            .in3(N__34666),
            .lcout(n2683),
            .ltout(),
            .carryin(n12379),
            .carryout(n12380),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_9_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_9_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_9_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_21_lut_LC_9_21_3 (
            .in0(_gnd_net_),
            .in1(N__38470),
            .in2(N__53870),
            .in3(N__34663),
            .lcout(n2682),
            .ltout(),
            .carryin(n12380),
            .carryout(n12381),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_9_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_9_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_9_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_22_lut_LC_9_21_4 (
            .in0(_gnd_net_),
            .in1(N__37245),
            .in2(N__53837),
            .in3(N__34732),
            .lcout(n2681),
            .ltout(),
            .carryin(n12381),
            .carryout(n12382),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_9_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_9_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_9_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_23_lut_LC_9_21_5 (
            .in0(_gnd_net_),
            .in1(N__53510),
            .in2(N__38557),
            .in3(N__34729),
            .lcout(n2680),
            .ltout(),
            .carryin(n12382),
            .carryout(n12383),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_9_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_9_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_9_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_24_lut_LC_9_21_6 (
            .in0(_gnd_net_),
            .in1(N__42474),
            .in2(N__53838),
            .in3(N__34726),
            .lcout(n2679),
            .ltout(),
            .carryin(n12383),
            .carryout(n12384),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_9_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_9_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_9_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_25_lut_LC_9_21_7 (
            .in0(_gnd_net_),
            .in1(N__38512),
            .in2(N__53871),
            .in3(N__34723),
            .lcout(n2678),
            .ltout(),
            .carryin(n12384),
            .carryout(n12385),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_9_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_9_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_9_22_0.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1771_26_lut_LC_9_22_0 (
            .in0(N__53523),
            .in1(N__37330),
            .in2(N__35184),
            .in3(N__34720),
            .lcout(n2709),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12965_1_lut_LC_9_22_1.C_ON=1'b0;
    defparam i12965_1_lut_LC_9_22_1.SEQ_MODE=4'b0000;
    defparam i12965_1_lut_LC_9_22_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12965_1_lut_LC_9_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42443),
            .lcout(n15437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_9_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_9_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_9_22_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1841_3_lut_LC_9_22_3 (
            .in0(N__47637),
            .in1(_gnd_net_),
            .in2(N__41572),
            .in3(N__40441),
            .lcout(n2809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_9_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_9_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_9_22_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2067_3_lut_LC_9_22_4 (
            .in0(_gnd_net_),
            .in1(N__44788),
            .in2(N__44764),
            .in3(N__49063),
            .lcout(n3131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_9_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_9_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_9_22_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2069_3_lut_LC_9_22_5 (
            .in0(_gnd_net_),
            .in1(N__44854),
            .in2(N__49082),
            .in3(N__44892),
            .lcout(n3133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_9_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_9_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_9_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2042_3_lut_LC_9_22_6 (
            .in0(_gnd_net_),
            .in1(N__45543),
            .in2(N__45517),
            .in3(N__49064),
            .lcout(n3106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_9_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_9_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_9_22_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2068_3_lut_LC_9_22_7 (
            .in0(N__44803),
            .in1(_gnd_net_),
            .in2(N__49081),
            .in3(N__44835),
            .lcout(n3132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10035_4_lut_LC_9_23_0.C_ON=1'b0;
    defparam i10035_4_lut_LC_9_23_0.SEQ_MODE=4'b0000;
    defparam i10035_4_lut_LC_9_23_0.LUT_INIT=16'b1111101011101010;
    LogicCell40 i10035_4_lut_LC_9_23_0 (
            .in0(N__51011),
            .in1(N__51176),
            .in2(N__51068),
            .in3(N__51110),
            .lcout(),
            .ltout(n11750_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_169_LC_9_23_1.C_ON=1'b0;
    defparam i1_4_lut_adj_169_LC_9_23_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_169_LC_9_23_1.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_169_LC_9_23_1 (
            .in0(N__50978),
            .in1(N__50928),
            .in2(N__34750),
            .in3(N__39637),
            .lcout(),
            .ltout(n13900_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_170_LC_9_23_2.C_ON=1'b0;
    defparam i1_4_lut_adj_170_LC_9_23_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_170_LC_9_23_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_170_LC_9_23_2 (
            .in0(N__52214),
            .in1(N__51588),
            .in2(N__34747),
            .in3(N__51639),
            .lcout(n13906),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_9_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_9_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_9_23_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2136_3_lut_LC_9_23_3 (
            .in0(_gnd_net_),
            .in1(N__51094),
            .in2(N__51117),
            .in3(N__50019),
            .lcout(n3232),
            .ltout(n3232_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9943_3_lut_LC_9_23_4.C_ON=1'b0;
    defparam i9943_3_lut_LC_9_23_4.SEQ_MODE=4'b0000;
    defparam i9943_3_lut_LC_9_23_4.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9943_3_lut_LC_9_23_4 (
            .in0(_gnd_net_),
            .in1(N__42818),
            .in2(N__34744),
            .in3(N__42761),
            .lcout(n11658),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_9_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_9_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_9_23_6.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2134_3_lut_LC_9_23_6 (
            .in0(N__51012),
            .in1(N__50998),
            .in2(N__50070),
            .in3(_gnd_net_),
            .lcout(n3230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_9_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_9_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_9_24_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2129_3_lut_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(N__51556),
            .in2(N__51520),
            .in3(N__50013),
            .lcout(n3225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_171_LC_9_24_1.C_ON=1'b0;
    defparam i1_4_lut_adj_171_LC_9_24_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_171_LC_9_24_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_171_LC_9_24_1 (
            .in0(N__52174),
            .in1(N__52140),
            .in2(N__52093),
            .in3(N__34741),
            .lcout(),
            .ltout(n13912_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12689_4_lut_LC_9_24_2.C_ON=1'b0;
    defparam i12689_4_lut_LC_9_24_2.SEQ_MODE=4'b0000;
    defparam i12689_4_lut_LC_9_24_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12689_4_lut_LC_9_24_2 (
            .in0(N__52040),
            .in1(N__51992),
            .in2(N__34735),
            .in3(N__51930),
            .lcout(n3138),
            .ltout(n3138_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_9_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_9_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_9_24_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i2137_3_lut_LC_9_24_3 (
            .in0(N__51181),
            .in1(_gnd_net_),
            .in2(N__34774),
            .in3(N__51139),
            .lcout(n3233),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_9_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_9_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_9_24_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2135_3_lut_LC_9_24_4 (
            .in0(_gnd_net_),
            .in1(N__51069),
            .in2(N__51040),
            .in3(N__50014),
            .lcout(n3231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_9_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_9_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_9_24_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2110_3_lut_LC_9_24_5 (
            .in0(N__52015),
            .in1(_gnd_net_),
            .in2(N__50069),
            .in3(N__52041),
            .lcout(n3206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_9_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_9_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_9_24_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2133_3_lut_LC_9_24_6 (
            .in0(_gnd_net_),
            .in1(N__50982),
            .in2(N__50950),
            .in3(N__50015),
            .lcout(n3229),
            .ltout(n3229_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_154_LC_9_24_7.C_ON=1'b0;
    defparam i1_4_lut_adj_154_LC_9_24_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_154_LC_9_24_7.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_154_LC_9_24_7 (
            .in0(N__42683),
            .in1(N__43094),
            .in2(N__34771),
            .in3(N__34768),
            .lcout(n13470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i0_LC_9_25_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i0_LC_9_25_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i0_LC_9_25_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i0_LC_9_25_0 (
            .in0(N__37876),
            .in1(N__36406),
            .in2(N__37924),
            .in3(N__34762),
            .lcout(encoder0_position_scaled_0),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(n12552),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i1_LC_9_25_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i1_LC_9_25_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i1_LC_9_25_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i1_LC_9_25_1 (
            .in0(N__43587),
            .in1(N__49618),
            .in2(N__36469),
            .in3(N__34759),
            .lcout(encoder0_position_scaled_1),
            .ltout(),
            .carryin(n12552),
            .carryout(n12553),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i2_LC_9_25_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i2_LC_9_25_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i2_LC_9_25_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i2_LC_9_25_2 (
            .in0(N__51951),
            .in1(N__50032),
            .in2(N__36473),
            .in3(N__34756),
            .lcout(encoder0_position_scaled_2),
            .ltout(),
            .carryin(n12553),
            .carryout(n12554),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i3_LC_9_25_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i3_LC_9_25_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i3_LC_9_25_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i3_LC_9_25_3 (
            .in0(N__45915),
            .in1(N__49080),
            .in2(N__36470),
            .in3(N__34753),
            .lcout(encoder0_position_scaled_3),
            .ltout(),
            .carryin(n12554),
            .carryout(n12555),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i4_LC_9_25_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i4_LC_9_25_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i4_LC_9_25_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i4_LC_9_25_4 (
            .in0(N__39763),
            .in1(N__43009),
            .in2(N__36474),
            .in3(N__35197),
            .lcout(encoder0_position_scaled_4),
            .ltout(),
            .carryin(n12555),
            .carryout(n12556),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i5_LC_9_25_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i5_LC_9_25_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i5_LC_9_25_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i5_LC_9_25_5 (
            .in0(N__49201),
            .in1(N__49374),
            .in2(N__36471),
            .in3(N__35194),
            .lcout(encoder0_position_scaled_5),
            .ltout(),
            .carryin(n12556),
            .carryout(n12557),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i6_LC_9_25_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i6_LC_9_25_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i6_LC_9_25_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i6_LC_9_25_6 (
            .in0(N__42283),
            .in1(N__36416),
            .in2(N__47644),
            .in3(N__35191),
            .lcout(encoder0_position_scaled_6),
            .ltout(),
            .carryin(n12557),
            .carryout(n12558),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i7_LC_9_25_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i7_LC_9_25_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i7_LC_9_25_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i7_LC_9_25_7 (
            .in0(N__35188),
            .in1(N__42448),
            .in2(N__36472),
            .in3(N__35167),
            .lcout(encoder0_position_scaled_7),
            .ltout(),
            .carryin(n12558),
            .carryout(n12559),
            .clk(N__56055),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i8_LC_9_26_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i8_LC_9_26_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i8_LC_9_26_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i8_LC_9_26_0 (
            .in0(N__35164),
            .in1(N__38944),
            .in2(N__36475),
            .in3(N__35140),
            .lcout(encoder0_position_scaled_8),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(n12560),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i9_LC_9_26_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i9_LC_9_26_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i9_LC_9_26_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i9_LC_9_26_1 (
            .in0(N__35137),
            .in1(N__35113),
            .in2(N__36479),
            .in3(N__34960),
            .lcout(encoder0_position_scaled_9),
            .ltout(),
            .carryin(n12560),
            .carryout(n12561),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i10_LC_9_26_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i10_LC_9_26_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i10_LC_9_26_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i10_LC_9_26_2 (
            .in0(N__34957),
            .in1(N__34939),
            .in2(N__36476),
            .in3(N__34801),
            .lcout(encoder0_position_scaled_10),
            .ltout(),
            .carryin(n12561),
            .carryout(n12562),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i11_LC_9_26_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i11_LC_9_26_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i11_LC_9_26_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i11_LC_9_26_3 (
            .in0(N__34798),
            .in1(N__39151),
            .in2(N__36480),
            .in3(N__34777),
            .lcout(encoder0_position_scaled_11),
            .ltout(),
            .carryin(n12562),
            .carryout(n12563),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i12_LC_9_26_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i12_LC_9_26_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i12_LC_9_26_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i12_LC_9_26_4 (
            .in0(N__36235),
            .in1(N__36211),
            .in2(N__36477),
            .in3(N__36076),
            .lcout(encoder0_position_scaled_12),
            .ltout(),
            .carryin(n12563),
            .carryout(n12564),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i13_LC_9_26_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i13_LC_9_26_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i13_LC_9_26_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i13_LC_9_26_5 (
            .in0(N__36073),
            .in1(N__36049),
            .in2(N__36481),
            .in3(N__35923),
            .lcout(encoder0_position_scaled_13),
            .ltout(),
            .carryin(n12564),
            .carryout(n12565),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i14_LC_9_26_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i14_LC_9_26_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i14_LC_9_26_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i14_LC_9_26_6 (
            .in0(N__35920),
            .in1(N__35899),
            .in2(N__36478),
            .in3(N__35788),
            .lcout(encoder0_position_scaled_14),
            .ltout(),
            .carryin(n12565),
            .carryout(n12566),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i15_LC_9_26_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i15_LC_9_26_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i15_LC_9_26_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i15_LC_9_26_7 (
            .in0(N__35785),
            .in1(N__35770),
            .in2(N__36482),
            .in3(N__35656),
            .lcout(encoder0_position_scaled_15),
            .ltout(),
            .carryin(n12566),
            .carryout(n12567),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i16_LC_9_27_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i16_LC_9_27_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i16_LC_9_27_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i16_LC_9_27_0 (
            .in0(N__35653),
            .in1(N__35629),
            .in2(N__36483),
            .in3(N__35530),
            .lcout(encoder0_position_scaled_16),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(n12568),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i17_LC_9_27_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i17_LC_9_27_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i17_LC_9_27_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i17_LC_9_27_1 (
            .in0(N__35527),
            .in1(N__36454),
            .in2(N__35503),
            .in3(N__35422),
            .lcout(encoder0_position_scaled_17),
            .ltout(),
            .carryin(n12568),
            .carryout(n12569),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i18_LC_9_27_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i18_LC_9_27_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i18_LC_9_27_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i18_LC_9_27_2 (
            .in0(N__35419),
            .in1(N__35398),
            .in2(N__36484),
            .in3(N__35320),
            .lcout(encoder0_position_scaled_18),
            .ltout(),
            .carryin(n12569),
            .carryout(n12570),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i19_LC_9_27_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i19_LC_9_27_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i19_LC_9_27_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i19_LC_9_27_3 (
            .in0(N__35317),
            .in1(N__36458),
            .in2(N__35293),
            .in3(N__35200),
            .lcout(encoder0_position_scaled_19),
            .ltout(),
            .carryin(n12570),
            .carryout(n12571),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i20_LC_9_27_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i20_LC_9_27_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i20_LC_9_27_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i20_LC_9_27_4 (
            .in0(N__36766),
            .in1(N__36745),
            .in2(N__36485),
            .in3(N__36673),
            .lcout(encoder0_position_scaled_20),
            .ltout(),
            .carryin(n12571),
            .carryout(n12572),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i21_LC_9_27_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i21_LC_9_27_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i21_LC_9_27_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i21_LC_9_27_5 (
            .in0(N__36670),
            .in1(N__36462),
            .in2(N__36646),
            .in3(N__36577),
            .lcout(encoder0_position_scaled_21),
            .ltout(),
            .carryin(n12572),
            .carryout(n12573),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i22_LC_9_27_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i22_LC_9_27_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i22_LC_9_27_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i22_LC_9_27_6 (
            .in0(N__36574),
            .in1(N__36550),
            .in2(N__36486),
            .in3(N__36490),
            .lcout(encoder0_position_scaled_22),
            .ltout(),
            .carryin(n12573),
            .carryout(n12574),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i23_LC_9_27_7.C_ON=1'b0;
    defparam encoder0_position_scaled_i23_LC_9_27_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i23_LC_9_27_7.LUT_INIT=16'b1100010111001010;
    LogicCell40 encoder0_position_scaled_i23_LC_9_27_7 (
            .in0(N__36970),
            .in1(N__36904),
            .in2(N__36487),
            .in3(N__36316),
            .lcout(encoder0_position_scaled_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i18_1_lut_LC_9_28_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i18_1_lut_LC_9_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i18_1_lut_LC_9_28_0.LUT_INIT=16'b0011001100110011;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i18_1_lut_LC_9_28_0 (
            .in0(_gnd_net_),
            .in1(N__36313),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n8_adj_562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i21_1_lut_LC_9_28_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i21_1_lut_LC_9_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i21_1_lut_LC_9_28_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i21_1_lut_LC_9_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36307),
            .lcout(n5_adj_565),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_9_28_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_9_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_9_28_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i26_3_lut_LC_9_28_2 (
            .in0(_gnd_net_),
            .in1(N__39542),
            .in2(N__36301),
            .in3(N__36271),
            .lcout(n294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i2_LC_9_28_4.C_ON=1'b0;
    defparam commutation_state_i2_LC_9_28_4.SEQ_MODE=4'b1000;
    defparam commutation_state_i2_LC_9_28_4.LUT_INIT=16'b1010001100100010;
    LogicCell40 commutation_state_i2_LC_9_28_4 (
            .in0(N__38150),
            .in1(N__38096),
            .in2(N__38203),
            .in3(N__56133),
            .lcout(commutation_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56061),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_9_28_6.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_9_28_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_9_28_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_2_lut_3_lut_LC_9_28_6 (
            .in0(N__38199),
            .in1(N__38148),
            .in2(_gnd_net_),
            .in3(N__38095),
            .lcout(commutation_state_7__N_261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i24_1_lut_LC_9_28_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i24_1_lut_LC_9_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i24_1_lut_LC_9_28_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i24_1_lut_LC_9_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36991),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_3_lut_LC_9_29_6.C_ON=1'b0;
    defparam i14_3_lut_LC_9_29_6.SEQ_MODE=4'b0000;
    defparam i14_3_lut_LC_9_29_6.LUT_INIT=16'b0111011111101110;
    LogicCell40 i14_3_lut_LC_9_29_6 (
            .in0(N__38192),
            .in1(N__38149),
            .in2(_gnd_net_),
            .in3(N__38097),
            .lcout(n6_adj_592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i0_LC_9_29_7 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i0_LC_9_29_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i0_LC_9_29_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.a_new_i0_LC_9_29_7  (
            .in0(N__36985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.a_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56064),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i16_3_lut_3_lut_LC_9_30_0.C_ON=1'b0;
    defparam LessThan_275_i16_3_lut_3_lut_LC_9_30_0.SEQ_MODE=4'b0000;
    defparam LessThan_275_i16_3_lut_3_lut_LC_9_30_0.LUT_INIT=16'b1101110101000100;
    LogicCell40 LessThan_275_i16_3_lut_3_lut_LC_9_30_0 (
            .in0(N__40177),
            .in1(N__39848),
            .in2(_gnd_net_),
            .in3(N__52771),
            .lcout(n16_adj_614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i10_4_lut_LC_9_30_2 .C_ON=1'b0;
    defparam \PWM.i10_4_lut_LC_9_30_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i10_4_lut_LC_9_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i10_4_lut_LC_9_30_2  (
            .in0(N__40176),
            .in1(N__44005),
            .in2(N__44035),
            .in3(N__40138),
            .lcout(\PWM.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12738_1_lut_LC_9_30_7.C_ON=1'b0;
    defparam i12738_1_lut_LC_9_30_7.SEQ_MODE=4'b0000;
    defparam i12738_1_lut_LC_9_30_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12738_1_lut_LC_9_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36966),
            .lcout(n15210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12064_4_lut_LC_9_31_1.C_ON=1'b0;
    defparam i12064_4_lut_LC_9_31_1.SEQ_MODE=4'b0000;
    defparam i12064_4_lut_LC_9_31_1.LUT_INIT=16'b1110101011111000;
    LogicCell40 i12064_4_lut_LC_9_31_1 (
            .in0(N__36832),
            .in1(N__36856),
            .in2(N__36793),
            .in3(N__36813),
            .lcout(),
            .ltout(n14536_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12065_3_lut_LC_9_31_2.C_ON=1'b0;
    defparam i12065_3_lut_LC_9_31_2.SEQ_MODE=4'b0000;
    defparam i12065_3_lut_LC_9_31_2.LUT_INIT=16'b0000111101010101;
    LogicCell40 i12065_3_lut_LC_9_31_2 (
            .in0(N__36772),
            .in1(_gnd_net_),
            .in2(N__36892),
            .in3(N__36889),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12063_4_lut_LC_9_31_4.C_ON=1'b0;
    defparam i12063_4_lut_LC_9_31_4.SEQ_MODE=4'b0000;
    defparam i12063_4_lut_LC_9_31_4.LUT_INIT=16'b1101010011000100;
    LogicCell40 i12063_4_lut_LC_9_31_4 (
            .in0(N__36855),
            .in1(N__36831),
            .in2(N__36814),
            .in3(N__36789),
            .lcout(n14535),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_62_LC_10_17_0.C_ON=1'b0;
    defparam i1_4_lut_adj_62_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_62_LC_10_17_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_62_LC_10_17_0 (
            .in0(N__37244),
            .in1(N__38549),
            .in2(N__38468),
            .in3(N__37159),
            .lcout(n14300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_10_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_10_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_10_17_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1789_3_lut_LC_10_17_1 (
            .in0(_gnd_net_),
            .in1(N__37153),
            .in2(N__42432),
            .in3(N__37143),
            .lcout(n2725),
            .ltout(n2725_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_51_LC_10_17_2.C_ON=1'b0;
    defparam i1_3_lut_adj_51_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_51_LC_10_17_2.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_51_LC_10_17_2 (
            .in0(N__42131),
            .in1(_gnd_net_),
            .in2(N__37129),
            .in3(N__44189),
            .lcout(),
            .ltout(n14040_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_53_LC_10_17_3.C_ON=1'b0;
    defparam i1_4_lut_adj_53_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_53_LC_10_17_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_53_LC_10_17_3 (
            .in0(N__40365),
            .in1(N__40341),
            .in2(N__37126),
            .in3(N__37252),
            .lcout(n14048),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_10_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_10_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_10_17_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1792_3_lut_LC_10_17_4 (
            .in0(_gnd_net_),
            .in1(N__37122),
            .in2(N__37102),
            .in3(N__42404),
            .lcout(n2728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_10_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_10_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_10_17_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1793_3_lut_LC_10_17_5 (
            .in0(_gnd_net_),
            .in1(N__37086),
            .in2(N__42431),
            .in3(N__37072),
            .lcout(n2729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_10_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_10_17_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1791_3_lut_LC_10_17_6 (
            .in0(_gnd_net_),
            .in1(N__37063),
            .in2(N__37053),
            .in3(N__42405),
            .lcout(n2727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_10_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_10_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_10_17_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1782_3_lut_LC_10_17_7 (
            .in0(N__42412),
            .in1(_gnd_net_),
            .in2(N__37027),
            .in3(N__37003),
            .lcout(n2718),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12350_3_lut_LC_10_18_0.C_ON=1'b0;
    defparam i12350_3_lut_LC_10_18_0.SEQ_MODE=4'b0000;
    defparam i12350_3_lut_LC_10_18_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 i12350_3_lut_LC_10_18_0 (
            .in0(N__37440),
            .in1(_gnd_net_),
            .in2(N__37414),
            .in3(N__42395),
            .lcout(n2726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_10_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_10_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_10_18_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1716_3_lut_LC_10_18_1 (
            .in0(N__37405),
            .in1(_gnd_net_),
            .in2(N__37375),
            .in3(N__38934),
            .lcout(n2620),
            .ltout(n2620_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_10_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_10_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_10_18_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1783_3_lut_LC_10_18_2 (
            .in0(_gnd_net_),
            .in1(N__37342),
            .in2(N__37333),
            .in3(N__42396),
            .lcout(n2719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12970_4_lut_LC_10_18_3.C_ON=1'b0;
    defparam i12970_4_lut_LC_10_18_3.SEQ_MODE=4'b0000;
    defparam i12970_4_lut_LC_10_18_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12970_4_lut_LC_10_18_3 (
            .in0(N__37326),
            .in1(N__38504),
            .in2(N__37306),
            .in3(N__42473),
            .lcout(n2643),
            .ltout(n2643_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_10_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_10_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_10_18_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1784_3_lut_LC_10_18_4 (
            .in0(N__37296),
            .in1(_gnd_net_),
            .in2(N__37276),
            .in3(N__37273),
            .lcout(n2720),
            .ltout(n2720_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_50_LC_10_18_5.C_ON=1'b0;
    defparam i1_4_lut_adj_50_LC_10_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_50_LC_10_18_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_50_LC_10_18_5 (
            .in0(N__41666),
            .in1(N__42173),
            .in2(N__37258),
            .in3(N__44486),
            .lcout(),
            .ltout(n14038_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_52_LC_10_18_6.C_ON=1'b0;
    defparam i1_4_lut_adj_52_LC_10_18_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_52_LC_10_18_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_52_LC_10_18_6 (
            .in0(N__40254),
            .in1(N__41879),
            .in2(N__37255),
            .in3(N__41951),
            .lcout(n14042),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_10_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_10_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_10_19_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1777_3_lut_LC_10_19_0 (
            .in0(_gnd_net_),
            .in1(N__37246),
            .in2(N__42442),
            .in3(N__37213),
            .lcout(n2713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_10_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_10_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_10_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1781_3_lut_LC_10_19_1 (
            .in0(_gnd_net_),
            .in1(N__37201),
            .in2(N__37192),
            .in3(N__42422),
            .lcout(n2717),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_10_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_10_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_10_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_10_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37780),
            .lcout(n27_adj_651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_19_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_19_4 (
            .in0(N__39564),
            .in1(N__37735),
            .in2(_gnd_net_),
            .in3(N__37720),
            .lcout(n310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_10_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_10_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_10_19_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i15_3_lut_LC_10_19_5 (
            .in0(N__37654),
            .in1(N__39562),
            .in2(_gnd_net_),
            .in3(N__37636),
            .lcout(n305),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_10_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_10_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_10_19_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i11_3_lut_LC_10_19_6 (
            .in0(N__39563),
            .in1(N__37570),
            .in2(_gnd_net_),
            .in3(N__37555),
            .lcout(n309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_10_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_10_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_10_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1779_3_lut_LC_10_19_7 (
            .in0(_gnd_net_),
            .in1(N__37482),
            .in2(N__37456),
            .in3(N__42423),
            .lcout(n2715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_166_LC_10_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_166_LC_10_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_166_LC_10_20_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_166_LC_10_20_0 (
            .in0(N__51498),
            .in1(N__50855),
            .in2(N__51406),
            .in3(N__51548),
            .lcout(),
            .ltout(n13884_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_167_LC_10_20_1.C_ON=1'b0;
    defparam i1_4_lut_adj_167_LC_10_20_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_167_LC_10_20_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_167_LC_10_20_1 (
            .in0(N__51750),
            .in1(N__37813),
            .in2(N__37444),
            .in3(N__37807),
            .lcout(n13894),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_10_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_10_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_10_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2055_3_lut_LC_10_20_2 (
            .in0(_gnd_net_),
            .in1(N__45422),
            .in2(N__45403),
            .in3(N__49069),
            .lcout(n3119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_10_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_10_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_10_20_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2053_3_lut_LC_10_20_3 (
            .in0(_gnd_net_),
            .in1(N__45338),
            .in2(N__49084),
            .in3(N__45322),
            .lcout(n3117),
            .ltout(n3117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_165_LC_10_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_165_LC_10_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_165_LC_10_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_165_LC_10_20_4 (
            .in0(N__51842),
            .in1(N__50799),
            .in2(N__37816),
            .in3(N__51273),
            .lcout(n13888),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_164_LC_10_20_5.C_ON=1'b0;
    defparam i1_4_lut_adj_164_LC_10_20_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_164_LC_10_20_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_164_LC_10_20_5 (
            .in0(N__51310),
            .in1(N__51434),
            .in2(N__51348),
            .in3(N__51212),
            .lcout(n13886),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_10_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_10_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_10_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_2_lut_LC_10_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47430),
            .in3(N__37801),
            .lcout(n3001),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(n12437),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_10_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_10_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_10_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_3_lut_LC_10_21_1 (
            .in0(_gnd_net_),
            .in1(N__54699),
            .in2(N__47407),
            .in3(N__37798),
            .lcout(n3000),
            .ltout(),
            .carryin(n12437),
            .carryout(n12438),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_10_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_10_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_10_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_4_lut_LC_10_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47464),
            .in3(N__37795),
            .lcout(n2999),
            .ltout(),
            .carryin(n12438),
            .carryout(n12439),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_10_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_10_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_10_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_5_lut_LC_10_21_3 (
            .in0(_gnd_net_),
            .in1(N__54700),
            .in2(N__47350),
            .in3(N__37792),
            .lcout(n2998),
            .ltout(),
            .carryin(n12439),
            .carryout(n12440),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_10_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_10_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_10_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_6_lut_LC_10_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47377),
            .in3(N__37789),
            .lcout(n2997),
            .ltout(),
            .carryin(n12440),
            .carryout(n12441),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_10_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_10_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_10_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_7_lut_LC_10_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47314),
            .in3(N__37786),
            .lcout(n2996),
            .ltout(),
            .carryin(n12441),
            .carryout(n12442),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_10_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_10_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_10_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_8_lut_LC_10_21_6 (
            .in0(_gnd_net_),
            .in1(N__54702),
            .in2(N__44572),
            .in3(N__37783),
            .lcout(n2995),
            .ltout(),
            .carryin(n12442),
            .carryout(n12443),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_10_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_10_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_10_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_9_lut_LC_10_21_7 (
            .in0(_gnd_net_),
            .in1(N__54701),
            .in2(N__44629),
            .in3(N__37843),
            .lcout(n2994),
            .ltout(),
            .carryin(n12443),
            .carryout(n12444),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_10_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_10_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_10_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_10_lut_LC_10_22_0 (
            .in0(_gnd_net_),
            .in1(N__44697),
            .in2(N__54321),
            .in3(N__37840),
            .lcout(n2993),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(n12445),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_10_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_10_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_10_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_11_lut_LC_10_22_1 (
            .in0(_gnd_net_),
            .in1(N__53858),
            .in2(N__44950),
            .in3(N__37837),
            .lcout(n2992),
            .ltout(),
            .carryin(n12445),
            .carryout(n12446),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_10_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_10_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_10_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_12_lut_LC_10_22_2 (
            .in0(_gnd_net_),
            .in1(N__53860),
            .in2(N__44467),
            .in3(N__37834),
            .lcout(n2991),
            .ltout(),
            .carryin(n12446),
            .carryout(n12447),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_10_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_10_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_10_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_13_lut_LC_10_22_3 (
            .in0(_gnd_net_),
            .in1(N__53859),
            .in2(N__44304),
            .in3(N__37831),
            .lcout(n2990),
            .ltout(),
            .carryin(n12447),
            .carryout(n12448),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_10_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_10_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_10_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_14_lut_LC_10_22_4 (
            .in0(_gnd_net_),
            .in1(N__53861),
            .in2(N__44545),
            .in3(N__37828),
            .lcout(n2989),
            .ltout(),
            .carryin(n12448),
            .carryout(n12449),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_10_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_10_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_10_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_15_lut_LC_10_22_5 (
            .in0(_gnd_net_),
            .in1(N__42117),
            .in2(N__54322),
            .in3(N__37825),
            .lcout(n2988),
            .ltout(),
            .carryin(n12449),
            .carryout(n12450),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_10_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_10_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_10_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_16_lut_LC_10_22_6 (
            .in0(_gnd_net_),
            .in1(N__53865),
            .in2(N__44667),
            .in3(N__37822),
            .lcout(n2987),
            .ltout(),
            .carryin(n12450),
            .carryout(n12451),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_10_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_10_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_10_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_17_lut_LC_10_22_7 (
            .in0(_gnd_net_),
            .in1(N__44601),
            .in2(N__54323),
            .in3(N__37819),
            .lcout(n2986),
            .ltout(),
            .carryin(n12451),
            .carryout(n12452),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_10_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_10_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_10_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_18_lut_LC_10_23_0 (
            .in0(_gnd_net_),
            .in1(N__42064),
            .in2(N__55185),
            .in3(N__37870),
            .lcout(n2985),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(n12453),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_10_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_10_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_10_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_19_lut_LC_10_23_1 (
            .in0(_gnd_net_),
            .in1(N__55034),
            .in2(N__42091),
            .in3(N__37867),
            .lcout(n2984),
            .ltout(),
            .carryin(n12453),
            .carryout(n12454),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_10_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_10_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_10_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_20_lut_LC_10_23_2 (
            .in0(_gnd_net_),
            .in1(N__42531),
            .in2(N__55186),
            .in3(N__37864),
            .lcout(n2983),
            .ltout(),
            .carryin(n12454),
            .carryout(n12455),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_10_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_10_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_10_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_21_lut_LC_10_23_3 (
            .in0(_gnd_net_),
            .in1(N__42559),
            .in2(N__54603),
            .in3(N__37861),
            .lcout(n2982),
            .ltout(),
            .carryin(n12455),
            .carryout(n12456),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_10_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_10_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_10_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_22_lut_LC_10_23_4 (
            .in0(_gnd_net_),
            .in1(N__44919),
            .in2(N__55187),
            .in3(N__37858),
            .lcout(n2981),
            .ltout(),
            .carryin(n12456),
            .carryout(n12457),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_10_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_10_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_10_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_23_lut_LC_10_23_5 (
            .in0(_gnd_net_),
            .in1(N__42606),
            .in2(N__54604),
            .in3(N__37855),
            .lcout(n2980),
            .ltout(),
            .carryin(n12457),
            .carryout(n12458),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_10_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_10_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_10_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_24_lut_LC_10_23_6 (
            .in0(_gnd_net_),
            .in1(N__54115),
            .in2(N__40522),
            .in3(N__37852),
            .lcout(n2979),
            .ltout(),
            .carryin(n12458),
            .carryout(n12459),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_10_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_10_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_10_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_25_lut_LC_10_23_7 (
            .in0(_gnd_net_),
            .in1(N__40545),
            .in2(N__54605),
            .in3(N__37849),
            .lcout(n2978),
            .ltout(),
            .carryin(n12459),
            .carryout(n12460),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_10_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_10_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_10_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_26_lut_LC_10_24_0 (
            .in0(_gnd_net_),
            .in1(N__47110),
            .in2(N__55188),
            .in3(N__37846),
            .lcout(n2977),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(n12461),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_10_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_10_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_10_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_27_lut_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(N__42261),
            .in2(N__54976),
            .in3(N__37885),
            .lcout(n2976),
            .ltout(),
            .carryin(n12461),
            .carryout(n12462),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_10_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_10_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_10_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_28_lut_LC_10_24_2 (
            .in0(_gnd_net_),
            .in1(N__40474),
            .in2(N__55189),
            .in3(N__37882),
            .lcout(n2975),
            .ltout(),
            .carryin(n12462),
            .carryout(n12463),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_10_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_10_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_10_24_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1972_29_lut_LC_10_24_3 (
            .in0(N__54593),
            .in1(N__39756),
            .in2(N__48766),
            .in3(N__37879),
            .lcout(n3006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_10_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_10_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_10_24_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2111_3_lut_LC_10_24_4 (
            .in0(_gnd_net_),
            .in1(N__52063),
            .in2(N__50071),
            .in3(N__52092),
            .lcout(n3207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_10_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_10_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_10_24_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2112_3_lut_LC_10_24_5 (
            .in0(_gnd_net_),
            .in1(N__52133),
            .in2(N__52114),
            .in3(N__50025),
            .lcout(n3208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_10_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_10_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_10_24_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2109_3_lut_LC_10_24_6 (
            .in0(_gnd_net_),
            .in1(N__51970),
            .in2(N__50072),
            .in3(N__51996),
            .lcout(n3205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_10_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_10_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_10_24_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2114_3_lut_LC_10_24_7 (
            .in0(N__52224),
            .in1(_gnd_net_),
            .in2(N__52189),
            .in3(N__50024),
            .lcout(n3210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12725_1_lut_LC_10_25_0.C_ON=1'b0;
    defparam i12725_1_lut_LC_10_25_0.SEQ_MODE=4'b0000;
    defparam i12725_1_lut_LC_10_25_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12725_1_lut_LC_10_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37923),
            .lcout(n15197),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_LC_10_25_1.C_ON=1'b0;
    defparam i16_4_lut_LC_10_25_1.SEQ_MODE=4'b0000;
    defparam i16_4_lut_LC_10_25_1.LUT_INIT=16'b1100101000001010;
    LogicCell40 i16_4_lut_LC_10_25_1 (
            .in0(N__43078),
            .in1(N__42687),
            .in2(N__49606),
            .in3(N__43104),
            .lcout(n5_adj_713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9879_4_lut_LC_10_25_2.C_ON=1'b0;
    defparam i9879_4_lut_LC_10_25_2.SEQ_MODE=4'b0000;
    defparam i9879_4_lut_LC_10_25_2.LUT_INIT=16'b1110111011111010;
    LogicCell40 i9879_4_lut_LC_10_25_2 (
            .in0(N__42849),
            .in1(N__42822),
            .in2(N__42787),
            .in3(N__49569),
            .lcout(),
            .ltout(n11593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9941_4_lut_LC_10_25_3.C_ON=1'b0;
    defparam i9941_4_lut_LC_10_25_3.SEQ_MODE=4'b0000;
    defparam i9941_4_lut_LC_10_25_3.LUT_INIT=16'b1110000001000000;
    LogicCell40 i9941_4_lut_LC_10_25_3 (
            .in0(N__49573),
            .in1(N__42745),
            .in2(N__37930),
            .in3(N__42765),
            .lcout(n11656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12686_1_lut_LC_10_25_4.C_ON=1'b0;
    defparam i12686_1_lut_LC_10_25_4.SEQ_MODE=4'b0000;
    defparam i12686_1_lut_LC_10_25_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12686_1_lut_LC_10_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50023),
            .lcout(n15158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12691_1_lut_LC_10_25_5.C_ON=1'b0;
    defparam i12691_1_lut_LC_10_25_5.SEQ_MODE=4'b0000;
    defparam i12691_1_lut_LC_10_25_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12691_1_lut_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49607),
            .in3(_gnd_net_),
            .lcout(n15163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_10_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_10_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2177_3_lut_LC_10_25_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i2177_3_lut_LC_10_25_6 (
            .in0(N__43642),
            .in1(N__43661),
            .in2(_gnd_net_),
            .in3(N__49577),
            .lcout(),
            .ltout(n59_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12728_4_lut_LC_10_25_7.C_ON=1'b0;
    defparam i12728_4_lut_LC_10_25_7.SEQ_MODE=4'b0000;
    defparam i12728_4_lut_LC_10_25_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12728_4_lut_LC_10_25_7 (
            .in0(N__39715),
            .in1(N__43570),
            .in2(N__37927),
            .in3(N__39802),
            .lcout(n11838),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i1_1_lut_LC_10_26_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i1_1_lut_LC_10_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i1_1_lut_LC_10_26_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i1_1_lut_LC_10_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37909),
            .lcout(n25_adj_545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i16_1_lut_LC_10_26_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i16_1_lut_LC_10_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i16_1_lut_LC_10_26_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i16_1_lut_LC_10_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37903),
            .lcout(n10_adj_560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i13_1_lut_LC_10_26_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i13_1_lut_LC_10_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i13_1_lut_LC_10_26_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i13_1_lut_LC_10_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37897),
            .lcout(n13_adj_557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i3_1_lut_LC_10_26_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i3_1_lut_LC_10_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i3_1_lut_LC_10_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i3_1_lut_LC_10_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37891),
            .lcout(n23_adj_547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i5_1_lut_LC_10_26_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i5_1_lut_LC_10_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i5_1_lut_LC_10_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i5_1_lut_LC_10_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38017),
            .lcout(n21_adj_549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12457_2_lut_LC_10_27_0.C_ON=1'b0;
    defparam i12457_2_lut_LC_10_27_0.SEQ_MODE=4'b0000;
    defparam i12457_2_lut_LC_10_27_0.LUT_INIT=16'b1111111100110011;
    LogicCell40 i12457_2_lut_LC_10_27_0 (
            .in0(_gnd_net_),
            .in1(N__55495),
            .in2(_gnd_net_),
            .in3(N__55469),
            .lcout(),
            .ltout(dti_N_333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_10_27_1.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_10_27_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_10_27_1.LUT_INIT=16'b1111111101101111;
    LogicCell40 i1_2_lut_4_lut_LC_10_27_1 (
            .in0(N__41066),
            .in1(N__56251),
            .in2(N__38011),
            .in3(N__41124),
            .lcout(n4828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i23_1_lut_LC_10_27_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i23_1_lut_LC_10_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i23_1_lut_LC_10_27_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i23_1_lut_LC_10_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38008),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_10_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_10_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_10_27_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i8_3_lut_LC_10_27_3 (
            .in0(N__38002),
            .in1(N__39558),
            .in2(_gnd_net_),
            .in3(N__37990),
            .lcout(n312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i20_1_lut_LC_10_27_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i20_1_lut_LC_10_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i20_1_lut_LC_10_27_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i20_1_lut_LC_10_27_4 (
            .in0(N__37960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n6_adj_564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i22_1_lut_LC_10_27_5.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i22_1_lut_LC_10_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i22_1_lut_LC_10_27_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i22_1_lut_LC_10_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37954),
            .lcout(n4_adj_566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i14_1_lut_LC_10_27_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i14_1_lut_LC_10_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i14_1_lut_LC_10_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i14_1_lut_LC_10_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37948),
            .lcout(n12_adj_558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_154_LC_10_28_3.C_ON=1'b0;
    defparam dti_154_LC_10_28_3.SEQ_MODE=4'b1000;
    defparam dti_154_LC_10_28_3.LUT_INIT=16'b1111111100110011;
    LogicCell40 dti_154_LC_10_28_3 (
            .in0(_gnd_net_),
            .in1(N__55506),
            .in2(_gnd_net_),
            .in3(N__55470),
            .lcout(dti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(N__37942),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_28_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38304),
            .lcout(n20_adj_644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38263),
            .lcout(n5_adj_629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i10_1_lut_LC_10_28_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i10_1_lut_LC_10_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i10_1_lut_LC_10_28_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i10_1_lut_LC_10_28_6 (
            .in0(N__38221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n16_adj_554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i11_1_lut_LC_10_28_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i11_1_lut_LC_10_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i11_1_lut_LC_10_28_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i11_1_lut_LC_10_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38212),
            .lcout(n15_adj_555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i0_LC_10_29_0.C_ON=1'b0;
    defparam commutation_state_i0_LC_10_29_0.SEQ_MODE=4'b1001;
    defparam commutation_state_i0_LC_10_29_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 commutation_state_i0_LC_10_29_0 (
            .in0(N__38198),
            .in1(N__38154),
            .in2(_gnd_net_),
            .in3(N__38098),
            .lcout(commutation_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56065),
            .ce(N__38041),
            .sr(N__38029));
    defparam LessThan_275_i13_2_lut_LC_10_29_2.C_ON=1'b0;
    defparam LessThan_275_i13_2_lut_LC_10_29_2.SEQ_MODE=4'b0000;
    defparam LessThan_275_i13_2_lut_LC_10_29_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i13_2_lut_LC_10_29_2 (
            .in0(_gnd_net_),
            .in1(N__41272),
            .in2(_gnd_net_),
            .in3(N__41164),
            .lcout(n13_adj_612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i23_2_lut_LC_10_29_3.C_ON=1'b0;
    defparam LessThan_275_i23_2_lut_LC_10_29_3.SEQ_MODE=4'b0000;
    defparam LessThan_275_i23_2_lut_LC_10_29_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i23_2_lut_LC_10_29_3 (
            .in0(_gnd_net_),
            .in1(N__41007),
            .in2(_gnd_net_),
            .in3(N__39947),
            .lcout(n23_adj_618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i11_4_lut_LC_10_30_0 .C_ON=1'b0;
    defparam \PWM.i11_4_lut_LC_10_30_0 .SEQ_MODE=4'b0000;
    defparam \PWM.i11_4_lut_LC_10_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i11_4_lut_LC_10_30_0  (
            .in0(N__40005),
            .in1(N__40974),
            .in2(N__39952),
            .in3(N__46766),
            .lcout(\PWM.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i41_2_lut_LC_10_30_1.C_ON=1'b0;
    defparam LessThan_275_i41_2_lut_LC_10_30_1.SEQ_MODE=4'b0000;
    defparam LessThan_275_i41_2_lut_LC_10_30_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i41_2_lut_LC_10_30_1 (
            .in0(_gnd_net_),
            .in1(N__41202),
            .in2(_gnd_net_),
            .in3(N__40004),
            .lcout(n41),
            .ltout(n41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12407_3_lut_LC_10_30_2.C_ON=1'b0;
    defparam i12407_3_lut_LC_10_30_2.SEQ_MODE=4'b0000;
    defparam i12407_3_lut_LC_10_30_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12407_3_lut_LC_10_30_2 (
            .in0(N__41203),
            .in1(_gnd_net_),
            .in2(N__38329),
            .in3(N__41362),
            .lcout(n40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12243_4_lut_LC_10_30_4.C_ON=1'b0;
    defparam i12243_4_lut_LC_10_30_4.SEQ_MODE=4'b0000;
    defparam i12243_4_lut_LC_10_30_4.LUT_INIT=16'b1111000011110001;
    LogicCell40 i12243_4_lut_LC_10_30_4 (
            .in0(N__38326),
            .in1(N__41386),
            .in2(N__38362),
            .in3(N__41743),
            .lcout(),
            .ltout(n14715_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12394_4_lut_LC_10_30_5.C_ON=1'b0;
    defparam i12394_4_lut_LC_10_30_5.SEQ_MODE=4'b0000;
    defparam i12394_4_lut_LC_10_30_5.LUT_INIT=16'b1100110111001000;
    LogicCell40 i12394_4_lut_LC_10_30_5 (
            .in0(N__38395),
            .in1(N__38371),
            .in2(N__38320),
            .in3(N__38317),
            .lcout(),
            .ltout(n14866_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.pwm_out_12_LC_10_30_6 .C_ON=1'b0;
    defparam \PWM.pwm_out_12_LC_10_30_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_out_12_LC_10_30_6 .LUT_INIT=16'b1100000011111100;
    LogicCell40 \PWM.pwm_out_12_LC_10_30_6  (
            .in0(_gnd_net_),
            .in1(N__43855),
            .in2(N__38311),
            .in3(N__44060),
            .lcout(pwm_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56069),
            .ce(),
            .sr(N__41251));
    defparam LessThan_275_i8_3_lut_3_lut_LC_10_31_0.C_ON=1'b0;
    defparam LessThan_275_i8_3_lut_3_lut_LC_10_31_0.SEQ_MODE=4'b0000;
    defparam LessThan_275_i8_3_lut_3_lut_LC_10_31_0.LUT_INIT=16'b1011101100100010;
    LogicCell40 LessThan_275_i8_3_lut_3_lut_LC_10_31_0 (
            .in0(N__40993),
            .in1(N__41531),
            .in2(_gnd_net_),
            .in3(N__40804),
            .lcout(n8_adj_607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i17_2_lut_LC_10_31_2.C_ON=1'b0;
    defparam LessThan_275_i17_2_lut_LC_10_31_2.SEQ_MODE=4'b0000;
    defparam LessThan_275_i17_2_lut_LC_10_31_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i17_2_lut_LC_10_31_2 (
            .in0(_gnd_net_),
            .in1(N__40992),
            .in2(_gnd_net_),
            .in3(N__41530),
            .lcout(n17_adj_615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_10_31_3.C_ON=1'b0;
    defparam i5_4_lut_LC_10_31_3.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_10_31_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_10_31_3 (
            .in0(N__40044),
            .in1(N__40107),
            .in2(N__40063),
            .in3(N__40227),
            .lcout(),
            .ltout(n12_adj_598_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_10_31_4.C_ON=1'b0;
    defparam i6_4_lut_LC_10_31_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_10_31_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_10_31_4 (
            .in0(N__40077),
            .in1(N__40212),
            .in2(N__38308),
            .in3(N__40092),
            .lcout(n4823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i45_2_lut_LC_10_31_5.C_ON=1'b0;
    defparam LessThan_275_i45_2_lut_LC_10_31_5.SEQ_MODE=4'b0000;
    defparam LessThan_275_i45_2_lut_LC_10_31_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i45_2_lut_LC_10_31_5 (
            .in0(_gnd_net_),
            .in1(N__43950),
            .in2(_gnd_net_),
            .in3(N__40130),
            .lcout(n45),
            .ltout(n45_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i24_3_lut_LC_10_31_6.C_ON=1'b0;
    defparam LessThan_275_i24_3_lut_LC_10_31_6.SEQ_MODE=4'b0000;
    defparam LessThan_275_i24_3_lut_LC_10_31_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 LessThan_275_i24_3_lut_LC_10_31_6 (
            .in0(N__43951),
            .in1(_gnd_net_),
            .in2(N__38422),
            .in3(N__38419),
            .lcout(n24_adj_619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i43_2_lut_LC_10_31_7.C_ON=1'b0;
    defparam LessThan_275_i43_2_lut_LC_10_31_7.SEQ_MODE=4'b0000;
    defparam LessThan_275_i43_2_lut_LC_10_31_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_275_i43_2_lut_LC_10_31_7 (
            .in0(N__39849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40175),
            .lcout(n43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12371_3_lut_LC_10_32_1.C_ON=1'b0;
    defparam i12371_3_lut_LC_10_32_1.SEQ_MODE=4'b0000;
    defparam i12371_3_lut_LC_10_32_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12371_3_lut_LC_10_32_1 (
            .in0(N__41828),
            .in1(N__41011),
            .in2(_gnd_net_),
            .in3(N__40948),
            .lcout(),
            .ltout(n14843_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12307_3_lut_LC_10_32_2.C_ON=1'b0;
    defparam i12307_3_lut_LC_10_32_2.SEQ_MODE=4'b0000;
    defparam i12307_3_lut_LC_10_32_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12307_3_lut_LC_10_32_2 (
            .in0(_gnd_net_),
            .in1(N__41731),
            .in2(N__38413),
            .in3(N__41691),
            .lcout(n14779),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12239_2_lut_4_lut_LC_10_32_3.C_ON=1'b0;
    defparam i12239_2_lut_4_lut_LC_10_32_3.SEQ_MODE=4'b0000;
    defparam i12239_2_lut_4_lut_LC_10_32_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i12239_2_lut_4_lut_LC_10_32_3 (
            .in0(N__39850),
            .in1(N__52770),
            .in2(N__41350),
            .in3(N__40168),
            .lcout(),
            .ltout(n14711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12354_4_lut_LC_10_32_4.C_ON=1'b0;
    defparam i12354_4_lut_LC_10_32_4.SEQ_MODE=4'b0000;
    defparam i12354_4_lut_LC_10_32_4.LUT_INIT=16'b1010101110101000;
    LogicCell40 i12354_4_lut_LC_10_32_4 (
            .in0(N__38410),
            .in1(N__38393),
            .in2(N__38404),
            .in3(N__38401),
            .lcout(),
            .ltout(n14826_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12392_4_lut_LC_10_32_5.C_ON=1'b0;
    defparam i12392_4_lut_LC_10_32_5.SEQ_MODE=4'b0000;
    defparam i12392_4_lut_LC_10_32_5.LUT_INIT=16'b1111000111100000;
    LogicCell40 i12392_4_lut_LC_10_32_5 (
            .in0(N__38394),
            .in1(N__38347),
            .in2(N__38380),
            .in3(N__38377),
            .lcout(n14864),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12241_4_lut_LC_10_32_7.C_ON=1'b0;
    defparam i12241_4_lut_LC_10_32_7.SEQ_MODE=4'b0000;
    defparam i12241_4_lut_LC_10_32_7.LUT_INIT=16'b1111111100000001;
    LogicCell40 i12241_4_lut_LC_10_32_7 (
            .in0(N__41692),
            .in1(N__41752),
            .in2(N__41833),
            .in3(N__38358),
            .lcout(n14713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_11_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_11_17_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1796_3_lut_LC_11_17_0 (
            .in0(_gnd_net_),
            .in1(N__38341),
            .in2(N__42427),
            .in3(N__38737),
            .lcout(n2732),
            .ltout(n2732_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9951_3_lut_LC_11_17_1.C_ON=1'b0;
    defparam i9951_3_lut_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam i9951_3_lut_LC_11_17_1.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9951_3_lut_LC_11_17_1 (
            .in0(_gnd_net_),
            .in1(N__47678),
            .in2(N__38662),
            .in3(N__44381),
            .lcout(),
            .ltout(n11666_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_54_LC_11_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_54_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_54_LC_11_17_2.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_54_LC_11_17_2 (
            .in0(N__41852),
            .in1(N__41981),
            .in2(N__38659),
            .in3(N__44423),
            .lcout(n13403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12346_3_lut_LC_11_17_3.C_ON=1'b0;
    defparam i12346_3_lut_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam i12346_3_lut_LC_11_17_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12346_3_lut_LC_11_17_3 (
            .in0(_gnd_net_),
            .in1(N__38656),
            .in2(N__38644),
            .in3(N__42382),
            .lcout(n2723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_11_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_11_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_11_17_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1780_3_lut_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(N__38611),
            .in2(N__42428),
            .in3(N__38581),
            .lcout(n2716),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_11_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_11_17_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1797_3_lut_LC_11_17_5 (
            .in0(N__38569),
            .in1(N__38776),
            .in2(_gnd_net_),
            .in3(N__42383),
            .lcout(n2733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_11_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_11_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_11_17_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1776_3_lut_LC_11_17_7 (
            .in0(_gnd_net_),
            .in1(N__38550),
            .in2(N__38527),
            .in3(N__42390),
            .lcout(n2712),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_11_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_11_18_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1774_3_lut_LC_11_18_0 (
            .in0(N__38511),
            .in1(N__38482),
            .in2(_gnd_net_),
            .in3(N__42403),
            .lcout(n2710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_11_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_11_18_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1848_3_lut_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(N__40340),
            .in2(N__40318),
            .in3(N__47628),
            .lcout(n2816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_11_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_11_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_11_18_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1778_3_lut_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(N__38469),
            .in2(N__38437),
            .in3(N__42402),
            .lcout(n2714),
            .ltout(n2714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_11_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_11_18_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1845_3_lut_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(N__40300),
            .in2(N__39271),
            .in3(N__47627),
            .lcout(n2813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12345_3_lut_LC_11_18_4.C_ON=1'b0;
    defparam i12345_3_lut_LC_11_18_4.SEQ_MODE=4'b0000;
    defparam i12345_3_lut_LC_11_18_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12345_3_lut_LC_11_18_4 (
            .in0(_gnd_net_),
            .in1(N__39264),
            .in2(N__39238),
            .in3(N__42397),
            .lcout(n2722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_11_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_11_18_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1794_3_lut_LC_11_18_5 (
            .in0(_gnd_net_),
            .in1(N__39223),
            .in2(N__42430),
            .in3(N__38704),
            .lcout(n2730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_11_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_11_18_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1795_3_lut_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(N__38790),
            .in2(N__39211),
            .in3(N__42398),
            .lcout(n2731),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_11_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_11_19_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1508_3_lut_LC_11_19_0 (
            .in0(_gnd_net_),
            .in1(N__39195),
            .in2(N__39166),
            .in3(N__39149),
            .lcout(n2316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_11_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_11_19_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1728_3_lut_LC_11_19_1 (
            .in0(_gnd_net_),
            .in1(N__38989),
            .in2(N__38962),
            .in3(N__38931),
            .lcout(n2632),
            .ltout(n2632_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10045_4_lut_LC_11_19_2.C_ON=1'b0;
    defparam i10045_4_lut_LC_11_19_2.SEQ_MODE=4'b0000;
    defparam i10045_4_lut_LC_11_19_2.LUT_INIT=16'b1111111111100000;
    LogicCell40 i10045_4_lut_LC_11_19_2 (
            .in0(N__38774),
            .in1(N__38729),
            .in2(N__38707),
            .in3(N__38696),
            .lcout(n11760),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_11_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_11_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_11_19_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1849_3_lut_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__40378),
            .in2(N__40354),
            .in3(N__47629),
            .lcout(n2817),
            .ltout(n2817_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_11_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_11_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_11_19_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1916_3_lut_LC_11_19_5 (
            .in0(_gnd_net_),
            .in1(N__48568),
            .in2(N__39601),
            .in3(N__49366),
            .lcout(n2916),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_11_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_11_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_11_20_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2000_3_lut_LC_11_20_0 (
            .in0(N__47406),
            .in1(N__39598),
            .in2(N__42997),
            .in3(_gnd_net_),
            .lcout(n3032),
            .ltout(n3032_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9945_3_lut_LC_11_20_1.C_ON=1'b0;
    defparam i9945_3_lut_LC_11_20_1.SEQ_MODE=4'b0000;
    defparam i9945_3_lut_LC_11_20_1.LUT_INIT=16'b1111000010100000;
    LogicCell40 i9945_3_lut_LC_11_20_1 (
            .in0(N__44888),
            .in1(_gnd_net_),
            .in2(N__39592),
            .in3(N__44819),
            .lcout(),
            .ltout(n11660_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_31_LC_11_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_31_LC_11_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_31_LC_11_20_2.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_31_LC_11_20_2 (
            .in0(N__45221),
            .in1(N__44732),
            .in2(N__39589),
            .in3(N__45180),
            .lcout(n13466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_11_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_11_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_11_20_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1986_3_lut_LC_11_20_3 (
            .in0(_gnd_net_),
            .in1(N__44602),
            .in2(N__39586),
            .in3(N__42960),
            .lcout(n3018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_11_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_11_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_11_20_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1997_3_lut_LC_11_20_4 (
            .in0(_gnd_net_),
            .in1(N__47376),
            .in2(N__42996),
            .in3(N__39574),
            .lcout(n3029),
            .ltout(n3029_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_11_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_11_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_11_20_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2064_3_lut_LC_11_20_5 (
            .in0(_gnd_net_),
            .in1(N__45169),
            .in2(N__39568),
            .in3(N__49075),
            .lcout(n3128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_11_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_11_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_11_20_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i5_3_lut_LC_11_20_6 (
            .in0(N__39565),
            .in1(N__39325),
            .in2(_gnd_net_),
            .in3(N__39313),
            .lcout(n315),
            .ltout(n315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_11_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_11_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_11_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2001_3_lut_LC_11_20_7 (
            .in0(_gnd_net_),
            .in1(N__39280),
            .in2(N__39274),
            .in3(N__42953),
            .lcout(n3033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_11_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_11_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_11_21_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1998_3_lut_LC_11_21_0 (
            .in0(_gnd_net_),
            .in1(N__39652),
            .in2(N__42998),
            .in3(N__47346),
            .lcout(n3030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_11_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_11_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_11_21_1.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2063_3_lut_LC_11_21_1 (
            .in0(N__45150),
            .in1(N__45130),
            .in2(N__49043),
            .in3(_gnd_net_),
            .lcout(n3127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_11_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_11_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_11_21_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2051_3_lut_LC_11_21_2 (
            .in0(_gnd_net_),
            .in1(N__45247),
            .in2(N__45273),
            .in3(N__49000),
            .lcout(n3115),
            .ltout(n3115_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_168_LC_11_21_3.C_ON=1'b0;
    defparam i1_3_lut_adj_168_LC_11_21_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_168_LC_11_21_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_168_LC_11_21_3 (
            .in0(_gnd_net_),
            .in1(N__51670),
            .in2(N__39646),
            .in3(N__39643),
            .lcout(n13898),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_11_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_11_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_11_21_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1988_3_lut_LC_11_21_4 (
            .in0(_gnd_net_),
            .in1(N__42118),
            .in2(N__42999),
            .in3(N__39625),
            .lcout(n3020),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_11_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_11_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_11_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1987_3_lut_LC_11_21_5 (
            .in0(_gnd_net_),
            .in1(N__39619),
            .in2(N__44668),
            .in3(N__42964),
            .lcout(n3019),
            .ltout(n3019_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_11_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_11_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_11_21_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2054_3_lut_LC_11_21_6 (
            .in0(_gnd_net_),
            .in1(N__45364),
            .in2(N__39613),
            .in3(N__48995),
            .lcout(n3118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_11_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_11_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_11_21_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i2060_3_lut_LC_11_21_7 (
            .in0(N__48999),
            .in1(N__45028),
            .in2(N__45054),
            .in3(_gnd_net_),
            .lcout(n3124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_11_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_11_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_11_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1983_3_lut_LC_11_22_0 (
            .in0(_gnd_net_),
            .in1(N__42532),
            .in2(N__39610),
            .in3(N__42971),
            .lcout(n3015),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_11_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_11_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_11_22_1.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1981_3_lut_LC_11_22_1 (
            .in0(N__44920),
            .in1(N__39709),
            .in2(N__43001),
            .in3(_gnd_net_),
            .lcout(n3013),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_11_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_11_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_11_22_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2065_3_lut_LC_11_22_2 (
            .in0(_gnd_net_),
            .in1(N__45225),
            .in2(N__45205),
            .in3(N__49019),
            .lcout(n3129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_11_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_11_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_11_22_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1984_3_lut_LC_11_22_3 (
            .in0(_gnd_net_),
            .in1(N__39703),
            .in2(N__43000),
            .in3(N__42090),
            .lcout(n3016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_11_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_11_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_11_22_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1912_3_lut_LC_11_22_4 (
            .in0(_gnd_net_),
            .in1(N__48429),
            .in2(N__49375),
            .in3(N__48397),
            .lcout(n2912),
            .ltout(n2912_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_11_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_11_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_11_22_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1979_3_lut_LC_11_22_5 (
            .in0(N__42975),
            .in1(_gnd_net_),
            .in2(N__39697),
            .in3(N__39694),
            .lcout(n3011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_11_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_11_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_11_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1975_3_lut_LC_11_22_6 (
            .in0(_gnd_net_),
            .in1(N__40470),
            .in2(N__39688),
            .in3(N__42979),
            .lcout(n3007),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_11_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_11_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_11_23_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1980_3_lut_LC_11_23_0 (
            .in0(_gnd_net_),
            .in1(N__42607),
            .in2(N__39676),
            .in3(N__43003),
            .lcout(n3012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_11_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_11_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_11_23_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1976_3_lut_LC_11_23_2 (
            .in0(_gnd_net_),
            .in1(N__42262),
            .in2(N__39667),
            .in3(N__43005),
            .lcout(n3008),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_11_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_11_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_11_23_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2116_3_lut_LC_11_23_3 (
            .in0(_gnd_net_),
            .in1(N__51632),
            .in2(N__51613),
            .in3(N__50086),
            .lcout(n3212),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_11_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_11_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_11_23_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1978_3_lut_LC_11_23_4 (
            .in0(_gnd_net_),
            .in1(N__39658),
            .in2(N__40549),
            .in3(N__43004),
            .lcout(n3010),
            .ltout(n3010_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_11_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_11_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_11_23_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2045_3_lut_LC_11_23_5 (
            .in0(_gnd_net_),
            .in1(N__45610),
            .in2(N__39766),
            .in3(N__49020),
            .lcout(n3109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12618_1_lut_LC_11_23_6.C_ON=1'b0;
    defparam i12618_1_lut_LC_11_23_6.SEQ_MODE=4'b0000;
    defparam i12618_1_lut_LC_11_23_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12618_1_lut_LC_11_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43002),
            .lcout(n15090),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_11_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_11_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_11_23_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2120_3_lut_LC_11_23_7 (
            .in0(_gnd_net_),
            .in1(N__51775),
            .in2(N__51805),
            .in3(N__50085),
            .lcout(n3216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_157_LC_11_24_0.C_ON=1'b0;
    defparam i1_4_lut_adj_157_LC_11_24_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_157_LC_11_24_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_157_LC_11_24_0 (
            .in0(N__43478),
            .in1(N__43433),
            .in2(N__43401),
            .in3(N__39730),
            .lcout(),
            .ltout(n14392_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_160_LC_11_24_1.C_ON=1'b0;
    defparam i1_4_lut_adj_160_LC_11_24_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_160_LC_11_24_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_160_LC_11_24_1 (
            .in0(N__43337),
            .in1(N__43298),
            .in2(N__39745),
            .in3(N__49428),
            .lcout(n14398),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_155_LC_11_24_2.C_ON=1'b0;
    defparam i1_4_lut_adj_155_LC_11_24_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_155_LC_11_24_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_155_LC_11_24_2 (
            .in0(N__43199),
            .in1(N__43229),
            .in2(N__45802),
            .in3(N__39742),
            .lcout(),
            .ltout(n14380_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_156_LC_11_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_156_LC_11_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_156_LC_11_24_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_156_LC_11_24_3 (
            .in0(N__43167),
            .in1(N__43132),
            .in2(N__39733),
            .in3(N__49930),
            .lcout(n14386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12724_4_lut_LC_11_24_4.C_ON=1'b0;
    defparam i12724_4_lut_LC_11_24_4.SEQ_MODE=4'b0000;
    defparam i12724_4_lut_LC_11_24_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12724_4_lut_LC_11_24_4 (
            .in0(N__51909),
            .in1(N__43619),
            .in2(N__43668),
            .in3(N__39724),
            .lcout(n3237),
            .ltout(n3237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_11_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_11_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2176_3_lut_LC_11_24_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i2176_3_lut_LC_11_24_5 (
            .in0(N__43620),
            .in1(_gnd_net_),
            .in2(N__39718),
            .in3(N__43606),
            .lcout(n61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_141_LC_11_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_141_LC_11_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_141_LC_11_25_1.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_141_LC_11_25_1 (
            .in0(N__43453),
            .in1(N__43482),
            .in2(N__49608),
            .in3(N__40618),
            .lcout(),
            .ltout(n13856_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_142_LC_11_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_142_LC_11_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_142_LC_11_25_2.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_142_LC_11_25_2 (
            .in0(N__43417),
            .in1(N__43441),
            .in2(N__39817),
            .in3(N__49581),
            .lcout(),
            .ltout(n13858_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_143_LC_11_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_143_LC_11_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_143_LC_11_25_3.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_143_LC_11_25_3 (
            .in0(N__49582),
            .in1(N__43375),
            .in2(N__39814),
            .in3(N__43394),
            .lcout(),
            .ltout(n13860_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_144_LC_11_25_4.C_ON=1'b0;
    defparam i1_4_lut_adj_144_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_144_LC_11_25_4.LUT_INIT=16'b1111111011110010;
    LogicCell40 i1_4_lut_adj_144_LC_11_25_4 (
            .in0(N__43360),
            .in1(N__49583),
            .in2(N__39811),
            .in3(N__49429),
            .lcout(),
            .ltout(n13862_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_145_LC_11_25_5.C_ON=1'b0;
    defparam i1_4_lut_adj_145_LC_11_25_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_145_LC_11_25_5.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_145_LC_11_25_5 (
            .in0(N__49584),
            .in1(N__43321),
            .in2(N__39808),
            .in3(N__43341),
            .lcout(),
            .ltout(n13864_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_146_LC_11_25_6.C_ON=1'b0;
    defparam i1_4_lut_adj_146_LC_11_25_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_146_LC_11_25_6.LUT_INIT=16'b1111111011110010;
    LogicCell40 i1_4_lut_adj_146_LC_11_25_6 (
            .in0(N__43282),
            .in1(N__49585),
            .in2(N__39805),
            .in3(N__43302),
            .lcout(n13866),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i6_1_lut_LC_11_25_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i6_1_lut_LC_11_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i6_1_lut_LC_11_25_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i6_1_lut_LC_11_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39796),
            .lcout(n20_adj_550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i9_1_lut_LC_11_26_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i9_1_lut_LC_11_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i9_1_lut_LC_11_26_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i9_1_lut_LC_11_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39784),
            .lcout(n17_adj_553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i12_1_lut_LC_11_26_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i12_1_lut_LC_11_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i12_1_lut_LC_11_26_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i12_1_lut_LC_11_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39775),
            .lcout(n14_adj_556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i8_1_lut_LC_11_26_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i8_1_lut_LC_11_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i8_1_lut_LC_11_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i8_1_lut_LC_11_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39877),
            .lcout(n18_adj_552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i22_1_lut_LC_11_26_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_11_26_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_11_26_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i22_1_lut_LC_11_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46347),
            .lcout(n4_adj_570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i2_1_lut_LC_11_26_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i2_1_lut_LC_11_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i2_1_lut_LC_11_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i2_1_lut_LC_11_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39865),
            .lcout(n24_adj_546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_77_LC_11_27_0.C_ON=1'b0;
    defparam i1_4_lut_adj_77_LC_11_27_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_77_LC_11_27_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_77_LC_11_27_0 (
            .in0(N__39892),
            .in1(N__56388),
            .in2(N__56174),
            .in3(N__55729),
            .lcout(n4_adj_698),
            .ltout(n4_adj_698_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12245_2_lut_4_lut_LC_11_27_1.C_ON=1'b0;
    defparam i12245_2_lut_4_lut_LC_11_27_1.SEQ_MODE=4'b0000;
    defparam i12245_2_lut_4_lut_LC_11_27_1.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12245_2_lut_4_lut_LC_11_27_1 (
            .in0(N__41055),
            .in1(N__56254),
            .in2(N__39853),
            .in3(N__40722),
            .lcout(n14700),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12282_2_lut_4_lut_LC_11_27_2.C_ON=1'b0;
    defparam i12282_2_lut_4_lut_LC_11_27_2.SEQ_MODE=4'b0000;
    defparam i12282_2_lut_4_lut_LC_11_27_2.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12282_2_lut_4_lut_LC_11_27_2 (
            .in0(N__56252),
            .in1(N__41057),
            .in2(N__41140),
            .in3(N__43546),
            .lcout(n14692),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12293_2_lut_4_lut_LC_11_27_3.C_ON=1'b0;
    defparam i12293_2_lut_4_lut_LC_11_27_3.SEQ_MODE=4'b0000;
    defparam i12293_2_lut_4_lut_LC_11_27_3.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12293_2_lut_4_lut_LC_11_27_3 (
            .in0(N__41059),
            .in1(N__41132),
            .in2(N__40831),
            .in3(N__56256),
            .lcout(n14687),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12283_2_lut_4_lut_LC_11_27_4.C_ON=1'b0;
    defparam i12283_2_lut_4_lut_LC_11_27_4.SEQ_MODE=4'b0000;
    defparam i12283_2_lut_4_lut_LC_11_27_4.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12283_2_lut_4_lut_LC_11_27_4 (
            .in0(N__56253),
            .in1(N__41058),
            .in2(N__41141),
            .in3(N__43527),
            .lcout(n14693),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12281_2_lut_4_lut_LC_11_27_5.C_ON=1'b0;
    defparam i12281_2_lut_4_lut_LC_11_27_5.SEQ_MODE=4'b0000;
    defparam i12281_2_lut_4_lut_LC_11_27_5.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12281_2_lut_4_lut_LC_11_27_5 (
            .in0(N__41056),
            .in1(N__41131),
            .in2(N__40675),
            .in3(N__56255),
            .lcout(n14691),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i21_LC_11_27_6.C_ON=1'b0;
    defparam pwm_setpoint_i21_LC_11_27_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i21_LC_11_27_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i21_LC_11_27_6 (
            .in0(N__55696),
            .in1(N__46348),
            .in2(_gnd_net_),
            .in3(N__43876),
            .lcout(pwm_setpoint_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i15_1_lut_LC_11_27_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i15_1_lut_LC_11_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i15_1_lut_LC_11_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i15_1_lut_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39928),
            .lcout(n11_adj_559),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i9_2_lut_LC_11_28_1.C_ON=1'b0;
    defparam LessThan_275_i9_2_lut_LC_11_28_1.SEQ_MODE=4'b0000;
    defparam LessThan_275_i9_2_lut_LC_11_28_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i9_2_lut_LC_11_28_1 (
            .in0(_gnd_net_),
            .in1(N__40797),
            .in2(_gnd_net_),
            .in3(N__39984),
            .lcout(n9_adj_608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i17_1_lut_LC_11_28_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i17_1_lut_LC_11_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i17_1_lut_LC_11_28_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i17_1_lut_LC_11_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39916),
            .lcout(n9_adj_561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i0_LC_11_28_3.C_ON=1'b0;
    defparam commutation_state_prev_i0_LC_11_28_3.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i0_LC_11_28_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 commutation_state_prev_i0_LC_11_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56250),
            .lcout(commutation_state_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i19_1_lut_LC_11_28_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i19_1_lut_LC_11_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i19_1_lut_LC_11_28_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i19_1_lut_LC_11_28_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39904),
            .lcout(n7_adj_563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i2_LC_11_28_7.C_ON=1'b0;
    defparam commutation_state_prev_i2_LC_11_28_7.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i2_LC_11_28_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i2_LC_11_28_7 (
            .in0(N__56145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.pwm_counter_635__i0_LC_11_29_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i0_LC_11_29_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i0_LC_11_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i0_LC_11_29_0  (
            .in0(_gnd_net_),
            .in1(N__46524),
            .in2(_gnd_net_),
            .in3(N__39886),
            .lcout(pwm_counter_0),
            .ltout(),
            .carryin(bfn_11_29_0_),
            .carryout(\PWM.n12686 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i1_LC_11_29_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i1_LC_11_29_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i1_LC_11_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i1_LC_11_29_1  (
            .in0(_gnd_net_),
            .in1(N__46542),
            .in2(_gnd_net_),
            .in3(N__39883),
            .lcout(pwm_counter_1),
            .ltout(),
            .carryin(\PWM.n12686 ),
            .carryout(\PWM.n12687 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i2_LC_11_29_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i2_LC_11_29_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i2_LC_11_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i2_LC_11_29_2  (
            .in0(_gnd_net_),
            .in1(N__40782),
            .in2(_gnd_net_),
            .in3(N__39880),
            .lcout(pwm_counter_2),
            .ltout(),
            .carryin(\PWM.n12687 ),
            .carryout(\PWM.n12688 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i3_LC_11_29_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i3_LC_11_29_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i3_LC_11_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i3_LC_11_29_3  (
            .in0(_gnd_net_),
            .in1(N__40768),
            .in2(_gnd_net_),
            .in3(N__39988),
            .lcout(pwm_counter_3),
            .ltout(),
            .carryin(\PWM.n12688 ),
            .carryout(\PWM.n12689 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i4_LC_11_29_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i4_LC_11_29_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i4_LC_11_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i4_LC_11_29_4  (
            .in0(_gnd_net_),
            .in1(N__39985),
            .in2(_gnd_net_),
            .in3(N__39973),
            .lcout(pwm_counter_4),
            .ltout(),
            .carryin(\PWM.n12689 ),
            .carryout(\PWM.n12690 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i5_LC_11_29_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i5_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i5_LC_11_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i5_LC_11_29_5  (
            .in0(_gnd_net_),
            .in1(N__41190),
            .in2(_gnd_net_),
            .in3(N__39970),
            .lcout(pwm_counter_5),
            .ltout(),
            .carryin(\PWM.n12690 ),
            .carryout(\PWM.n12691 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i6_LC_11_29_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i6_LC_11_29_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i6_LC_11_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i6_LC_11_29_6  (
            .in0(_gnd_net_),
            .in1(N__41169),
            .in2(_gnd_net_),
            .in3(N__39967),
            .lcout(pwm_counter_6),
            .ltout(),
            .carryin(\PWM.n12691 ),
            .carryout(\PWM.n12692 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i7_LC_11_29_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i7_LC_11_29_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i7_LC_11_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i7_LC_11_29_7  (
            .in0(_gnd_net_),
            .in1(N__47029),
            .in2(_gnd_net_),
            .in3(N__39964),
            .lcout(pwm_counter_7),
            .ltout(),
            .carryin(\PWM.n12692 ),
            .carryout(\PWM.n12693 ),
            .clk(N__56070),
            .ce(),
            .sr(N__41423));
    defparam \PWM.pwm_counter_635__i8_LC_11_30_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i8_LC_11_30_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i8_LC_11_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i8_LC_11_30_0  (
            .in0(_gnd_net_),
            .in1(N__41533),
            .in2(_gnd_net_),
            .in3(N__39961),
            .lcout(pwm_counter_8),
            .ltout(),
            .carryin(bfn_11_30_0_),
            .carryout(\PWM.n12694 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i9_LC_11_30_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i9_LC_11_30_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i9_LC_11_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i9_LC_11_30_1  (
            .in0(_gnd_net_),
            .in1(N__41341),
            .in2(_gnd_net_),
            .in3(N__39958),
            .lcout(pwm_counter_9),
            .ltout(),
            .carryin(\PWM.n12694 ),
            .carryout(\PWM.n12695 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i10_LC_11_30_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i10_LC_11_30_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i10_LC_11_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i10_LC_11_30_2  (
            .in0(_gnd_net_),
            .in1(N__40975),
            .in2(_gnd_net_),
            .in3(N__39955),
            .lcout(pwm_counter_10),
            .ltout(),
            .carryin(\PWM.n12695 ),
            .carryout(\PWM.n12696 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i11_LC_11_30_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i11_LC_11_30_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i11_LC_11_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i11_LC_11_30_3  (
            .in0(_gnd_net_),
            .in1(N__39951),
            .in2(_gnd_net_),
            .in3(N__39931),
            .lcout(pwm_counter_11),
            .ltout(),
            .carryin(\PWM.n12696 ),
            .carryout(\PWM.n12697 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i12_LC_11_30_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i12_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i12_LC_11_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i12_LC_11_30_4  (
            .in0(_gnd_net_),
            .in1(N__41712),
            .in2(_gnd_net_),
            .in3(N__40030),
            .lcout(pwm_counter_12),
            .ltout(),
            .carryin(\PWM.n12697 ),
            .carryout(\PWM.n12698 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i13_LC_11_30_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i13_LC_11_30_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i13_LC_11_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i13_LC_11_30_5  (
            .in0(_gnd_net_),
            .in1(N__46742),
            .in2(_gnd_net_),
            .in3(N__40027),
            .lcout(pwm_counter_13),
            .ltout(),
            .carryin(\PWM.n12698 ),
            .carryout(\PWM.n12699 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i14_LC_11_30_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i14_LC_11_30_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i14_LC_11_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i14_LC_11_30_6  (
            .in0(_gnd_net_),
            .in1(N__46767),
            .in2(_gnd_net_),
            .in3(N__40024),
            .lcout(pwm_counter_14),
            .ltout(),
            .carryin(\PWM.n12699 ),
            .carryout(\PWM.n12700 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i15_LC_11_30_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i15_LC_11_30_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i15_LC_11_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i15_LC_11_30_7  (
            .in0(_gnd_net_),
            .in1(N__44030),
            .in2(_gnd_net_),
            .in3(N__40021),
            .lcout(pwm_counter_15),
            .ltout(),
            .carryin(\PWM.n12700 ),
            .carryout(\PWM.n12701 ),
            .clk(N__56074),
            .ce(),
            .sr(N__41440));
    defparam \PWM.pwm_counter_635__i16_LC_11_31_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i16_LC_11_31_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i16_LC_11_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i16_LC_11_31_0  (
            .in0(_gnd_net_),
            .in1(N__46828),
            .in2(_gnd_net_),
            .in3(N__40018),
            .lcout(pwm_counter_16),
            .ltout(),
            .carryin(bfn_11_31_0_),
            .carryout(\PWM.n12702 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i17_LC_11_31_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i17_LC_11_31_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i17_LC_11_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i17_LC_11_31_1  (
            .in0(_gnd_net_),
            .in1(N__44270),
            .in2(_gnd_net_),
            .in3(N__40015),
            .lcout(pwm_counter_17),
            .ltout(),
            .carryin(\PWM.n12702 ),
            .carryout(\PWM.n12703 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i18_LC_11_31_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i18_LC_11_31_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i18_LC_11_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i18_LC_11_31_2  (
            .in0(_gnd_net_),
            .in1(N__44004),
            .in2(_gnd_net_),
            .in3(N__40012),
            .lcout(pwm_counter_18),
            .ltout(),
            .carryin(\PWM.n12703 ),
            .carryout(\PWM.n12704 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i19_LC_11_31_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i19_LC_11_31_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i19_LC_11_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i19_LC_11_31_3  (
            .in0(_gnd_net_),
            .in1(N__41401),
            .in2(_gnd_net_),
            .in3(N__40009),
            .lcout(pwm_counter_19),
            .ltout(),
            .carryin(\PWM.n12704 ),
            .carryout(\PWM.n12705 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i20_LC_11_31_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i20_LC_11_31_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i20_LC_11_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i20_LC_11_31_4  (
            .in0(_gnd_net_),
            .in1(N__40006),
            .in2(_gnd_net_),
            .in3(N__39991),
            .lcout(pwm_counter_20),
            .ltout(),
            .carryin(\PWM.n12705 ),
            .carryout(\PWM.n12706 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i21_LC_11_31_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i21_LC_11_31_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i21_LC_11_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i21_LC_11_31_5  (
            .in0(_gnd_net_),
            .in1(N__40169),
            .in2(_gnd_net_),
            .in3(N__40141),
            .lcout(pwm_counter_21),
            .ltout(),
            .carryin(\PWM.n12706 ),
            .carryout(\PWM.n12707 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i22_LC_11_31_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i22_LC_11_31_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i22_LC_11_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i22_LC_11_31_6  (
            .in0(_gnd_net_),
            .in1(N__40134),
            .in2(_gnd_net_),
            .in3(N__40114),
            .lcout(pwm_counter_22),
            .ltout(),
            .carryin(\PWM.n12707 ),
            .carryout(\PWM.n12708 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i23_LC_11_31_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i23_LC_11_31_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i23_LC_11_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i23_LC_11_31_7  (
            .in0(_gnd_net_),
            .in1(N__44062),
            .in2(_gnd_net_),
            .in3(N__40111),
            .lcout(pwm_counter_23),
            .ltout(),
            .carryin(\PWM.n12708 ),
            .carryout(\PWM.n12709 ),
            .clk(N__56077),
            .ce(),
            .sr(N__41429));
    defparam \PWM.pwm_counter_635__i24_LC_11_32_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i24_LC_11_32_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i24_LC_11_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i24_LC_11_32_0  (
            .in0(_gnd_net_),
            .in1(N__40108),
            .in2(_gnd_net_),
            .in3(N__40096),
            .lcout(pwm_counter_24),
            .ltout(),
            .carryin(bfn_11_32_0_),
            .carryout(\PWM.n12710 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i25_LC_11_32_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i25_LC_11_32_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i25_LC_11_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i25_LC_11_32_1  (
            .in0(_gnd_net_),
            .in1(N__40093),
            .in2(_gnd_net_),
            .in3(N__40081),
            .lcout(pwm_counter_25),
            .ltout(),
            .carryin(\PWM.n12710 ),
            .carryout(\PWM.n12711 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i26_LC_11_32_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i26_LC_11_32_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i26_LC_11_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i26_LC_11_32_2  (
            .in0(_gnd_net_),
            .in1(N__40078),
            .in2(_gnd_net_),
            .in3(N__40066),
            .lcout(pwm_counter_26),
            .ltout(),
            .carryin(\PWM.n12711 ),
            .carryout(\PWM.n12712 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i27_LC_11_32_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i27_LC_11_32_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i27_LC_11_32_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i27_LC_11_32_3  (
            .in0(_gnd_net_),
            .in1(N__40062),
            .in2(_gnd_net_),
            .in3(N__40048),
            .lcout(pwm_counter_27),
            .ltout(),
            .carryin(\PWM.n12712 ),
            .carryout(\PWM.n12713 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i28_LC_11_32_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i28_LC_11_32_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i28_LC_11_32_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i28_LC_11_32_4  (
            .in0(_gnd_net_),
            .in1(N__40045),
            .in2(_gnd_net_),
            .in3(N__40033),
            .lcout(pwm_counter_28),
            .ltout(),
            .carryin(\PWM.n12713 ),
            .carryout(\PWM.n12714 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i29_LC_11_32_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i29_LC_11_32_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i29_LC_11_32_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i29_LC_11_32_5  (
            .in0(_gnd_net_),
            .in1(N__40228),
            .in2(_gnd_net_),
            .in3(N__40216),
            .lcout(pwm_counter_29),
            .ltout(),
            .carryin(\PWM.n12714 ),
            .carryout(\PWM.n12715 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i30_LC_11_32_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_635__i30_LC_11_32_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i30_LC_11_32_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i30_LC_11_32_6  (
            .in0(_gnd_net_),
            .in1(N__40213),
            .in2(_gnd_net_),
            .in3(N__40201),
            .lcout(pwm_counter_30),
            .ltout(),
            .carryin(\PWM.n12715 ),
            .carryout(\PWM.n12716 ),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam \PWM.pwm_counter_635__i31_LC_11_32_7 .C_ON=1'b0;
    defparam \PWM.pwm_counter_635__i31_LC_11_32_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_635__i31_LC_11_32_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_635__i31_LC_11_32_7  (
            .in0(_gnd_net_),
            .in1(N__41475),
            .in2(_gnd_net_),
            .in3(N__40198),
            .lcout(pwm_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56081),
            .ce(),
            .sr(N__41436));
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_12_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_12_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_2_lut_LC_12_17_0 (
            .in0(_gnd_net_),
            .in1(N__47683),
            .in2(_gnd_net_),
            .in3(N__40195),
            .lcout(n2801),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(n12386),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_12_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_12_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_3_lut_LC_12_17_1 (
            .in0(_gnd_net_),
            .in1(N__53560),
            .in2(N__44385),
            .in3(N__40192),
            .lcout(n2800),
            .ltout(),
            .carryin(n12386),
            .carryout(n12387),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_12_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_12_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_4_lut_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44346),
            .in3(N__40189),
            .lcout(n2799),
            .ltout(),
            .carryin(n12387),
            .carryout(n12388),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_12_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_12_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_5_lut_LC_12_17_3 (
            .in0(_gnd_net_),
            .in1(N__53561),
            .in2(N__41985),
            .in3(N__40186),
            .lcout(n2798),
            .ltout(),
            .carryin(n12388),
            .carryout(n12389),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_12_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_12_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_6_lut_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41856),
            .in3(N__40183),
            .lcout(n2797),
            .ltout(),
            .carryin(n12389),
            .carryout(n12390),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_12_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_12_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_7_lut_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44430),
            .in3(N__40180),
            .lcout(n2796),
            .ltout(),
            .carryin(n12390),
            .carryout(n12391),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_12_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_12_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_12_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_8_lut_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(N__53569),
            .in2(N__41962),
            .in3(N__40282),
            .lcout(n2795),
            .ltout(),
            .carryin(n12391),
            .carryout(n12392),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_12_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_12_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_12_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_9_lut_LC_12_17_7 (
            .in0(_gnd_net_),
            .in1(N__53562),
            .in2(N__44193),
            .in3(N__40279),
            .lcout(n2794),
            .ltout(),
            .carryin(n12392),
            .carryout(n12393),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_12_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_12_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_12_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_10_lut_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(N__53839),
            .in2(N__44499),
            .in3(N__40276),
            .lcout(n2793),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(n12394),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_12_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_12_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_12_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_11_lut_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__53563),
            .in2(N__41641),
            .in3(N__40273),
            .lcout(n2792),
            .ltout(),
            .carryin(n12394),
            .carryout(n12395),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_12_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_12_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_12_lut_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(N__53840),
            .in2(N__42184),
            .in3(N__40270),
            .lcout(n2791),
            .ltout(),
            .carryin(n12395),
            .carryout(n12396),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_12_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_12_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_12_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_13_lut_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(N__53564),
            .in2(N__41673),
            .in3(N__40267),
            .lcout(n2790),
            .ltout(),
            .carryin(n12396),
            .carryout(n12397),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_12_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_12_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_12_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_14_lut_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(N__53841),
            .in2(N__41886),
            .in3(N__40264),
            .lcout(n2789),
            .ltout(),
            .carryin(n12397),
            .carryout(n12398),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_12_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_12_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_15_lut_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__53565),
            .in2(N__40261),
            .in3(N__40234),
            .lcout(n2788),
            .ltout(),
            .carryin(n12398),
            .carryout(n12399),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_12_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_12_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_16_lut_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(N__41919),
            .in2(N__53877),
            .in3(N__40231),
            .lcout(n2787),
            .ltout(),
            .carryin(n12399),
            .carryout(n12400),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_12_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_12_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_17_lut_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(N__42138),
            .in2(N__54308),
            .in3(N__40381),
            .lcout(n2786),
            .ltout(),
            .carryin(n12400),
            .carryout(n12401),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_12_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_12_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_12_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_18_lut_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(N__40377),
            .in2(N__54336),
            .in3(N__40345),
            .lcout(n2785),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(n12402),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_12_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_12_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_12_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_19_lut_LC_12_19_1 (
            .in0(_gnd_net_),
            .in1(N__40342),
            .in2(N__54767),
            .in3(N__40309),
            .lcout(n2784),
            .ltout(),
            .carryin(n12402),
            .carryout(n12403),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_12_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_12_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_12_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_20_lut_LC_12_19_2 (
            .in0(_gnd_net_),
            .in1(N__44167),
            .in2(N__54337),
            .in3(N__40306),
            .lcout(n2783),
            .ltout(),
            .carryin(n12403),
            .carryout(n12404),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_12_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_12_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_12_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_21_lut_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(N__44111),
            .in2(N__54768),
            .in3(N__40303),
            .lcout(n2782),
            .ltout(),
            .carryin(n12404),
            .carryout(n12405),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_12_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_12_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_12_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_22_lut_LC_12_19_4 (
            .in0(_gnd_net_),
            .in1(N__41589),
            .in2(N__54338),
            .in3(N__40294),
            .lcout(n2781),
            .ltout(),
            .carryin(n12405),
            .carryout(n12406),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_12_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_12_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_23_lut_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(N__42227),
            .in2(N__54769),
            .in3(N__40291),
            .lcout(n2780),
            .ltout(),
            .carryin(n12406),
            .carryout(n12407),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_12_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_12_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_12_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_24_lut_LC_12_19_6 (
            .in0(_gnd_net_),
            .in1(N__44250),
            .in2(N__54339),
            .in3(N__40288),
            .lcout(n2779),
            .ltout(),
            .carryin(n12407),
            .carryout(n12408),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_12_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_12_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_12_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_25_lut_LC_12_19_7 (
            .in0(_gnd_net_),
            .in1(N__53890),
            .in2(N__42309),
            .in3(N__40285),
            .lcout(n2778),
            .ltout(),
            .carryin(n12408),
            .carryout(n12409),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_12_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_12_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_12_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_26_lut_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(N__41567),
            .in2(N__54770),
            .in3(N__40429),
            .lcout(n2777),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(n12410),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_12_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_12_20_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1838_27_lut_LC_12_20_1 (
            .in0(N__53891),
            .in1(N__42273),
            .in2(N__42028),
            .in3(N__40426),
            .lcout(n2808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_12_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_12_20_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2043_3_lut_LC_12_20_3 (
            .in0(_gnd_net_),
            .in1(N__45588),
            .in2(N__45562),
            .in3(N__49074),
            .lcout(n3107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_12_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_12_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_12_20_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1911_3_lut_LC_12_20_4 (
            .in0(_gnd_net_),
            .in1(N__48377),
            .in2(N__48355),
            .in3(N__49367),
            .lcout(n2911),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_12_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_12_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_12_20_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1985_3_lut_LC_12_20_6 (
            .in0(_gnd_net_),
            .in1(N__40423),
            .in2(N__42063),
            .in3(N__42980),
            .lcout(n3017),
            .ltout(n3017_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_12_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_12_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_12_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2052_3_lut_LC_12_20_7 (
            .in0(_gnd_net_),
            .in1(N__45289),
            .in2(N__40411),
            .in3(N__49073),
            .lcout(n3116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_12_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_12_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_12_21_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1977_3_lut_LC_12_21_0 (
            .in0(N__47103),
            .in1(_gnd_net_),
            .in2(N__42993),
            .in3(N__40408),
            .lcout(n3009),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_12_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_12_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_12_21_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1993_3_lut_LC_12_21_1 (
            .in0(N__44698),
            .in1(_gnd_net_),
            .in2(N__40396),
            .in3(N__42940),
            .lcout(n3025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_41_LC_12_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_41_LC_12_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_41_LC_12_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_41_LC_12_21_2 (
            .in0(N__44912),
            .in1(N__42594),
            .in2(N__47275),
            .in3(N__42505),
            .lcout(),
            .ltout(n13948_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_42_LC_12_21_3.C_ON=1'b0;
    defparam i1_4_lut_adj_42_LC_12_21_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_42_LC_12_21_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_42_LC_12_21_3 (
            .in0(N__40533),
            .in1(N__40518),
            .in2(N__40507),
            .in3(N__47102),
            .lcout(),
            .ltout(n13954_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12622_4_lut_LC_12_21_4.C_ON=1'b0;
    defparam i12622_4_lut_LC_12_21_4.SEQ_MODE=4'b0000;
    defparam i12622_4_lut_LC_12_21_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12622_4_lut_LC_12_21_4 (
            .in0(N__42248),
            .in1(N__48759),
            .in2(N__40504),
            .in3(N__40466),
            .lcout(n2940),
            .ltout(n2940_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_12_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_12_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_12_21_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1999_3_lut_LC_12_21_5 (
            .in0(N__40501),
            .in1(_gnd_net_),
            .in2(N__40492),
            .in3(N__47460),
            .lcout(n3031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_12_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_12_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_12_21_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1996_3_lut_LC_12_21_7 (
            .in0(_gnd_net_),
            .in1(N__47313),
            .in2(N__40489),
            .in3(N__42941),
            .lcout(n3028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_33_LC_12_22_0.C_ON=1'b0;
    defparam i1_4_lut_adj_33_LC_12_22_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_33_LC_12_22_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_33_LC_12_22_0 (
            .in0(N__45705),
            .in1(N__49463),
            .in2(N__45668),
            .in3(N__40561),
            .lcout(),
            .ltout(n14340_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_34_LC_12_22_1.C_ON=1'b0;
    defparam i1_4_lut_adj_34_LC_12_22_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_34_LC_12_22_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_34_LC_12_22_1 (
            .in0(N__45621),
            .in1(N__49173),
            .in2(N__40477),
            .in3(N__43015),
            .lcout(n14344),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_12_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_12_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_12_22_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1908_3_lut_LC_12_22_2 (
            .in0(N__48823),
            .in1(_gnd_net_),
            .in2(N__48863),
            .in3(N__49371),
            .lcout(n2908),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12655_4_lut_LC_12_22_4.C_ON=1'b0;
    defparam i12655_4_lut_LC_12_22_4.SEQ_MODE=4'b0000;
    defparam i12655_4_lut_LC_12_22_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12655_4_lut_LC_12_22_4 (
            .in0(N__45578),
            .in1(N__45533),
            .in2(N__45940),
            .in3(N__40450),
            .lcout(n3039),
            .ltout(n3039_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_12_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_12_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_12_22_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2059_3_lut_LC_12_22_5 (
            .in0(_gnd_net_),
            .in1(N__44992),
            .in2(N__40444),
            .in3(N__45012),
            .lcout(n3123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_32_LC_12_22_6.C_ON=1'b0;
    defparam i1_4_lut_adj_32_LC_12_22_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_32_LC_12_22_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_32_LC_12_22_6 (
            .in0(N__49118),
            .in1(N__45303),
            .in2(N__42193),
            .in3(N__40570),
            .lcout(n14334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12651_1_lut_LC_12_22_7.C_ON=1'b0;
    defparam i12651_1_lut_LC_12_22_7.SEQ_MODE=4'b0000;
    defparam i12651_1_lut_LC_12_22_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12651_1_lut_LC_12_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49079),
            .in3(_gnd_net_),
            .lcout(n15123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_12_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_12_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_12_23_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2047_3_lut_LC_12_23_0 (
            .in0(N__45670),
            .in1(N__45646),
            .in2(N__49039),
            .in3(_gnd_net_),
            .lcout(n3111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_12_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_12_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_12_23_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2057_3_lut_LC_12_23_1 (
            .in0(_gnd_net_),
            .in1(N__45495),
            .in2(N__45475),
            .in3(N__48980),
            .lcout(n3121),
            .ltout(n3121_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_12_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_12_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_12_23_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2124_3_lut_LC_12_23_2 (
            .in0(_gnd_net_),
            .in1(N__51289),
            .in2(N__40555),
            .in3(N__50073),
            .lcout(n3220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_12_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_12_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_12_23_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2049_3_lut_LC_12_23_3 (
            .in0(_gnd_net_),
            .in1(N__45721),
            .in2(N__45736),
            .in3(N__48981),
            .lcout(n3113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_12_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_12_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_12_23_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2121_3_lut_LC_12_23_4 (
            .in0(_gnd_net_),
            .in1(N__51852),
            .in2(N__51826),
            .in3(N__50077),
            .lcout(n3217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_12_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_12_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_12_23_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2127_3_lut_LC_12_23_5 (
            .in0(N__51418),
            .in1(_gnd_net_),
            .in2(N__50105),
            .in3(N__51444),
            .lcout(n3223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_12_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_12_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_12_23_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2048_3_lut_LC_12_23_6 (
            .in0(_gnd_net_),
            .in1(N__45682),
            .in2(N__49040),
            .in3(N__45704),
            .lcout(n3112),
            .ltout(n3112_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_12_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_12_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_12_23_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i2115_3_lut_LC_12_23_7 (
            .in0(N__50078),
            .in1(_gnd_net_),
            .in2(N__40552),
            .in3(N__51571),
            .lcout(n3211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_12_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_12_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_12_24_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2195_3_lut_LC_12_24_0 (
            .in0(_gnd_net_),
            .in1(N__45766),
            .in2(N__43042),
            .in3(N__49563),
            .lcout(),
            .ltout(n23_adj_707_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_132_LC_12_24_1.C_ON=1'b0;
    defparam i1_4_lut_adj_132_LC_12_24_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_132_LC_12_24_1.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_132_LC_12_24_1 (
            .in0(N__49565),
            .in1(N__43264),
            .in2(N__40600),
            .in3(N__45871),
            .lcout(n13828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_12_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_12_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2194_3_lut_LC_12_24_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2194_3_lut_LC_12_24_2 (
            .in0(_gnd_net_),
            .in1(N__46134),
            .in2(N__43030),
            .in3(N__49564),
            .lcout(),
            .ltout(n25_adj_708_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_133_LC_12_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_133_LC_12_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_133_LC_12_24_3.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_133_LC_12_24_3 (
            .in0(N__49566),
            .in1(N__45837),
            .in2(N__40597),
            .in3(N__43249),
            .lcout(n13826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_131_LC_12_24_4.C_ON=1'b0;
    defparam i1_4_lut_adj_131_LC_12_24_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_131_LC_12_24_4.LUT_INIT=16'b1111101011101110;
    LogicCell40 i1_4_lut_adj_131_LC_12_24_4 (
            .in0(N__40612),
            .in1(N__43054),
            .in2(N__49402),
            .in3(N__49567),
            .lcout(),
            .ltout(n13832_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_135_LC_12_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_135_LC_12_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_135_LC_12_24_5.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_135_LC_12_24_5 (
            .in0(N__49568),
            .in1(N__43183),
            .in2(N__40594),
            .in3(N__43203),
            .lcout(),
            .ltout(n13840_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_136_LC_12_24_6.C_ON=1'b0;
    defparam i1_4_lut_adj_136_LC_12_24_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_136_LC_12_24_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_136_LC_12_24_6 (
            .in0(N__40591),
            .in1(N__40585),
            .in2(N__40579),
            .in3(N__48652),
            .lcout(n13846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i5_1_lut_LC_12_25_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_12_25_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_12_25_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i5_1_lut_LC_12_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46002),
            .lcout(n21_adj_587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_137_LC_12_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_137_LC_12_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_137_LC_12_25_1.LUT_INIT=16'b1111111110101100;
    LogicCell40 i1_4_lut_adj_137_LC_12_25_1 (
            .in0(N__43171),
            .in1(N__43141),
            .in2(N__49605),
            .in3(N__40576),
            .lcout(),
            .ltout(n13848_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_138_LC_12_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_138_LC_12_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_138_LC_12_25_2.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_138_LC_12_25_2 (
            .in0(N__43501),
            .in1(N__43131),
            .in2(N__40645),
            .in3(N__49561),
            .lcout(),
            .ltout(n13850_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_139_LC_12_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_139_LC_12_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_139_LC_12_25_3.LUT_INIT=16'b1111110011111000;
    LogicCell40 i1_4_lut_adj_139_LC_12_25_3 (
            .in0(N__40606),
            .in1(N__40642),
            .in2(N__40633),
            .in3(N__40630),
            .lcout(),
            .ltout(n13852_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_140_LC_12_25_4.C_ON=1'b0;
    defparam i1_4_lut_adj_140_LC_12_25_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_140_LC_12_25_4.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_140_LC_12_25_4 (
            .in0(N__49929),
            .in1(N__43492),
            .in2(N__40621),
            .in3(N__49562),
            .lcout(n13854),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_12_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_12_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_12_25_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2126_3_lut_LC_12_25_5 (
            .in0(_gnd_net_),
            .in1(N__51395),
            .in2(N__51367),
            .in3(N__50106),
            .lcout(n3222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_12_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_12_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2188_3_lut_LC_12_25_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2188_3_lut_LC_12_25_6 (
            .in0(_gnd_net_),
            .in1(N__43216),
            .in2(N__43240),
            .in3(N__49554),
            .lcout(n37_adj_710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_12_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_12_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2203_3_lut_LC_12_25_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2203_3_lut_LC_12_25_7 (
            .in0(_gnd_net_),
            .in1(N__42706),
            .in2(N__49604),
            .in3(N__42727),
            .lcout(n7_adj_703),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_12_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_12_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_12_26_0.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i2118_3_lut_LC_12_26_0 (
            .in0(N__50107),
            .in1(N__51685),
            .in2(N__51715),
            .in3(_gnd_net_),
            .lcout(n3214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12280_2_lut_4_lut_LC_12_26_1.C_ON=1'b0;
    defparam i12280_2_lut_4_lut_LC_12_26_1.SEQ_MODE=4'b0000;
    defparam i12280_2_lut_4_lut_LC_12_26_1.LUT_INIT=16'b0000100000000100;
    LogicCell40 i12280_2_lut_4_lut_LC_12_26_1 (
            .in0(N__56277),
            .in1(N__40925),
            .in2(N__41143),
            .in3(N__41068),
            .lcout(n14690),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9490_2_lut_LC_12_26_2.C_ON=1'b0;
    defparam i9490_2_lut_LC_12_26_2.SEQ_MODE=4'b0000;
    defparam i9490_2_lut_LC_12_26_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9490_2_lut_LC_12_26_2 (
            .in0(N__55508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55447),
            .lcout(n11202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12268_2_lut_4_lut_LC_12_26_3.C_ON=1'b0;
    defparam i12268_2_lut_4_lut_LC_12_26_3.SEQ_MODE=4'b0000;
    defparam i12268_2_lut_4_lut_LC_12_26_3.LUT_INIT=16'b0000100000000100;
    LogicCell40 i12268_2_lut_4_lut_LC_12_26_3 (
            .in0(N__56276),
            .in1(N__40893),
            .in2(N__41142),
            .in3(N__41067),
            .lcout(n14688),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i12_1_lut_LC_12_26_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_12_26_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_12_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i12_1_lut_LC_12_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46197),
            .lcout(n14_adj_580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_76_LC_12_26_5.C_ON=1'b0;
    defparam i6_4_lut_adj_76_LC_12_26_5.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_76_LC_12_26_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_76_LC_12_26_5 (
            .in0(N__41084),
            .in1(N__40892),
            .in2(N__40927),
            .in3(N__40820),
            .lcout(),
            .ltout(n14_adj_679_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_12_26_6.C_ON=1'b0;
    defparam i7_4_lut_LC_12_26_6.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_12_26_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_12_26_6 (
            .in0(N__40664),
            .in1(N__40718),
            .in2(N__40741),
            .in3(N__43507),
            .lcout(n4781),
            .ltout(n4781_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9491_1_lut_2_lut_LC_12_26_7.C_ON=1'b0;
    defparam i9491_1_lut_2_lut_LC_12_26_7.SEQ_MODE=4'b0000;
    defparam i9491_1_lut_2_lut_LC_12_26_7.LUT_INIT=16'b0000111111111111;
    LogicCell40 i9491_1_lut_2_lut_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40738),
            .in3(N__55507),
            .lcout(n1259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i0_LC_12_27_0.C_ON=1'b1;
    defparam dti_counter_633__i0_LC_12_27_0.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i0_LC_12_27_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 dti_counter_633__i0_LC_12_27_0 (
            .in0(N__40735),
            .in1(N__40729),
            .in2(N__40723),
            .in3(N__40702),
            .lcout(dti_counter_0),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(n12742),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i1_LC_12_27_1.C_ON=1'b1;
    defparam dti_counter_633__i1_LC_12_27_1.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i1_LC_12_27_1.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_633__i1_LC_12_27_1 (
            .in0(N__40699),
            .in1(N__40855),
            .in2(N__43528),
            .in3(N__40693),
            .lcout(dti_counter_1),
            .ltout(),
            .carryin(n12742),
            .carryout(n12743),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i2_LC_12_27_2.C_ON=1'b1;
    defparam dti_counter_633__i2_LC_12_27_2.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i2_LC_12_27_2.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_633__i2_LC_12_27_2 (
            .in0(N__40690),
            .in1(N__43545),
            .in2(N__40868),
            .in3(N__40684),
            .lcout(dti_counter_2),
            .ltout(),
            .carryin(n12743),
            .carryout(n12744),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i3_LC_12_27_3.C_ON=1'b1;
    defparam dti_counter_633__i3_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i3_LC_12_27_3.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_633__i3_LC_12_27_3 (
            .in0(N__40681),
            .in1(N__40859),
            .in2(N__40674),
            .in3(N__40648),
            .lcout(dti_counter_3),
            .ltout(),
            .carryin(n12744),
            .carryout(n12745),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i4_LC_12_27_4.C_ON=1'b1;
    defparam dti_counter_633__i4_LC_12_27_4.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i4_LC_12_27_4.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_633__i4_LC_12_27_4 (
            .in0(N__40936),
            .in1(N__40926),
            .in2(N__40869),
            .in3(N__40906),
            .lcout(dti_counter_4),
            .ltout(),
            .carryin(n12745),
            .carryout(n12746),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i5_LC_12_27_5.C_ON=1'b1;
    defparam dti_counter_633__i5_LC_12_27_5.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i5_LC_12_27_5.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_633__i5_LC_12_27_5 (
            .in0(N__41026),
            .in1(N__40863),
            .in2(N__41094),
            .in3(N__40903),
            .lcout(dti_counter_5),
            .ltout(),
            .carryin(n12746),
            .carryout(n12747),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i6_LC_12_27_6.C_ON=1'b1;
    defparam dti_counter_633__i6_LC_12_27_6.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i6_LC_12_27_6.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_633__i6_LC_12_27_6 (
            .in0(N__40900),
            .in1(N__40894),
            .in2(N__40870),
            .in3(N__40879),
            .lcout(dti_counter_6),
            .ltout(),
            .carryin(n12747),
            .carryout(n12748),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_633__i7_LC_12_27_7.C_ON=1'b0;
    defparam dti_counter_633__i7_LC_12_27_7.SEQ_MODE=4'b1000;
    defparam dti_counter_633__i7_LC_12_27_7.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_633__i7_LC_12_27_7 (
            .in0(N__40876),
            .in1(N__40867),
            .in2(N__40830),
            .in3(N__40834),
            .lcout(dti_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56067),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i4_LC_12_28_1.C_ON=1'b0;
    defparam pwm_setpoint_i4_LC_12_28_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i4_LC_12_28_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i4_LC_12_28_1 (
            .in0(N__55711),
            .in1(N__43714),
            .in2(_gnd_net_),
            .in3(N__46003),
            .lcout(pwm_setpoint_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56071),
            .ce(),
            .sr(_gnd_net_));
    defparam i12273_3_lut_4_lut_LC_12_28_2.C_ON=1'b0;
    defparam i12273_3_lut_4_lut_LC_12_28_2.SEQ_MODE=4'b0000;
    defparam i12273_3_lut_4_lut_LC_12_28_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i12273_3_lut_4_lut_LC_12_28_2 (
            .in0(N__41019),
            .in1(N__40749),
            .in2(N__40786),
            .in3(N__40766),
            .lcout(n14745),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i6_LC_12_28_3.C_ON=1'b0;
    defparam pwm_setpoint_i6_LC_12_28_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i6_LC_12_28_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i6_LC_12_28_3 (
            .in0(N__55712),
            .in1(N__43681),
            .in2(_gnd_net_),
            .in3(N__46321),
            .lcout(pwm_setpoint_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56071),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i3_LC_12_28_4.C_ON=1'b0;
    defparam pwm_setpoint_i3_LC_12_28_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i3_LC_12_28_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 pwm_setpoint_i3_LC_12_28_4 (
            .in0(N__43735),
            .in1(N__50197),
            .in2(_gnd_net_),
            .in3(N__55713),
            .lcout(pwm_setpoint_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56071),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i6_3_lut_3_lut_LC_12_28_5.C_ON=1'b0;
    defparam LessThan_275_i6_3_lut_3_lut_LC_12_28_5.SEQ_MODE=4'b0000;
    defparam LessThan_275_i6_3_lut_3_lut_LC_12_28_5.LUT_INIT=16'b1111010101010000;
    LogicCell40 LessThan_275_i6_3_lut_3_lut_LC_12_28_5 (
            .in0(N__40767),
            .in1(_gnd_net_),
            .in2(N__40753),
            .in3(N__41020),
            .lcout(n6_adj_606),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12279_2_lut_4_lut_LC_12_28_6.C_ON=1'b0;
    defparam i12279_2_lut_4_lut_LC_12_28_6.SEQ_MODE=4'b0000;
    defparam i12279_2_lut_4_lut_LC_12_28_6.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12279_2_lut_4_lut_LC_12_28_6 (
            .in0(N__56275),
            .in1(N__41139),
            .in2(N__41095),
            .in3(N__41060),
            .lcout(n14689),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i2_LC_12_28_7.C_ON=1'b0;
    defparam pwm_setpoint_i2_LC_12_28_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i2_LC_12_28_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i2_LC_12_28_7 (
            .in0(N__55710),
            .in1(N__43744),
            .in2(_gnd_net_),
            .in3(N__46048),
            .lcout(pwm_setpoint_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56071),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i5_LC_12_29_0.C_ON=1'b0;
    defparam pwm_setpoint_i5_LC_12_29_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i5_LC_12_29_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i5_LC_12_29_0 (
            .in0(N__55698),
            .in1(N__43699),
            .in2(_gnd_net_),
            .in3(N__45961),
            .lcout(pwm_setpoint_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i11_LC_12_29_1.C_ON=1'b0;
    defparam pwm_setpoint_i11_LC_12_29_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i11_LC_12_29_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i11_LC_12_29_1 (
            .in0(N__46198),
            .in1(N__55700),
            .in2(_gnd_net_),
            .in3(N__43798),
            .lcout(pwm_setpoint_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i12_LC_12_29_2.C_ON=1'b0;
    defparam pwm_setpoint_i12_LC_12_29_2.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i12_LC_12_29_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 pwm_setpoint_i12_LC_12_29_2 (
            .in0(N__55697),
            .in1(_gnd_net_),
            .in2(N__43789),
            .in3(N__46795),
            .lcout(pwm_setpoint_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i8_LC_12_29_3.C_ON=1'b0;
    defparam pwm_setpoint_i8_LC_12_29_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i8_LC_12_29_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 pwm_setpoint_i8_LC_12_29_3 (
            .in0(N__52732),
            .in1(N__43837),
            .in2(_gnd_net_),
            .in3(N__55701),
            .lcout(pwm_setpoint_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i8_1_lut_LC_12_29_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_12_29_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_12_29_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i8_1_lut_LC_12_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46948),
            .lcout(n18_adj_584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i21_2_lut_LC_12_29_5.C_ON=1'b0;
    defparam LessThan_275_i21_2_lut_LC_12_29_5.SEQ_MODE=4'b0000;
    defparam LessThan_275_i21_2_lut_LC_12_29_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i21_2_lut_LC_12_29_5 (
            .in0(_gnd_net_),
            .in1(N__41292),
            .in2(_gnd_net_),
            .in3(N__40973),
            .lcout(n21_adj_617),
            .ltout(n21_adj_617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12370_3_lut_LC_12_29_6.C_ON=1'b0;
    defparam i12370_3_lut_LC_12_29_6.SEQ_MODE=4'b0000;
    defparam i12370_3_lut_LC_12_29_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12370_3_lut_LC_12_29_6 (
            .in0(N__41293),
            .in1(_gnd_net_),
            .in2(N__40957),
            .in3(N__40954),
            .lcout(n14842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i10_LC_12_29_7.C_ON=1'b0;
    defparam pwm_setpoint_i10_LC_12_29_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i10_LC_12_29_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i10_LC_12_29_7 (
            .in0(N__43816),
            .in1(N__55699),
            .in2(_gnd_net_),
            .in3(N__46234),
            .lcout(pwm_setpoint_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i11_2_lut_LC_12_30_0.C_ON=1'b0;
    defparam LessThan_275_i11_2_lut_LC_12_30_0.SEQ_MODE=4'b0000;
    defparam LessThan_275_i11_2_lut_LC_12_30_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i11_2_lut_LC_12_30_0 (
            .in0(_gnd_net_),
            .in1(N__41280),
            .in2(_gnd_net_),
            .in3(N__41186),
            .lcout(n11_adj_610),
            .ltout(n11_adj_610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12256_4_lut_LC_12_30_1.C_ON=1'b0;
    defparam i12256_4_lut_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam i12256_4_lut_LC_12_30_1.LUT_INIT=16'b1111111100000001;
    LogicCell40 i12256_4_lut_LC_12_30_1 (
            .in0(N__41235),
            .in1(N__41304),
            .in2(N__41284),
            .in3(N__46713),
            .lcout(n14728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i19_LC_12_30_2.C_ON=1'b0;
    defparam pwm_setpoint_i19_LC_12_30_2.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i19_LC_12_30_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i19_LC_12_30_2 (
            .in0(N__50281),
            .in1(N__55702),
            .in2(_gnd_net_),
            .in3(N__43906),
            .lcout(pwm_setpoint_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56078),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i10_3_lut_3_lut_LC_12_30_3.C_ON=1'b0;
    defparam LessThan_275_i10_3_lut_3_lut_LC_12_30_3.SEQ_MODE=4'b0000;
    defparam LessThan_275_i10_3_lut_3_lut_LC_12_30_3.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_275_i10_3_lut_3_lut_LC_12_30_3 (
            .in0(N__41281),
            .in1(N__41271),
            .in2(_gnd_net_),
            .in3(N__41165),
            .lcout(n10_adj_609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_67_LC_12_30_5.C_ON=1'b0;
    defparam i1_2_lut_adj_67_LC_12_30_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_67_LC_12_30_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_67_LC_12_30_5 (
            .in0(_gnd_net_),
            .in1(N__41476),
            .in2(_gnd_net_),
            .in3(N__41500),
            .lcout(n4825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12332_4_lut_LC_12_30_6.C_ON=1'b0;
    defparam i12332_4_lut_LC_12_30_6.SEQ_MODE=4'b0000;
    defparam i12332_4_lut_LC_12_30_6.LUT_INIT=16'b1111110011111101;
    LogicCell40 i12332_4_lut_LC_12_30_6 (
            .in0(N__41778),
            .in1(N__41236),
            .in2(N__41221),
            .in3(N__41212),
            .lcout(n14804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i20_LC_12_30_7.C_ON=1'b0;
    defparam pwm_setpoint_i20_LC_12_30_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i20_LC_12_30_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 pwm_setpoint_i20_LC_12_30_7 (
            .in0(N__47065),
            .in1(_gnd_net_),
            .in2(N__55714),
            .in3(N__43897),
            .lcout(pwm_setpoint_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56078),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i2_3_lut_LC_12_31_0 .C_ON=1'b0;
    defparam \PWM.i2_3_lut_LC_12_31_0 .SEQ_MODE=4'b0000;
    defparam \PWM.i2_3_lut_LC_12_31_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \PWM.i2_3_lut_LC_12_31_0  (
            .in0(N__41191),
            .in1(N__41170),
            .in2(_gnd_net_),
            .in3(N__47031),
            .lcout(),
            .ltout(\PWM.n13596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i1_4_lut_LC_12_31_1 .C_ON=1'b0;
    defparam \PWM.i1_4_lut_LC_12_31_1 .SEQ_MODE=4'b0000;
    defparam \PWM.i1_4_lut_LC_12_31_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \PWM.i1_4_lut_LC_12_31_1  (
            .in0(N__41400),
            .in1(N__41342),
            .in2(N__41536),
            .in3(N__41532),
            .lcout(),
            .ltout(\PWM.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i13_4_lut_LC_12_31_2 .C_ON=1'b0;
    defparam \PWM.i13_4_lut_LC_12_31_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i13_4_lut_LC_12_31_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i13_4_lut_LC_12_31_2  (
            .in0(N__41512),
            .in1(N__41496),
            .in2(N__41479),
            .in3(N__41711),
            .lcout(),
            .ltout(\PWM.n29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i9623_4_lut_LC_12_31_3 .C_ON=1'b0;
    defparam \PWM.i9623_4_lut_LC_12_31_3 .SEQ_MODE=4'b0000;
    defparam \PWM.i9623_4_lut_LC_12_31_3 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \PWM.i9623_4_lut_LC_12_31_3  (
            .in0(N__41474),
            .in1(N__44041),
            .in2(N__41455),
            .in3(N__41452),
            .lcout(\PWM.pwm_counter_31__N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i15_2_lut_LC_12_31_4.C_ON=1'b0;
    defparam LessThan_275_i15_2_lut_LC_12_31_4.SEQ_MODE=4'b0000;
    defparam LessThan_275_i15_2_lut_LC_12_31_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i15_2_lut_LC_12_31_4 (
            .in0(_gnd_net_),
            .in1(N__47030),
            .in2(_gnd_net_),
            .in3(N__46927),
            .lcout(n15_adj_613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i39_2_lut_LC_12_31_6.C_ON=1'b0;
    defparam LessThan_275_i39_2_lut_LC_12_31_6.SEQ_MODE=4'b0000;
    defparam LessThan_275_i39_2_lut_LC_12_31_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i39_2_lut_LC_12_31_6 (
            .in0(_gnd_net_),
            .in1(N__41373),
            .in2(_gnd_net_),
            .in3(N__41399),
            .lcout(n39),
            .ltout(n39_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12411_3_lut_LC_12_31_7.C_ON=1'b0;
    defparam i12411_3_lut_LC_12_31_7.SEQ_MODE=4'b0000;
    defparam i12411_3_lut_LC_12_31_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12411_3_lut_LC_12_31_7 (
            .in0(N__41374),
            .in1(_gnd_net_),
            .in2(N__41365),
            .in3(N__43963),
            .lcout(n14883),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i19_2_lut_LC_12_32_1.C_ON=1'b0;
    defparam LessThan_275_i19_2_lut_LC_12_32_1.SEQ_MODE=4'b0000;
    defparam LessThan_275_i19_2_lut_LC_12_32_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i19_2_lut_LC_12_32_1 (
            .in0(_gnd_net_),
            .in1(N__52763),
            .in2(_gnd_net_),
            .in3(N__41343),
            .lcout(n19_adj_616),
            .ltout(n19_adj_616_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12328_4_lut_LC_12_32_2.C_ON=1'b0;
    defparam i12328_4_lut_LC_12_32_2.SEQ_MODE=4'b0000;
    defparam i12328_4_lut_LC_12_32_2.LUT_INIT=16'b1111110011111101;
    LogicCell40 i12328_4_lut_LC_12_32_2 (
            .in0(N__41317),
            .in1(N__41799),
            .in2(N__41308),
            .in3(N__41305),
            .lcout(),
            .ltout(n14800_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12398_4_lut_LC_12_32_3.C_ON=1'b0;
    defparam i12398_4_lut_LC_12_32_3.SEQ_MODE=4'b0000;
    defparam i12398_4_lut_LC_12_32_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12398_4_lut_LC_12_32_3 (
            .in0(N__41763),
            .in1(N__41832),
            .in2(N__41809),
            .in3(N__41685),
            .lcout(n14870),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12262_4_lut_LC_12_32_4.C_ON=1'b0;
    defparam i12262_4_lut_LC_12_32_4.SEQ_MODE=4'b0000;
    defparam i12262_4_lut_LC_12_32_4.LUT_INIT=16'b1111111100000001;
    LogicCell40 i12262_4_lut_LC_12_32_4 (
            .in0(N__41806),
            .in1(N__41800),
            .in2(N__41785),
            .in3(N__41764),
            .lcout(n14734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12402_4_lut_LC_12_32_6.C_ON=1'b0;
    defparam i12402_4_lut_LC_12_32_6.SEQ_MODE=4'b0000;
    defparam i12402_4_lut_LC_12_32_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12402_4_lut_LC_12_32_6 (
            .in0(N__43981),
            .in1(N__43924),
            .in2(N__46891),
            .in3(N__46804),
            .lcout(n14874),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i25_2_lut_LC_12_32_7.C_ON=1'b0;
    defparam LessThan_275_i25_2_lut_LC_12_32_7.SEQ_MODE=4'b0000;
    defparam LessThan_275_i25_2_lut_LC_12_32_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_275_i25_2_lut_LC_12_32_7 (
            .in0(N__41727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41713),
            .lcout(n25_adj_620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12347_3_lut_LC_13_17_0.C_ON=1'b0;
    defparam i12347_3_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam i12347_3_lut_LC_13_17_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12347_3_lut_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(N__41674),
            .in2(N__41650),
            .in3(N__47568),
            .lcout(n2822),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_13_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_13_17_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1856_3_lut_LC_13_17_1 (
            .in0(N__41637),
            .in1(_gnd_net_),
            .in2(N__47605),
            .in3(N__41617),
            .lcout(n2824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_55_LC_13_17_2.C_ON=1'b0;
    defparam i1_4_lut_adj_55_LC_13_17_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_55_LC_13_17_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_55_LC_13_17_2 (
            .in0(N__44165),
            .in1(N__41611),
            .in2(N__44116),
            .in3(N__41602),
            .lcout(),
            .ltout(n14054_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_56_LC_13_17_3.C_ON=1'b0;
    defparam i1_4_lut_adj_56_LC_13_17_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_56_LC_13_17_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_56_LC_13_17_3 (
            .in0(N__42231),
            .in1(N__41593),
            .in2(N__41575),
            .in3(N__44246),
            .lcout(),
            .ltout(n14060_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13000_4_lut_LC_13_17_4.C_ON=1'b0;
    defparam i13000_4_lut_LC_13_17_4.SEQ_MODE=4'b0000;
    defparam i13000_4_lut_LC_13_17_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13000_4_lut_LC_13_17_4 (
            .in0(N__42305),
            .in1(N__41568),
            .in2(N__41539),
            .in3(N__42027),
            .lcout(n2742),
            .ltout(n2742_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_13_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_13_17_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1862_3_lut_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(N__41998),
            .in2(N__41992),
            .in3(N__41989),
            .lcout(n2830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_13_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_13_17_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1859_3_lut_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__41961),
            .in2(N__41938),
            .in3(N__47567),
            .lcout(n2827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_44_LC_13_18_0.C_ON=1'b0;
    defparam i1_4_lut_adj_44_LC_13_18_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_44_LC_13_18_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_44_LC_13_18_0 (
            .in0(N__47762),
            .in1(N__48128),
            .in2(N__48224),
            .in3(N__47726),
            .lcout(),
            .ltout(n14238_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_45_LC_13_18_1.C_ON=1'b0;
    defparam i1_3_lut_adj_45_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_45_LC_13_18_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_45_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__48176),
            .in2(N__41929),
            .in3(N__48303),
            .lcout(),
            .ltout(n14240_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_46_LC_13_18_2.C_ON=1'b0;
    defparam i1_4_lut_adj_46_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_46_LC_13_18_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_46_LC_13_18_2 (
            .in0(N__48038),
            .in1(N__47999),
            .in2(N__41926),
            .in3(N__48080),
            .lcout(n14246),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_13_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_13_18_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1851_3_lut_LC_13_18_3 (
            .in0(N__47577),
            .in1(_gnd_net_),
            .in2(N__41923),
            .in3(N__41905),
            .lcout(n2819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_13_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_13_18_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1853_3_lut_LC_13_18_4 (
            .in0(N__41896),
            .in1(_gnd_net_),
            .in2(N__41890),
            .in3(N__47572),
            .lcout(n2821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_13_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_13_18_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1861_3_lut_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__41863),
            .in2(N__47606),
            .in3(N__41857),
            .lcout(n2829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12349_3_lut_LC_13_18_6.C_ON=1'b0;
    defparam i12349_3_lut_LC_13_18_6.SEQ_MODE=4'b0000;
    defparam i12349_3_lut_LC_13_18_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12349_3_lut_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(N__42183),
            .in2(N__42160),
            .in3(N__47573),
            .lcout(n2823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_13_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_13_18_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1850_3_lut_LC_13_18_7 (
            .in0(_gnd_net_),
            .in1(N__42148),
            .in2(N__47607),
            .in3(N__42142),
            .lcout(n2818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_13_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_13_19_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1921_3_lut_LC_13_19_0 (
            .in0(N__48186),
            .in1(_gnd_net_),
            .in2(N__48160),
            .in3(N__49312),
            .lcout(n2921),
            .ltout(n2921_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_36_LC_13_19_1.C_ON=1'b0;
    defparam i1_2_lut_adj_36_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_36_LC_13_19_1.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_36_LC_13_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42100),
            .in3(N__44528),
            .lcout(n13926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_13_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_13_19_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1915_3_lut_LC_13_19_2 (
            .in0(_gnd_net_),
            .in1(N__48553),
            .in2(N__48523),
            .in3(N__49316),
            .lcout(n2915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_13_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_13_19_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1918_3_lut_LC_13_19_3 (
            .in0(_gnd_net_),
            .in1(N__48042),
            .in2(N__49353),
            .in3(N__48022),
            .lcout(n2918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_13_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_13_19_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1842_3_lut_LC_13_19_4 (
            .in0(_gnd_net_),
            .in1(N__42097),
            .in2(N__42310),
            .in3(N__47594),
            .lcout(n2810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_13_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_13_19_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1917_3_lut_LC_13_19_5 (
            .in0(_gnd_net_),
            .in1(N__48604),
            .in2(N__49354),
            .in3(N__48003),
            .lcout(n2917),
            .ltout(n2917_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_38_LC_13_19_6.C_ON=1'b0;
    defparam i1_4_lut_adj_38_LC_13_19_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_38_LC_13_19_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_38_LC_13_19_6 (
            .in0(N__42053),
            .in1(N__42037),
            .in2(N__42031),
            .in3(N__44456),
            .lcout(),
            .ltout(n13934_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_39_LC_13_19_7.C_ON=1'b0;
    defparam i1_4_lut_adj_39_LC_13_19_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_39_LC_13_19_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_39_LC_13_19_7 (
            .in0(N__42548),
            .in1(N__42524),
            .in2(N__42508),
            .in3(N__44704),
            .lcout(n13942),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_13_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_13_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_13_20_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1775_3_lut_LC_13_20_0 (
            .in0(_gnd_net_),
            .in1(N__42496),
            .in2(N__42484),
            .in3(N__42444),
            .lcout(n2711),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12995_1_lut_LC_13_20_1.C_ON=1'b0;
    defparam i12995_1_lut_LC_13_20_1.SEQ_MODE=4'b0000;
    defparam i12995_1_lut_LC_13_20_1.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12995_1_lut_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47625),
            .in3(_gnd_net_),
            .lcout(n15467),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_13_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_13_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_13_20_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1909_3_lut_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(N__49336),
            .in2(N__48906),
            .in3(N__48880),
            .lcout(n2909),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_13_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_13_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_13_20_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2119_3_lut_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(N__51730),
            .in2(N__50118),
            .in3(N__51749),
            .lcout(n3215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_13_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_13_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_13_20_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2122_3_lut_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(N__51222),
            .in2(N__51199),
            .in3(N__50109),
            .lcout(n3218),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_13_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_13_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_13_20_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1844_3_lut_LC_13_20_7 (
            .in0(_gnd_net_),
            .in1(N__42232),
            .in2(N__47626),
            .in3(N__42202),
            .lcout(n2812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_29_LC_13_21_0.C_ON=1'b0;
    defparam i1_4_lut_adj_29_LC_13_21_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_29_LC_13_21_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_29_LC_13_21_0 (
            .in0(N__45491),
            .in1(N__45146),
            .in2(N__45456),
            .in3(N__45113),
            .lcout(),
            .ltout(n14322_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_30_LC_13_21_1.C_ON=1'b0;
    defparam i1_4_lut_adj_30_LC_13_21_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_30_LC_13_21_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_30_LC_13_21_1 (
            .in0(N__45423),
            .in1(N__45378),
            .in2(N__42196),
            .in3(N__42637),
            .lcout(n14328),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_13_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_13_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_13_21_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1992_3_lut_LC_13_21_2 (
            .in0(N__42664),
            .in1(N__44943),
            .in2(_gnd_net_),
            .in3(N__42946),
            .lcout(n3024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_13_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_13_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_13_21_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1991_3_lut_LC_13_21_3 (
            .in0(N__44460),
            .in1(_gnd_net_),
            .in2(N__42994),
            .in3(N__42652),
            .lcout(n3023),
            .ltout(n3023_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_28_LC_13_21_4.C_ON=1'b0;
    defparam i1_4_lut_adj_28_LC_13_21_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_28_LC_13_21_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_28_LC_13_21_4 (
            .in0(N__45044),
            .in1(N__45008),
            .in2(N__42640),
            .in3(N__45083),
            .lcout(n14320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_13_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_13_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_13_21_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1995_3_lut_LC_13_21_5 (
            .in0(_gnd_net_),
            .in1(N__42631),
            .in2(N__42995),
            .in3(N__44571),
            .lcout(n3027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_13_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_13_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_13_21_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1994_3_lut_LC_13_21_6 (
            .in0(_gnd_net_),
            .in1(N__44625),
            .in2(N__42622),
            .in3(N__42945),
            .lcout(n3026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_13_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_13_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_13_22_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1913_3_lut_LC_13_22_0 (
            .in0(_gnd_net_),
            .in1(N__48442),
            .in2(N__48469),
            .in3(N__49359),
            .lcout(n2913),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_13_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_13_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_13_22_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2061_3_lut_LC_13_22_1 (
            .in0(_gnd_net_),
            .in1(N__45067),
            .in2(N__49041),
            .in3(N__45087),
            .lcout(n3125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_13_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_13_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_13_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1990_3_lut_LC_13_22_2 (
            .in0(_gnd_net_),
            .in1(N__42583),
            .in2(N__44308),
            .in3(N__42961),
            .lcout(n3022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_13_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_13_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_13_22_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1982_3_lut_LC_13_22_3 (
            .in0(N__42963),
            .in1(_gnd_net_),
            .in2(N__42574),
            .in3(N__42558),
            .lcout(n3014),
            .ltout(n3014_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_13_22_4.C_ON=1'b0;
    defparam i1_3_lut_LC_13_22_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_13_22_4.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_LC_13_22_4 (
            .in0(N__45345),
            .in1(_gnd_net_),
            .in2(N__43018),
            .in3(N__45269),
            .lcout(n14408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_13_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_13_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_13_22_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1989_3_lut_LC_13_22_5 (
            .in0(N__42962),
            .in1(N__42862),
            .in2(N__44544),
            .in3(_gnd_net_),
            .lcout(n3021),
            .ltout(n3021_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_13_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_13_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_13_22_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2056_3_lut_LC_13_22_6 (
            .in0(_gnd_net_),
            .in1(N__45439),
            .in2(N__42853),
            .in3(N__48988),
            .lcout(n3120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_13_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_13_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_13_22_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2066_3_lut_LC_13_22_7 (
            .in0(_gnd_net_),
            .in1(N__44716),
            .in2(N__49042),
            .in3(N__44742),
            .lcout(n3130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_2_LC_13_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_2_LC_13_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_2_LC_13_23_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 encoder0_position_31__I_0_add_2173_2_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(N__42850),
            .in2(N__54865),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(n12521),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_13_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_13_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_13_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_3_lut_LC_13_23_1 (
            .in0(_gnd_net_),
            .in1(N__42823),
            .in2(_gnd_net_),
            .in3(N__42772),
            .lcout(n3301),
            .ltout(),
            .carryin(n12521),
            .carryout(n12522),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_13_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_13_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_13_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_4_lut_LC_13_23_2 (
            .in0(_gnd_net_),
            .in1(N__42769),
            .in2(N__54866),
            .in3(N__42730),
            .lcout(n3300),
            .ltout(),
            .carryin(n12522),
            .carryout(n12523),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_13_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_13_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_13_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_5_lut_LC_13_23_3 (
            .in0(_gnd_net_),
            .in1(N__42723),
            .in2(_gnd_net_),
            .in3(N__42694),
            .lcout(n3299),
            .ltout(),
            .carryin(n12523),
            .carryout(n12524),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_13_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_13_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_13_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_6_lut_LC_13_23_4 (
            .in0(_gnd_net_),
            .in1(N__42691),
            .in2(N__54867),
            .in3(N__42667),
            .lcout(n3298),
            .ltout(),
            .carryin(n12524),
            .carryout(n12525),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_13_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_13_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_13_23_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 encoder0_position_31__I_0_add_2173_7_lut_LC_13_23_5 (
            .in0(N__43111),
            .in1(_gnd_net_),
            .in2(N__43105),
            .in3(N__43066),
            .lcout(n14697),
            .ltout(),
            .carryin(n12525),
            .carryout(n12526),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_13_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_13_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_13_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_8_lut_LC_13_23_6 (
            .in0(_gnd_net_),
            .in1(N__48682),
            .in2(_gnd_net_),
            .in3(N__43063),
            .lcout(n3296),
            .ltout(),
            .carryin(n12526),
            .carryout(n12527),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_13_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_13_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_13_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_9_lut_LC_13_23_7 (
            .in0(_gnd_net_),
            .in1(N__54403),
            .in2(N__45787),
            .in3(N__43060),
            .lcout(n3295),
            .ltout(),
            .carryin(n12527),
            .carryout(n12528),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_13_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_13_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_13_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_10_lut_LC_13_24_0 (
            .in0(_gnd_net_),
            .in1(N__46107),
            .in2(N__54868),
            .in3(N__43057),
            .lcout(n3294),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(n12529),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_13_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_13_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_13_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_11_lut_LC_13_24_1 (
            .in0(_gnd_net_),
            .in1(N__49398),
            .in2(N__54872),
            .in3(N__43048),
            .lcout(n3293),
            .ltout(),
            .carryin(n12529),
            .carryout(n12530),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_13_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_13_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_13_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_12_lut_LC_13_24_2 (
            .in0(_gnd_net_),
            .in1(N__49656),
            .in2(N__54869),
            .in3(N__43045),
            .lcout(n3292),
            .ltout(),
            .carryin(n12530),
            .carryout(n12531),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_13_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_13_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_13_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_13_lut_LC_13_24_3 (
            .in0(_gnd_net_),
            .in1(N__45765),
            .in2(N__54873),
            .in3(N__43033),
            .lcout(n3291),
            .ltout(),
            .carryin(n12531),
            .carryout(n12532),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_13_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_13_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_13_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_14_lut_LC_13_24_4 (
            .in0(_gnd_net_),
            .in1(N__46133),
            .in2(N__54870),
            .in3(N__43021),
            .lcout(n3290),
            .ltout(),
            .carryin(n12532),
            .carryout(n12533),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_13_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_13_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_13_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_15_lut_LC_13_24_5 (
            .in0(_gnd_net_),
            .in1(N__48635),
            .in2(N__54874),
            .in3(N__43267),
            .lcout(n3289),
            .ltout(),
            .carryin(n12533),
            .carryout(n12534),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_13_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_13_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_13_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_16_lut_LC_13_24_6 (
            .in0(_gnd_net_),
            .in1(N__45870),
            .in2(N__54871),
            .in3(N__43258),
            .lcout(n3288),
            .ltout(),
            .carryin(n12534),
            .carryout(n12535),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_13_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_13_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_13_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_17_lut_LC_13_24_7 (
            .in0(_gnd_net_),
            .in1(N__48734),
            .in2(N__54875),
            .in3(N__43255),
            .lcout(n3287),
            .ltout(),
            .carryin(n12535),
            .carryout(n12536),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_13_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_13_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_13_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_18_lut_LC_13_25_0 (
            .in0(_gnd_net_),
            .in1(N__49689),
            .in2(N__54876),
            .in3(N__43252),
            .lcout(n3286),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(n12537),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_13_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_13_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_13_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_19_lut_LC_13_25_1 (
            .in0(_gnd_net_),
            .in1(N__54431),
            .in2(N__45838),
            .in3(N__43243),
            .lcout(n3285),
            .ltout(),
            .carryin(n12537),
            .carryout(n12538),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_13_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_13_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_13_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_20_lut_LC_13_25_2 (
            .in0(_gnd_net_),
            .in1(N__43236),
            .in2(N__54877),
            .in3(N__43210),
            .lcout(n3284),
            .ltout(),
            .carryin(n12538),
            .carryout(n12539),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_13_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_13_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_13_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_21_lut_LC_13_25_3 (
            .in0(_gnd_net_),
            .in1(N__43207),
            .in2(N__54880),
            .in3(N__43174),
            .lcout(n3283),
            .ltout(),
            .carryin(n12539),
            .carryout(n12540),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_13_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_13_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_13_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_22_lut_LC_13_25_4 (
            .in0(_gnd_net_),
            .in1(N__43166),
            .in2(N__54878),
            .in3(N__43135),
            .lcout(n3282),
            .ltout(),
            .carryin(n12540),
            .carryout(n12541),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_13_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_13_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_13_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_23_lut_LC_13_25_5 (
            .in0(_gnd_net_),
            .in1(N__43130),
            .in2(N__54881),
            .in3(N__43495),
            .lcout(n3281),
            .ltout(),
            .carryin(n12541),
            .carryout(n12542),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_13_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_13_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_13_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_24_lut_LC_13_25_6 (
            .in0(_gnd_net_),
            .in1(N__49928),
            .in2(N__54879),
            .in3(N__43486),
            .lcout(n3280),
            .ltout(),
            .carryin(n12542),
            .carryout(n12543),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_13_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_13_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_13_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_25_lut_LC_13_25_7 (
            .in0(_gnd_net_),
            .in1(N__43483),
            .in2(N__54882),
            .in3(N__43444),
            .lcout(n3279),
            .ltout(),
            .carryin(n12543),
            .carryout(n12544),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_13_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_13_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_13_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_26_lut_LC_13_26_0 (
            .in0(_gnd_net_),
            .in1(N__43440),
            .in2(N__54883),
            .in3(N__43405),
            .lcout(n3278),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(n12545),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_13_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_13_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_13_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_27_lut_LC_13_26_1 (
            .in0(_gnd_net_),
            .in1(N__43402),
            .in2(N__54887),
            .in3(N__43363),
            .lcout(n3277),
            .ltout(),
            .carryin(n12545),
            .carryout(n12546),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_13_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_13_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_13_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_28_lut_LC_13_26_2 (
            .in0(_gnd_net_),
            .in1(N__49427),
            .in2(N__54884),
            .in3(N__43348),
            .lcout(n3276),
            .ltout(),
            .carryin(n12546),
            .carryout(n12547),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_13_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_13_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_13_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_29_lut_LC_13_26_3 (
            .in0(_gnd_net_),
            .in1(N__43345),
            .in2(N__54888),
            .in3(N__43309),
            .lcout(n3275),
            .ltout(),
            .carryin(n12547),
            .carryout(n12548),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_13_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_13_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_13_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_30_lut_LC_13_26_4 (
            .in0(_gnd_net_),
            .in1(N__43306),
            .in2(N__54885),
            .in3(N__43270),
            .lcout(n3274),
            .ltout(),
            .carryin(n12548),
            .carryout(n12549),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_13_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_13_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_13_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_31_lut_LC_13_26_5 (
            .in0(_gnd_net_),
            .in1(N__43672),
            .in2(N__54889),
            .in3(N__43630),
            .lcout(n3273),
            .ltout(),
            .carryin(n12549),
            .carryout(n12550),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_13_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_13_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_13_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_32_lut_LC_13_26_6 (
            .in0(_gnd_net_),
            .in1(N__43627),
            .in2(N__54886),
            .in3(N__43594),
            .lcout(n3272),
            .ltout(),
            .carryin(n12550),
            .carryout(n12551),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_13_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_13_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_13_26_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_2173_33_lut_LC_13_26_7 (
            .in0(N__54471),
            .in1(N__43591),
            .in2(N__51910),
            .in3(N__43573),
            .lcout(n14461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i7_1_lut_LC_13_27_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_13_27_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_13_27_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i7_1_lut_LC_13_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46314),
            .lcout(n19_adj_585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 unary_minus_13_inv_0_i3_1_lut_LC_13_27_1 (
            .in0(N__46041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n23_adj_589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i11_1_lut_LC_13_27_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_13_27_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_13_27_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i11_1_lut_LC_13_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46227),
            .lcout(n15_adj_581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i6_1_lut_LC_13_27_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_13_27_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_13_27_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i6_1_lut_LC_13_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45954),
            .lcout(n20_adj_586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i4_1_lut_LC_13_27_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i4_1_lut_LC_13_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i4_1_lut_LC_13_27_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i4_1_lut_LC_13_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43558),
            .lcout(n22_adj_548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_13_27_5.C_ON=1'b0;
    defparam i2_2_lut_LC_13_27_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_13_27_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_LC_13_27_5 (
            .in0(_gnd_net_),
            .in1(N__43544),
            .in2(_gnd_net_),
            .in3(N__43523),
            .lcout(n10_adj_680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i1_1_lut_LC_13_27_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_13_27_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_13_27_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i1_1_lut_LC_13_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46473),
            .lcout(n25_adj_591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i15_1_lut_LC_13_27_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_13_27_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_13_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i15_1_lut_LC_13_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46560),
            .lcout(n11_adj_577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_2_lut_LC_13_28_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_2_lut_LC_13_28_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_2_lut_LC_13_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_2_lut_LC_13_28_0 (
            .in0(_gnd_net_),
            .in1(N__43762),
            .in2(_gnd_net_),
            .in3(N__43756),
            .lcout(pwm_setpoint_23_N_171_0),
            .ltout(),
            .carryin(bfn_13_28_0_),
            .carryout(n12050),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_3_lut_LC_13_28_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_3_lut_LC_13_28_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_3_lut_LC_13_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_3_lut_LC_13_28_1 (
            .in0(_gnd_net_),
            .in1(N__50206),
            .in2(_gnd_net_),
            .in3(N__43753),
            .lcout(pwm_setpoint_23_N_171_1),
            .ltout(),
            .carryin(n12050),
            .carryout(n12051),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_4_lut_LC_13_28_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_4_lut_LC_13_28_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_4_lut_LC_13_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_4_lut_LC_13_28_2 (
            .in0(_gnd_net_),
            .in1(N__43750),
            .in2(_gnd_net_),
            .in3(N__43738),
            .lcout(pwm_setpoint_23_N_171_2),
            .ltout(),
            .carryin(n12051),
            .carryout(n12052),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_5_lut_LC_13_28_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_5_lut_LC_13_28_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_5_lut_LC_13_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_5_lut_LC_13_28_3 (
            .in0(_gnd_net_),
            .in1(N__50173),
            .in2(_gnd_net_),
            .in3(N__43729),
            .lcout(pwm_setpoint_23_N_171_3),
            .ltout(),
            .carryin(n12052),
            .carryout(n12053),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_6_lut_LC_13_28_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_6_lut_LC_13_28_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_6_lut_LC_13_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_6_lut_LC_13_28_4 (
            .in0(_gnd_net_),
            .in1(N__43726),
            .in2(_gnd_net_),
            .in3(N__43708),
            .lcout(pwm_setpoint_23_N_171_4),
            .ltout(),
            .carryin(n12053),
            .carryout(n12054),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_7_lut_LC_13_28_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_7_lut_LC_13_28_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_7_lut_LC_13_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_7_lut_LC_13_28_5 (
            .in0(_gnd_net_),
            .in1(N__43705),
            .in2(_gnd_net_),
            .in3(N__43690),
            .lcout(pwm_setpoint_23_N_171_5),
            .ltout(),
            .carryin(n12054),
            .carryout(n12055),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_8_lut_LC_13_28_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_8_lut_LC_13_28_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_8_lut_LC_13_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_8_lut_LC_13_28_6 (
            .in0(_gnd_net_),
            .in1(N__43687),
            .in2(_gnd_net_),
            .in3(N__43675),
            .lcout(pwm_setpoint_23_N_171_6),
            .ltout(),
            .carryin(n12055),
            .carryout(n12056),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_9_lut_LC_13_28_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_9_lut_LC_13_28_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_9_lut_LC_13_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_9_lut_LC_13_28_7 (
            .in0(_gnd_net_),
            .in1(N__43846),
            .in2(_gnd_net_),
            .in3(N__43840),
            .lcout(pwm_setpoint_23_N_171_7),
            .ltout(),
            .carryin(n12056),
            .carryout(n12057),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_10_lut_LC_13_29_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_10_lut_LC_13_29_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_10_lut_LC_13_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_10_lut_LC_13_29_0 (
            .in0(_gnd_net_),
            .in1(N__52711),
            .in2(_gnd_net_),
            .in3(N__43831),
            .lcout(pwm_setpoint_23_N_171_8),
            .ltout(),
            .carryin(bfn_13_29_0_),
            .carryout(n12058),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_11_lut_LC_13_29_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_11_lut_LC_13_29_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_11_lut_LC_13_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_11_lut_LC_13_29_1 (
            .in0(_gnd_net_),
            .in1(N__46510),
            .in2(_gnd_net_),
            .in3(N__43828),
            .lcout(pwm_setpoint_23_N_171_9),
            .ltout(),
            .carryin(n12058),
            .carryout(n12059),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_12_lut_LC_13_29_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_12_lut_LC_13_29_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_12_lut_LC_13_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_12_lut_LC_13_29_2 (
            .in0(_gnd_net_),
            .in1(N__43825),
            .in2(_gnd_net_),
            .in3(N__43810),
            .lcout(pwm_setpoint_23_N_171_10),
            .ltout(),
            .carryin(n12059),
            .carryout(n12060),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_13_lut_LC_13_29_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_13_lut_LC_13_29_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_13_lut_LC_13_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_13_lut_LC_13_29_3 (
            .in0(_gnd_net_),
            .in1(N__43807),
            .in2(_gnd_net_),
            .in3(N__43792),
            .lcout(pwm_setpoint_23_N_171_11),
            .ltout(),
            .carryin(n12060),
            .carryout(n12061),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_14_lut_LC_13_29_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_14_lut_LC_13_29_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_14_lut_LC_13_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_14_lut_LC_13_29_4 (
            .in0(_gnd_net_),
            .in1(N__46774),
            .in2(_gnd_net_),
            .in3(N__43780),
            .lcout(pwm_setpoint_23_N_171_12),
            .ltout(),
            .carryin(n12061),
            .carryout(n12062),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_15_lut_LC_13_29_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_15_lut_LC_13_29_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_15_lut_LC_13_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_15_lut_LC_13_29_5 (
            .in0(_gnd_net_),
            .in1(N__46489),
            .in2(_gnd_net_),
            .in3(N__43777),
            .lcout(pwm_setpoint_23_N_171_13),
            .ltout(),
            .carryin(n12062),
            .carryout(n12063),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_16_lut_LC_13_29_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_16_lut_LC_13_29_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_16_lut_LC_13_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_16_lut_LC_13_29_6 (
            .in0(_gnd_net_),
            .in1(N__43774),
            .in2(_gnd_net_),
            .in3(N__43765),
            .lcout(pwm_setpoint_23_N_171_14),
            .ltout(),
            .carryin(n12063),
            .carryout(n12064),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_17_lut_LC_13_29_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_17_lut_LC_13_29_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_17_lut_LC_13_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_17_lut_LC_13_29_7 (
            .in0(_gnd_net_),
            .in1(N__46570),
            .in2(_gnd_net_),
            .in3(N__43918),
            .lcout(pwm_setpoint_23_N_171_15),
            .ltout(),
            .carryin(n12064),
            .carryout(n12065),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_18_lut_LC_13_30_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_18_lut_LC_13_30_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_18_lut_LC_13_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_18_lut_LC_13_30_0 (
            .in0(_gnd_net_),
            .in1(N__46645),
            .in2(_gnd_net_),
            .in3(N__43915),
            .lcout(pwm_setpoint_23_N_171_16),
            .ltout(),
            .carryin(bfn_13_30_0_),
            .carryout(n12066),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_19_lut_LC_13_30_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_19_lut_LC_13_30_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_19_lut_LC_13_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_19_lut_LC_13_30_1 (
            .in0(_gnd_net_),
            .in1(N__47134),
            .in2(_gnd_net_),
            .in3(N__43912),
            .lcout(pwm_setpoint_23_N_171_17),
            .ltout(),
            .carryin(n12066),
            .carryout(n12067),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_20_lut_LC_13_30_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_20_lut_LC_13_30_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_20_lut_LC_13_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_20_lut_LC_13_30_2 (
            .in0(_gnd_net_),
            .in1(N__50233),
            .in2(_gnd_net_),
            .in3(N__43909),
            .lcout(pwm_setpoint_23_N_171_18),
            .ltout(),
            .carryin(n12067),
            .carryout(n12068),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_21_lut_LC_13_30_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_21_lut_LC_13_30_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_21_lut_LC_13_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_21_lut_LC_13_30_3 (
            .in0(_gnd_net_),
            .in1(N__50260),
            .in2(_gnd_net_),
            .in3(N__43900),
            .lcout(pwm_setpoint_23_N_171_19),
            .ltout(),
            .carryin(n12068),
            .carryout(n12069),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_22_lut_LC_13_30_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_22_lut_LC_13_30_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_22_lut_LC_13_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_22_lut_LC_13_30_4 (
            .in0(_gnd_net_),
            .in1(N__47044),
            .in2(_gnd_net_),
            .in3(N__43891),
            .lcout(pwm_setpoint_23_N_171_20),
            .ltout(),
            .carryin(n12069),
            .carryout(n12070),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_23_lut_LC_13_30_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_23_lut_LC_13_30_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_23_lut_LC_13_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_23_lut_LC_13_30_5 (
            .in0(_gnd_net_),
            .in1(N__43888),
            .in2(_gnd_net_),
            .in3(N__43864),
            .lcout(pwm_setpoint_23_N_171_21),
            .ltout(),
            .carryin(n12070),
            .carryout(n12071),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_24_lut_LC_13_30_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_24_lut_LC_13_30_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_24_lut_LC_13_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_24_lut_LC_13_30_6 (
            .in0(_gnd_net_),
            .in1(N__46651),
            .in2(_gnd_net_),
            .in3(N__43861),
            .lcout(pwm_setpoint_23_N_171_22),
            .ltout(),
            .carryin(n12071),
            .carryout(n12072),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i23_LC_13_30_7.C_ON=1'b0;
    defparam pwm_setpoint_i23_LC_13_30_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i23_LC_13_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 pwm_setpoint_i23_LC_13_30_7 (
            .in0(_gnd_net_),
            .in1(N__55563),
            .in2(_gnd_net_),
            .in3(N__43858),
            .lcout(pwm_setpoint_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56082),
            .ce(),
            .sr(N__55567));
    defparam pwm_setpoint_i15_LC_13_31_0.C_ON=1'b0;
    defparam pwm_setpoint_i15_LC_13_31_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i15_LC_13_31_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i15_LC_13_31_0 (
            .in0(N__44077),
            .in1(N__55656),
            .in2(_gnd_net_),
            .in3(N__46588),
            .lcout(pwm_setpoint_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i18_LC_13_31_1.C_ON=1'b0;
    defparam pwm_setpoint_i18_LC_13_31_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i18_LC_13_31_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i18_LC_13_31_1 (
            .in0(N__55655),
            .in1(N__50251),
            .in2(_gnd_net_),
            .in3(N__44068),
            .lcout(pwm_setpoint_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i12_4_lut_LC_13_31_2 .C_ON=1'b0;
    defparam \PWM.i12_4_lut_LC_13_31_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i12_4_lut_LC_13_31_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i12_4_lut_LC_13_31_2  (
            .in0(N__44061),
            .in1(N__44274),
            .in2(N__46843),
            .in3(N__46747),
            .lcout(\PWM.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i31_2_lut_LC_13_31_3.C_ON=1'b0;
    defparam LessThan_275_i31_2_lut_LC_13_31_3.SEQ_MODE=4'b0000;
    defparam LessThan_275_i31_2_lut_LC_13_31_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i31_2_lut_LC_13_31_3 (
            .in0(_gnd_net_),
            .in1(N__46980),
            .in2(_gnd_net_),
            .in3(N__44031),
            .lcout(n31_adj_624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i37_2_lut_LC_13_31_4.C_ON=1'b0;
    defparam LessThan_275_i37_2_lut_LC_13_31_4.SEQ_MODE=4'b0000;
    defparam LessThan_275_i37_2_lut_LC_13_31_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i37_2_lut_LC_13_31_4 (
            .in0(_gnd_net_),
            .in1(N__43974),
            .in2(_gnd_net_),
            .in3(N__44000),
            .lcout(n37),
            .ltout(n37_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12415_3_lut_LC_13_31_5.C_ON=1'b0;
    defparam i12415_3_lut_LC_13_31_5.SEQ_MODE=4'b0000;
    defparam i12415_3_lut_LC_13_31_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12415_3_lut_LC_13_31_5 (
            .in0(N__43975),
            .in1(_gnd_net_),
            .in2(N__43966),
            .in3(N__46987),
            .lcout(n14887),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i22_LC_13_31_6.C_ON=1'b0;
    defparam pwm_setpoint_i22_LC_13_31_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i22_LC_13_31_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i22_LC_13_31_6 (
            .in0(N__55709),
            .in1(N__46666),
            .in2(_gnd_net_),
            .in3(N__43957),
            .lcout(pwm_setpoint_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i17_LC_13_32_0.C_ON=1'b0;
    defparam pwm_setpoint_i17_LC_13_32_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i17_LC_13_32_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i17_LC_13_32_0 (
            .in0(N__47152),
            .in1(N__55708),
            .in2(_gnd_net_),
            .in3(N__43939),
            .lcout(pwm_setpoint_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56090),
            .ce(),
            .sr(_gnd_net_));
    defparam i12360_4_lut_LC_13_32_3.C_ON=1'b0;
    defparam i12360_4_lut_LC_13_32_3.SEQ_MODE=4'b0000;
    defparam i12360_4_lut_LC_13_32_3.LUT_INIT=16'b1111111111111101;
    LogicCell40 i12360_4_lut_LC_13_32_3 (
            .in0(N__43930),
            .in1(N__47179),
            .in2(N__46720),
            .in3(N__47212),
            .lcout(n14832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i35_2_lut_LC_13_32_4.C_ON=1'b0;
    defparam LessThan_275_i35_2_lut_LC_13_32_4.SEQ_MODE=4'b0000;
    defparam LessThan_275_i35_2_lut_LC_13_32_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i35_2_lut_LC_13_32_4 (
            .in0(_gnd_net_),
            .in1(N__46905),
            .in2(_gnd_net_),
            .in3(N__44275),
            .lcout(n35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_14_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_14_17_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1843_3_lut_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(N__44251),
            .in2(N__44224),
            .in3(N__47562),
            .lcout(n2811),
            .ltout(n2811_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_48_LC_14_17_1.C_ON=1'b0;
    defparam i1_4_lut_adj_48_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_48_LC_14_17_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_48_LC_14_17_1 (
            .in0(N__48384),
            .in1(N__44083),
            .in2(N__44209),
            .in3(N__48425),
            .lcout(n14266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_14_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_14_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1858_3_lut_LC_14_17_2 (
            .in0(_gnd_net_),
            .in1(N__44206),
            .in2(N__44197),
            .in3(N__47554),
            .lcout(n2826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_14_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_14_17_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1933_3_lut_LC_14_17_3 (
            .in0(N__47227),
            .in1(N__47260),
            .in2(_gnd_net_),
            .in3(N__49273),
            .lcout(n2933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_14_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_14_17_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1847_3_lut_LC_14_17_4 (
            .in0(_gnd_net_),
            .in1(N__44166),
            .in2(N__44143),
            .in3(N__47558),
            .lcout(n2815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_14_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_14_17_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1846_3_lut_LC_14_17_5 (
            .in0(_gnd_net_),
            .in1(N__44128),
            .in2(N__47603),
            .in3(N__44115),
            .lcout(n2814),
            .ltout(n2814_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_43_LC_14_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_43_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_43_LC_14_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_43_LC_14_17_6 (
            .in0(N__47810),
            .in1(N__48263),
            .in2(N__44086),
            .in3(N__48494),
            .lcout(n14260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_14_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_14_17_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1860_3_lut_LC_14_17_7 (
            .in0(N__44440),
            .in1(_gnd_net_),
            .in2(N__47602),
            .in3(N__44431),
            .lcout(n2828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_14_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_14_18_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1864_3_lut_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(N__44404),
            .in2(N__44392),
            .in3(N__47563),
            .lcout(n2832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_14_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_14_18_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1863_3_lut_LC_14_18_1 (
            .in0(_gnd_net_),
            .in1(N__44362),
            .in2(N__47604),
            .in3(N__44350),
            .lcout(n2831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_14_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_14_18_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1929_3_lut_LC_14_18_2 (
            .in0(N__47866),
            .in1(_gnd_net_),
            .in2(N__47889),
            .in3(N__49320),
            .lcout(n2929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_47_LC_14_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_47_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_47_LC_14_18_3.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_47_LC_14_18_3 (
            .in0(N__47470),
            .in1(N__47882),
            .in2(N__47850),
            .in3(N__44329),
            .lcout(),
            .ltout(n14248_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_49_LC_14_18_4.C_ON=1'b0;
    defparam i1_4_lut_adj_49_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_49_LC_14_18_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_49_LC_14_18_4 (
            .in0(N__48545),
            .in1(N__48585),
            .in2(N__44323),
            .in3(N__48864),
            .lcout(),
            .ltout(n14254_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12452_4_lut_LC_14_18_5.C_ON=1'b0;
    defparam i12452_4_lut_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam i12452_4_lut_LC_14_18_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12452_4_lut_LC_14_18_5 (
            .in0(N__48800),
            .in1(N__48896),
            .in2(N__44320),
            .in3(N__44317),
            .lcout(n2841),
            .ltout(n2841_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_14_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_14_18_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1923_3_lut_LC_14_18_6 (
            .in0(N__48247),
            .in1(_gnd_net_),
            .in2(N__44311),
            .in3(N__48273),
            .lcout(n2923),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_35_LC_14_19_0.C_ON=1'b0;
    defparam i1_4_lut_adj_35_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_35_LC_14_19_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_35_LC_14_19_0 (
            .in0(N__44556),
            .in1(N__44286),
            .in2(N__44654),
            .in3(N__44939),
            .lcout(),
            .ltout(n13932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_37_LC_14_19_1.C_ON=1'b0;
    defparam i1_4_lut_adj_37_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_37_LC_14_19_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_37_LC_14_19_1 (
            .in0(N__44615),
            .in1(N__44684),
            .in2(N__44707),
            .in3(N__44588),
            .lcout(n13936),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_14_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_14_19_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1926_3_lut_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(N__47746),
            .in2(N__47782),
            .in3(N__49296),
            .lcout(n2926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_14_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_14_19_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1920_3_lut_LC_14_19_3 (
            .in0(N__49293),
            .in1(_gnd_net_),
            .in2(N__48138),
            .in3(N__48112),
            .lcout(n2920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_14_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_14_19_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1927_3_lut_LC_14_19_4 (
            .in0(N__47814),
            .in1(N__47791),
            .in2(_gnd_net_),
            .in3(N__49295),
            .lcout(n2927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_14_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_14_19_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1919_3_lut_LC_14_19_5 (
            .in0(N__49297),
            .in1(N__48061),
            .in2(N__48100),
            .in3(_gnd_net_),
            .lcout(n2919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_14_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_14_19_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1928_3_lut_LC_14_19_6 (
            .in0(N__47824),
            .in1(N__47846),
            .in2(_gnd_net_),
            .in3(N__49292),
            .lcout(n2928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_14_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_14_19_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1922_3_lut_LC_14_19_7 (
            .in0(N__49294),
            .in1(_gnd_net_),
            .in2(N__48234),
            .in3(N__48202),
            .lcout(n2922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12351_3_lut_LC_14_20_1.C_ON=1'b0;
    defparam i12351_3_lut_LC_14_20_1.SEQ_MODE=4'b0000;
    defparam i12351_3_lut_LC_14_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12351_3_lut_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(N__44515),
            .in2(N__44503),
            .in3(N__47595),
            .lcout(n2825),
            .ltout(n2825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_14_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_14_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_14_20_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1924_3_lut_LC_14_20_2 (
            .in0(N__49326),
            .in1(_gnd_net_),
            .in2(N__44470),
            .in3(N__48286),
            .lcout(n2924),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_14_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_14_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_14_20_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1925_3_lut_LC_14_20_3 (
            .in0(_gnd_net_),
            .in1(N__47736),
            .in2(N__47707),
            .in3(N__49325),
            .lcout(n2925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_14_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_14_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_14_20_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2058_3_lut_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(N__44979),
            .in2(N__44965),
            .in3(N__49065),
            .lcout(n3122),
            .ltout(n3122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_14_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_14_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_14_20_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i2125_3_lut_LC_14_20_5 (
            .in0(N__51325),
            .in1(_gnd_net_),
            .in2(N__44923),
            .in3(N__50108),
            .lcout(n3221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_14_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_14_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_14_20_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1914_3_lut_LC_14_20_6 (
            .in0(_gnd_net_),
            .in1(N__48504),
            .in2(N__49358),
            .in3(N__48481),
            .lcout(n2914),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_14_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_14_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_14_20_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2062_3_lut_LC_14_20_7 (
            .in0(N__45097),
            .in1(_gnd_net_),
            .in2(N__49083),
            .in3(N__45117),
            .lcout(n3126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_14_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_14_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_14_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_2_lut_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(N__44893),
            .in2(_gnd_net_),
            .in3(N__44839),
            .lcout(n3101),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(n12464),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_14_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_14_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_14_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_3_lut_LC_14_21_1 (
            .in0(_gnd_net_),
            .in1(N__55190),
            .in2(N__44836),
            .in3(N__44791),
            .lcout(n3100),
            .ltout(),
            .carryin(n12464),
            .carryout(n12465),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_14_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_14_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_14_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_4_lut_LC_14_21_2 (
            .in0(_gnd_net_),
            .in1(N__44787),
            .in2(_gnd_net_),
            .in3(N__44746),
            .lcout(n3099),
            .ltout(),
            .carryin(n12465),
            .carryout(n12466),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_14_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_14_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_14_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_5_lut_LC_14_21_3 (
            .in0(_gnd_net_),
            .in1(N__55191),
            .in2(N__44743),
            .in3(N__44710),
            .lcout(n3098),
            .ltout(),
            .carryin(n12466),
            .carryout(n12467),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_14_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_14_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_14_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_6_lut_LC_14_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45229),
            .in3(N__45190),
            .lcout(n3097),
            .ltout(),
            .carryin(n12467),
            .carryout(n12468),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_14_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_14_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_14_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_7_lut_LC_14_21_5 (
            .in0(_gnd_net_),
            .in1(N__45187),
            .in2(_gnd_net_),
            .in3(N__45157),
            .lcout(n3096),
            .ltout(),
            .carryin(n12468),
            .carryout(n12469),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_14_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_14_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_14_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_8_lut_LC_14_21_6 (
            .in0(_gnd_net_),
            .in1(N__55060),
            .in2(N__45154),
            .in3(N__45121),
            .lcout(n3095),
            .ltout(),
            .carryin(n12469),
            .carryout(n12470),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_14_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_14_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_14_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_9_lut_LC_14_21_7 (
            .in0(_gnd_net_),
            .in1(N__55192),
            .in2(N__45118),
            .in3(N__45091),
            .lcout(n3094),
            .ltout(),
            .carryin(n12470),
            .carryout(n12471),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_14_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_14_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_14_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_10_lut_LC_14_22_0 (
            .in0(_gnd_net_),
            .in1(N__54618),
            .in2(N__45088),
            .in3(N__45061),
            .lcout(n3093),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(n12472),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_14_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_14_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_14_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_11_lut_LC_14_22_1 (
            .in0(_gnd_net_),
            .in1(N__54340),
            .in2(N__45058),
            .in3(N__45016),
            .lcout(n3092),
            .ltout(),
            .carryin(n12472),
            .carryout(n12473),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_14_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_14_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_14_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_12_lut_LC_14_22_2 (
            .in0(_gnd_net_),
            .in1(N__54619),
            .in2(N__45013),
            .in3(N__44983),
            .lcout(n3091),
            .ltout(),
            .carryin(n12473),
            .carryout(n12474),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_14_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_14_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_13_lut_LC_14_22_3 (
            .in0(_gnd_net_),
            .in1(N__54341),
            .in2(N__44980),
            .in3(N__44953),
            .lcout(n3090),
            .ltout(),
            .carryin(n12474),
            .carryout(n12475),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_14_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_14_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_14_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_14_lut_LC_14_22_4 (
            .in0(_gnd_net_),
            .in1(N__54620),
            .in2(N__45496),
            .in3(N__45460),
            .lcout(n3089),
            .ltout(),
            .carryin(n12475),
            .carryout(n12476),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_14_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_14_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_14_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_15_lut_LC_14_22_5 (
            .in0(_gnd_net_),
            .in1(N__54342),
            .in2(N__45457),
            .in3(N__45433),
            .lcout(n3088),
            .ltout(),
            .carryin(n12476),
            .carryout(n12477),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_14_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_14_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_14_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_16_lut_LC_14_22_6 (
            .in0(_gnd_net_),
            .in1(N__54621),
            .in2(N__45430),
            .in3(N__45385),
            .lcout(n3087),
            .ltout(),
            .carryin(n12477),
            .carryout(n12478),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_14_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_14_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_14_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_17_lut_LC_14_22_7 (
            .in0(_gnd_net_),
            .in1(N__45382),
            .in2(N__54979),
            .in3(N__45352),
            .lcout(n3086),
            .ltout(),
            .carryin(n12478),
            .carryout(n12479),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_14_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_14_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_14_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_18_lut_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(N__54649),
            .in2(N__45349),
            .in3(N__45310),
            .lcout(n3085),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(n12480),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_14_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_14_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_14_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_19_lut_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(N__45307),
            .in2(N__54988),
            .in3(N__45277),
            .lcout(n3084),
            .ltout(),
            .carryin(n12480),
            .carryout(n12481),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_14_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_14_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_14_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_20_lut_LC_14_23_2 (
            .in0(_gnd_net_),
            .in1(N__45274),
            .in2(N__55247),
            .in3(N__45235),
            .lcout(n3083),
            .ltout(),
            .carryin(n12481),
            .carryout(n12482),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_14_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_14_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_14_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_21_lut_LC_14_23_3 (
            .in0(_gnd_net_),
            .in1(N__49125),
            .in2(N__54989),
            .in3(N__45232),
            .lcout(n3082),
            .ltout(),
            .carryin(n12482),
            .carryout(n12483),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_14_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_14_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_14_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_22_lut_LC_14_23_4 (
            .in0(_gnd_net_),
            .in1(N__45732),
            .in2(N__55248),
            .in3(N__45712),
            .lcout(n3081),
            .ltout(),
            .carryin(n12483),
            .carryout(n12484),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_14_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_14_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_14_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_23_lut_LC_14_23_5 (
            .in0(_gnd_net_),
            .in1(N__45709),
            .in2(N__54990),
            .in3(N__45673),
            .lcout(n3080),
            .ltout(),
            .carryin(n12484),
            .carryout(n12485),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_14_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_14_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_14_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_24_lut_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__45669),
            .in2(N__55249),
            .in3(N__45637),
            .lcout(n3079),
            .ltout(),
            .carryin(n12485),
            .carryout(n12486),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_14_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_14_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_14_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_25_lut_LC_14_23_7 (
            .in0(_gnd_net_),
            .in1(N__49470),
            .in2(N__54991),
            .in3(N__45634),
            .lcout(n3078),
            .ltout(),
            .carryin(n12486),
            .carryout(n12487),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_14_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_14_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_14_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_26_lut_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__54669),
            .in2(N__45631),
            .in3(N__45595),
            .lcout(n3077),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(n12488),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_14_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_14_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_14_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_27_lut_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(N__49185),
            .in2(N__54994),
            .in3(N__45592),
            .lcout(n3076),
            .ltout(),
            .carryin(n12488),
            .carryout(n12489),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_14_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_14_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_14_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_28_lut_LC_14_24_2 (
            .in0(_gnd_net_),
            .in1(N__45589),
            .in2(N__54978),
            .in3(N__45547),
            .lcout(n3075),
            .ltout(),
            .carryin(n12489),
            .carryout(n12490),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_14_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_14_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_29_lut_LC_14_24_3 (
            .in0(_gnd_net_),
            .in1(N__45544),
            .in2(N__54995),
            .in3(N__45499),
            .lcout(n3074),
            .ltout(),
            .carryin(n12490),
            .carryout(n12491),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_14_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_14_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_14_24_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_2039_30_lut_LC_14_24_4 (
            .in0(N__54609),
            .in1(N__45939),
            .in2(N__45916),
            .in3(N__45889),
            .lcout(n3105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_14_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_14_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_14_24_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2128_3_lut_LC_14_24_5 (
            .in0(_gnd_net_),
            .in1(N__51497),
            .in2(N__51466),
            .in3(N__50068),
            .lcout(n3224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2199_3_lut_LC_14_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2199_3_lut_LC_14_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2199_3_lut_LC_14_24_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2199_3_lut_LC_14_24_6 (
            .in0(_gnd_net_),
            .in1(N__45886),
            .in2(N__49612),
            .in3(N__45783),
            .lcout(n15_adj_704),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_14_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_14_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_14_24_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2198_3_lut_LC_14_24_7 (
            .in0(_gnd_net_),
            .in1(N__46108),
            .in2(N__45880),
            .in3(N__49589),
            .lcout(n17_adj_705),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_152_LC_14_25_0.C_ON=1'b0;
    defparam i1_4_lut_adj_152_LC_14_25_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_152_LC_14_25_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_152_LC_14_25_0 (
            .in0(N__49655),
            .in1(N__46106),
            .in2(N__45745),
            .in3(N__45863),
            .lcout(),
            .ltout(n14368_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_153_LC_14_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_153_LC_14_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_153_LC_14_25_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_153_LC_14_25_1 (
            .in0(N__45833),
            .in1(N__49688),
            .in2(N__45805),
            .in3(N__46114),
            .lcout(n14374),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_14_25_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_14_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_14_25_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2132_3_lut_LC_14_25_3 (
            .in0(_gnd_net_),
            .in1(N__50929),
            .in2(N__50896),
            .in3(N__50113),
            .lcout(n3228),
            .ltout(n3228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_150_LC_14_25_4.C_ON=1'b0;
    defparam i1_2_lut_adj_150_LC_14_25_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_150_LC_14_25_4.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_150_LC_14_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45769),
            .in3(N__45758),
            .lcout(n14362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_151_LC_14_25_5.C_ON=1'b0;
    defparam i1_4_lut_adj_151_LC_14_25_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_151_LC_14_25_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_151_LC_14_25_5 (
            .in0(N__49386),
            .in1(N__48741),
            .in2(N__46141),
            .in3(N__48639),
            .lcout(n14366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_14_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_14_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_14_25_6.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i2131_3_lut_LC_14_25_6 (
            .in0(N__50877),
            .in1(N__50839),
            .in2(N__50119),
            .in3(_gnd_net_),
            .lcout(n3227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_14_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_14_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_14_25_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2123_3_lut_LC_14_25_7 (
            .in0(_gnd_net_),
            .in1(N__51272),
            .in2(N__51241),
            .in3(N__50117),
            .lcout(n3219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i0_LC_14_26_0.C_ON=1'b1;
    defparam duty_i0_LC_14_26_0.SEQ_MODE=4'b1000;
    defparam duty_i0_LC_14_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i0_LC_14_26_0 (
            .in0(_gnd_net_),
            .in1(N__51880),
            .in2(N__46090),
            .in3(N__46078),
            .lcout(duty_0),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(n12073),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i1_LC_14_26_1.C_ON=1'b1;
    defparam duty_i1_LC_14_26_1.SEQ_MODE=4'b1000;
    defparam duty_i1_LC_14_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i1_LC_14_26_1 (
            .in0(_gnd_net_),
            .in1(N__52474),
            .in2(N__46075),
            .in3(N__46063),
            .lcout(duty_1),
            .ltout(),
            .carryin(n12073),
            .carryout(n12074),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i2_LC_14_26_2.C_ON=1'b1;
    defparam duty_i2_LC_14_26_2.SEQ_MODE=4'b1000;
    defparam duty_i2_LC_14_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i2_LC_14_26_2 (
            .in0(_gnd_net_),
            .in1(N__46060),
            .in2(N__52447),
            .in3(N__46030),
            .lcout(duty_2),
            .ltout(),
            .carryin(n12074),
            .carryout(n12075),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i3_LC_14_26_3.C_ON=1'b1;
    defparam duty_i3_LC_14_26_3.SEQ_MODE=4'b1000;
    defparam duty_i3_LC_14_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i3_LC_14_26_3 (
            .in0(_gnd_net_),
            .in1(N__52414),
            .in2(N__46027),
            .in3(N__46018),
            .lcout(duty_3),
            .ltout(),
            .carryin(n12075),
            .carryout(n12076),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i4_LC_14_26_4.C_ON=1'b1;
    defparam duty_i4_LC_14_26_4.SEQ_MODE=4'b1000;
    defparam duty_i4_LC_14_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i4_LC_14_26_4 (
            .in0(_gnd_net_),
            .in1(N__52387),
            .in2(N__46015),
            .in3(N__45979),
            .lcout(duty_4),
            .ltout(),
            .carryin(n12076),
            .carryout(n12077),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i5_LC_14_26_5.C_ON=1'b1;
    defparam duty_i5_LC_14_26_5.SEQ_MODE=4'b1000;
    defparam duty_i5_LC_14_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i5_LC_14_26_5 (
            .in0(_gnd_net_),
            .in1(N__52357),
            .in2(N__45976),
            .in3(N__45943),
            .lcout(duty_5),
            .ltout(),
            .carryin(n12077),
            .carryout(n12078),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i6_LC_14_26_6.C_ON=1'b1;
    defparam duty_i6_LC_14_26_6.SEQ_MODE=4'b1000;
    defparam duty_i6_LC_14_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i6_LC_14_26_6 (
            .in0(_gnd_net_),
            .in1(N__52332),
            .in2(N__55531),
            .in3(N__46303),
            .lcout(duty_6),
            .ltout(),
            .carryin(n12078),
            .carryout(n12079),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i7_LC_14_26_7.C_ON=1'b1;
    defparam duty_i7_LC_14_26_7.SEQ_MODE=4'b1000;
    defparam duty_i7_LC_14_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i7_LC_14_26_7 (
            .in0(_gnd_net_),
            .in1(N__52306),
            .in2(N__46300),
            .in3(N__46288),
            .lcout(duty_7),
            .ltout(),
            .carryin(n12079),
            .carryout(n12080),
            .clk(N__56072),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i8_LC_14_27_0.C_ON=1'b1;
    defparam duty_i8_LC_14_27_0.SEQ_MODE=4'b1000;
    defparam duty_i8_LC_14_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i8_LC_14_27_0 (
            .in0(_gnd_net_),
            .in1(N__52281),
            .in2(N__46285),
            .in3(N__46270),
            .lcout(duty_8),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(n12081),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i9_LC_14_27_1.C_ON=1'b1;
    defparam duty_i9_LC_14_27_1.SEQ_MODE=4'b1000;
    defparam duty_i9_LC_14_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i9_LC_14_27_1 (
            .in0(_gnd_net_),
            .in1(N__52252),
            .in2(N__46267),
            .in3(N__46252),
            .lcout(duty_9),
            .ltout(),
            .carryin(n12081),
            .carryout(n12082),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i10_LC_14_27_2.C_ON=1'b1;
    defparam duty_i10_LC_14_27_2.SEQ_MODE=4'b1000;
    defparam duty_i10_LC_14_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i10_LC_14_27_2 (
            .in0(_gnd_net_),
            .in1(N__52701),
            .in2(N__46249),
            .in3(N__46216),
            .lcout(duty_10),
            .ltout(),
            .carryin(n12082),
            .carryout(n12083),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i11_LC_14_27_3.C_ON=1'b1;
    defparam duty_i11_LC_14_27_3.SEQ_MODE=4'b1000;
    defparam duty_i11_LC_14_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i11_LC_14_27_3 (
            .in0(_gnd_net_),
            .in1(N__52675),
            .in2(N__46213),
            .in3(N__46174),
            .lcout(duty_11),
            .ltout(),
            .carryin(n12083),
            .carryout(n12084),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i12_LC_14_27_4.C_ON=1'b1;
    defparam duty_i12_LC_14_27_4.SEQ_MODE=4'b1000;
    defparam duty_i12_LC_14_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i12_LC_14_27_4 (
            .in0(_gnd_net_),
            .in1(N__46171),
            .in2(N__52651),
            .in3(N__46159),
            .lcout(duty_12),
            .ltout(),
            .carryin(n12084),
            .carryout(n12085),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i13_LC_14_27_5.C_ON=1'b1;
    defparam duty_i13_LC_14_27_5.SEQ_MODE=4'b1000;
    defparam duty_i13_LC_14_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i13_LC_14_27_5 (
            .in0(_gnd_net_),
            .in1(N__52617),
            .in2(N__46156),
            .in3(N__46144),
            .lcout(duty_13),
            .ltout(),
            .carryin(n12085),
            .carryout(n12086),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i14_LC_14_27_6.C_ON=1'b1;
    defparam duty_i14_LC_14_27_6.SEQ_MODE=4'b1000;
    defparam duty_i14_LC_14_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i14_LC_14_27_6 (
            .in0(_gnd_net_),
            .in1(N__52591),
            .in2(N__46456),
            .in3(N__46444),
            .lcout(duty_14),
            .ltout(),
            .carryin(n12086),
            .carryout(n12087),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i15_LC_14_27_7.C_ON=1'b1;
    defparam duty_i15_LC_14_27_7.SEQ_MODE=4'b1000;
    defparam duty_i15_LC_14_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i15_LC_14_27_7 (
            .in0(_gnd_net_),
            .in1(N__46441),
            .in2(N__52558),
            .in3(N__46429),
            .lcout(duty_15),
            .ltout(),
            .carryin(n12087),
            .carryout(n12088),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i16_LC_14_28_0.C_ON=1'b1;
    defparam duty_i16_LC_14_28_0.SEQ_MODE=4'b1000;
    defparam duty_i16_LC_14_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i16_LC_14_28_0 (
            .in0(_gnd_net_),
            .in1(N__52531),
            .in2(N__46426),
            .in3(N__46414),
            .lcout(duty_16),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(n12089),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i17_LC_14_28_1.C_ON=1'b1;
    defparam duty_i17_LC_14_28_1.SEQ_MODE=4'b1000;
    defparam duty_i17_LC_14_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i17_LC_14_28_1 (
            .in0(_gnd_net_),
            .in1(N__46411),
            .in2(N__52507),
            .in3(N__46402),
            .lcout(duty_17),
            .ltout(),
            .carryin(n12089),
            .carryout(n12090),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i18_LC_14_28_2.C_ON=1'b1;
    defparam duty_i18_LC_14_28_2.SEQ_MODE=4'b1000;
    defparam duty_i18_LC_14_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i18_LC_14_28_2 (
            .in0(_gnd_net_),
            .in1(N__46399),
            .in2(N__55396),
            .in3(N__46390),
            .lcout(duty_18),
            .ltout(),
            .carryin(n12090),
            .carryout(n12091),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i19_LC_14_28_3.C_ON=1'b1;
    defparam duty_i19_LC_14_28_3.SEQ_MODE=4'b1000;
    defparam duty_i19_LC_14_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i19_LC_14_28_3 (
            .in0(_gnd_net_),
            .in1(N__46387),
            .in2(N__55366),
            .in3(N__46375),
            .lcout(duty_19),
            .ltout(),
            .carryin(n12091),
            .carryout(n12092),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i20_LC_14_28_4.C_ON=1'b1;
    defparam duty_i20_LC_14_28_4.SEQ_MODE=4'b1000;
    defparam duty_i20_LC_14_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i20_LC_14_28_4 (
            .in0(_gnd_net_),
            .in1(N__46372),
            .in2(N__55333),
            .in3(N__46363),
            .lcout(duty_20),
            .ltout(),
            .carryin(n12092),
            .carryout(n12093),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i21_LC_14_28_5.C_ON=1'b1;
    defparam duty_i21_LC_14_28_5.SEQ_MODE=4'b1000;
    defparam duty_i21_LC_14_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i21_LC_14_28_5 (
            .in0(_gnd_net_),
            .in1(N__46360),
            .in2(N__55306),
            .in3(N__46324),
            .lcout(duty_21),
            .ltout(),
            .carryin(n12093),
            .carryout(n12094),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i22_LC_14_28_6.C_ON=1'b1;
    defparam duty_i22_LC_14_28_6.SEQ_MODE=4'b1000;
    defparam duty_i22_LC_14_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i22_LC_14_28_6 (
            .in0(_gnd_net_),
            .in1(N__46621),
            .in2(N__55276),
            .in3(N__46609),
            .lcout(duty_22),
            .ltout(),
            .carryin(n12094),
            .carryout(n12095),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i23_LC_14_28_7.C_ON=1'b0;
    defparam duty_i23_LC_14_28_7.SEQ_MODE=4'b1000;
    defparam duty_i23_LC_14_28_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 duty_i23_LC_14_28_7 (
            .in0(N__52918),
            .in1(N__46606),
            .in2(_gnd_net_),
            .in3(N__46597),
            .lcout(duty_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i13_LC_14_29_0.C_ON=1'b0;
    defparam pwm_setpoint_i13_LC_14_29_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i13_LC_14_29_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i13_LC_14_29_0 (
            .in0(N__55652),
            .in1(N__46504),
            .in2(_gnd_net_),
            .in3(N__46594),
            .lcout(pwm_setpoint_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56083),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i16_1_lut_LC_14_29_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_14_29_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_14_29_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i16_1_lut_LC_14_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46584),
            .lcout(n10_adj_576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i14_LC_14_29_2.C_ON=1'b0;
    defparam pwm_setpoint_i14_LC_14_29_2.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i14_LC_14_29_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i14_LC_14_29_2 (
            .in0(N__55653),
            .in1(N__46564),
            .in2(_gnd_net_),
            .in3(N__46549),
            .lcout(pwm_setpoint_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56083),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i4_4_lut_LC_14_29_3.C_ON=1'b0;
    defparam LessThan_275_i4_4_lut_LC_14_29_3.SEQ_MODE=4'b0000;
    defparam LessThan_275_i4_4_lut_LC_14_29_3.LUT_INIT=16'b0100110101000100;
    LogicCell40 LessThan_275_i4_4_lut_LC_14_29_3 (
            .in0(N__46543),
            .in1(N__50128),
            .in2(N__46528),
            .in3(N__46462),
            .lcout(n4_adj_605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i10_1_lut_LC_14_29_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_14_29_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_14_29_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i10_1_lut_LC_14_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52788),
            .lcout(n16_adj_582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i14_1_lut_LC_14_29_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_14_29_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_14_29_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i14_1_lut_LC_14_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46503),
            .lcout(n12_adj_578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i0_LC_14_29_6.C_ON=1'b0;
    defparam pwm_setpoint_i0_LC_14_29_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i0_LC_14_29_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i0_LC_14_29_6 (
            .in0(N__55651),
            .in1(N__46483),
            .in2(_gnd_net_),
            .in3(N__46477),
            .lcout(pwm_setpoint_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56083),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i13_1_lut_LC_14_29_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_14_29_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_14_29_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i13_1_lut_LC_14_29_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46791),
            .lcout(n13_adj_579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i29_2_lut_LC_14_30_0.C_ON=1'b0;
    defparam LessThan_275_i29_2_lut_LC_14_30_0.SEQ_MODE=4'b0000;
    defparam LessThan_275_i29_2_lut_LC_14_30_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_275_i29_2_lut_LC_14_30_0 (
            .in0(N__46768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46677),
            .lcout(n29_adj_622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i27_2_lut_LC_14_30_1.C_ON=1'b0;
    defparam LessThan_275_i27_2_lut_LC_14_30_1.SEQ_MODE=4'b0000;
    defparam LessThan_275_i27_2_lut_LC_14_30_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_275_i27_2_lut_LC_14_30_1 (
            .in0(_gnd_net_),
            .in1(N__46695),
            .in2(_gnd_net_),
            .in3(N__46743),
            .lcout(n27_adj_621),
            .ltout(n27_adj_621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12368_3_lut_LC_14_30_2.C_ON=1'b0;
    defparam i12368_3_lut_LC_14_30_2.SEQ_MODE=4'b0000;
    defparam i12368_3_lut_LC_14_30_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12368_3_lut_LC_14_30_2 (
            .in0(N__46696),
            .in1(_gnd_net_),
            .in2(N__46687),
            .in3(N__46684),
            .lcout(),
            .ltout(n14840_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12369_3_lut_LC_14_30_3.C_ON=1'b0;
    defparam i12369_3_lut_LC_14_30_3.SEQ_MODE=4'b0000;
    defparam i12369_3_lut_LC_14_30_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 i12369_3_lut_LC_14_30_3 (
            .in0(N__46678),
            .in1(_gnd_net_),
            .in2(N__46669),
            .in3(N__47171),
            .lcout(n14841),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i23_1_lut_LC_14_30_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_14_30_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_14_30_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i23_1_lut_LC_14_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46665),
            .lcout(n3_adj_569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i17_1_lut_LC_14_30_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_14_30_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_14_30_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 unary_minus_13_inv_0_i17_1_lut_LC_14_30_5 (
            .in0(N__46638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n9_adj_575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i16_LC_14_30_6.C_ON=1'b0;
    defparam pwm_setpoint_i16_LC_14_30_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i16_LC_14_30_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i16_LC_14_30_6 (
            .in0(N__55654),
            .in1(N__46639),
            .in2(_gnd_net_),
            .in3(N__46627),
            .lcout(pwm_setpoint_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56087),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i21_1_lut_LC_14_30_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_14_30_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_14_30_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i21_1_lut_LC_14_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47061),
            .lcout(n5_adj_571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12250_2_lut_4_lut_LC_14_31_0.C_ON=1'b0;
    defparam i12250_2_lut_4_lut_LC_14_31_0.SEQ_MODE=4'b0000;
    defparam i12250_2_lut_4_lut_LC_14_31_0.LUT_INIT=16'b0110111111110110;
    LogicCell40 i12250_2_lut_4_lut_LC_14_31_0 (
            .in0(N__46842),
            .in1(N__46859),
            .in2(N__47038),
            .in3(N__46926),
            .lcout(),
            .ltout(n14722_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12404_4_lut_LC_14_31_1.C_ON=1'b0;
    defparam i12404_4_lut_LC_14_31_1.SEQ_MODE=4'b0000;
    defparam i12404_4_lut_LC_14_31_1.LUT_INIT=16'b1111111000000010;
    LogicCell40 i12404_4_lut_LC_14_31_1 (
            .in0(N__47005),
            .in1(N__46886),
            .in2(N__46993),
            .in3(N__46867),
            .lcout(),
            .ltout(n14876_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12414_4_lut_LC_14_31_2.C_ON=1'b0;
    defparam i12414_4_lut_LC_14_31_2.SEQ_MODE=4'b0000;
    defparam i12414_4_lut_LC_14_31_2.LUT_INIT=16'b1111000111100000;
    LogicCell40 i12414_4_lut_LC_14_31_2 (
            .in0(N__46887),
            .in1(N__47158),
            .in2(N__46990),
            .in3(N__46963),
            .lcout(n14886),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12309_3_lut_LC_14_31_6.C_ON=1'b0;
    defparam i12309_3_lut_LC_14_31_6.SEQ_MODE=4'b0000;
    defparam i12309_3_lut_LC_14_31_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12309_3_lut_LC_14_31_6 (
            .in0(N__47210),
            .in1(N__46981),
            .in2(_gnd_net_),
            .in3(N__46969),
            .lcout(n14781),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i7_LC_14_31_7.C_ON=1'b0;
    defparam pwm_setpoint_i7_LC_14_31_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i7_LC_14_31_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i7_LC_14_31_7 (
            .in0(N__55694),
            .in1(N__46957),
            .in2(_gnd_net_),
            .in3(N__46947),
            .lcout(pwm_setpoint_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56091),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i12_3_lut_3_lut_LC_14_32_0.C_ON=1'b0;
    defparam LessThan_275_i12_3_lut_3_lut_LC_14_32_0.SEQ_MODE=4'b0000;
    defparam LessThan_275_i12_3_lut_3_lut_LC_14_32_0.LUT_INIT=16'b1101110101000100;
    LogicCell40 LessThan_275_i12_3_lut_3_lut_LC_14_32_0 (
            .in0(N__46840),
            .in1(N__46860),
            .in2(_gnd_net_),
            .in3(N__46922),
            .lcout(),
            .ltout(n12_adj_611_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i30_3_lut_LC_14_32_1.C_ON=1'b0;
    defparam LessThan_275_i30_3_lut_LC_14_32_1.SEQ_MODE=4'b0000;
    defparam LessThan_275_i30_3_lut_LC_14_32_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 LessThan_275_i30_3_lut_LC_14_32_1 (
            .in0(_gnd_net_),
            .in1(N__46906),
            .in2(N__46894),
            .in3(N__46885),
            .lcout(n30_adj_623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_275_i33_2_lut_LC_14_32_3.C_ON=1'b0;
    defparam LessThan_275_i33_2_lut_LC_14_32_3.SEQ_MODE=4'b0000;
    defparam LessThan_275_i33_2_lut_LC_14_32_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_275_i33_2_lut_LC_14_32_3 (
            .in0(N__46861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46841),
            .lcout(n33_adj_625),
            .ltout(n33_adj_625_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12252_4_lut_LC_14_32_4.C_ON=1'b0;
    defparam i12252_4_lut_LC_14_32_4.SEQ_MODE=4'b0000;
    defparam i12252_4_lut_LC_14_32_4.LUT_INIT=16'b1111000011110001;
    LogicCell40 i12252_4_lut_LC_14_32_4 (
            .in0(N__47211),
            .in1(N__47194),
            .in2(N__47182),
            .in3(N__47178),
            .lcout(n14724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i18_1_lut_LC_14_32_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_14_32_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_14_32_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i18_1_lut_LC_14_32_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47148),
            .lcout(n8_adj_574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_162_LC_15_17_0.C_ON=1'b0;
    defparam i10_4_lut_adj_162_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_162_LC_15_17_0.LUT_INIT=16'b1111111111111101;
    LogicCell40 i10_4_lut_adj_162_LC_15_17_0 (
            .in0(N__50535),
            .in1(N__50220),
            .in2(N__50572),
            .in3(N__50601),
            .lcout(n28_adj_597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_15_17_7.C_ON=1'b0;
    defparam i13_4_lut_LC_15_17_7.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_15_17_7.LUT_INIT=16'b1111111110111111;
    LogicCell40 i13_4_lut_LC_15_17_7 (
            .in0(N__50649),
            .in1(N__50745),
            .in2(N__50716),
            .in3(N__50586),
            .lcout(n31_adj_594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_3_lut_adj_163_LC_15_18_1.C_ON=1'b0;
    defparam i14_3_lut_adj_163_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam i14_3_lut_adj_163_LC_15_18_1.LUT_INIT=16'b1101110111111111;
    LogicCell40 i14_3_lut_adj_163_LC_15_18_1 (
            .in0(N__50661),
            .in1(N__47125),
            .in2(_gnd_net_),
            .in3(N__50730),
            .lcout(),
            .ltout(n32_adj_593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12759_4_lut_LC_15_18_2.C_ON=1'b0;
    defparam i12759_4_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam i12759_4_lut_LC_15_18_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12759_4_lut_LC_15_18_2 (
            .in0(N__47119),
            .in1(N__47077),
            .in2(N__47113),
            .in3(N__47071),
            .lcout(n4856),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_15_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_15_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_15_18_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1910_3_lut_LC_15_18_3 (
            .in0(_gnd_net_),
            .in1(N__48316),
            .in2(N__48336),
            .in3(N__49324),
            .lcout(n2910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_LC_15_18_5.C_ON=1'b0;
    defparam i12_4_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam i12_4_lut_LC_15_18_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_LC_15_18_5 (
            .in0(N__50616),
            .in1(N__50520),
            .in2(N__50635),
            .in3(N__50760),
            .lcout(n30_adj_595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_15_18_6.C_ON=1'b0;
    defparam i11_4_lut_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_15_18_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_LC_15_18_6 (
            .in0(N__50679),
            .in1(N__50775),
            .in2(N__50698),
            .in3(N__50550),
            .lcout(n29_adj_596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_15_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_15_19_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1865_3_lut_LC_15_19_0 (
            .in0(N__47695),
            .in1(N__47682),
            .in2(_gnd_net_),
            .in3(N__47616),
            .lcout(n2833),
            .ltout(n2833_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10041_4_lut_LC_15_19_1.C_ON=1'b0;
    defparam i10041_4_lut_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam i10041_4_lut_LC_15_19_1.LUT_INIT=16'b1111111010101010;
    LogicCell40 i10041_4_lut_LC_15_19_1 (
            .in0(N__47921),
            .in1(N__47256),
            .in2(N__47473),
            .in3(N__47951),
            .lcout(n11756),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_15_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_15_19_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1931_3_lut_LC_15_19_2 (
            .in0(N__47952),
            .in1(_gnd_net_),
            .in2(N__49340),
            .in3(N__47935),
            .lcout(n2931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_15_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_15_19_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1932_3_lut_LC_15_19_3 (
            .in0(_gnd_net_),
            .in1(N__47982),
            .in2(N__47968),
            .in3(N__49298),
            .lcout(n2932),
            .ltout(n2932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9947_3_lut_LC_15_19_4.C_ON=1'b0;
    defparam i9947_3_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam i9947_3_lut_LC_15_19_4.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9947_3_lut_LC_15_19_4 (
            .in0(_gnd_net_),
            .in1(N__47434),
            .in2(N__47410),
            .in3(N__47396),
            .lcout(n11662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_15_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_15_19_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1930_3_lut_LC_15_19_5 (
            .in0(N__47922),
            .in1(_gnd_net_),
            .in2(N__47905),
            .in3(N__49302),
            .lcout(n2930),
            .ltout(n2930_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_40_LC_15_19_6.C_ON=1'b0;
    defparam i1_4_lut_adj_40_LC_15_19_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_40_LC_15_19_6.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_40_LC_15_19_6 (
            .in0(N__47333),
            .in1(N__47303),
            .in2(N__47284),
            .in3(N__47281),
            .lcout(n13417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_15_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_15_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_15_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_2_lut_LC_15_20_0 (
            .in0(_gnd_net_),
            .in1(N__47249),
            .in2(_gnd_net_),
            .in3(N__47215),
            .lcout(n2901),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(n12411),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_15_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_15_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_3_lut_LC_15_20_1 (
            .in0(_gnd_net_),
            .in1(N__54610),
            .in2(N__47983),
            .in3(N__47959),
            .lcout(n2900),
            .ltout(),
            .carryin(n12411),
            .carryout(n12412),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_15_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_15_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_15_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_4_lut_LC_15_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47956),
            .in3(N__47929),
            .lcout(n2899),
            .ltout(),
            .carryin(n12412),
            .carryout(n12413),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_15_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_15_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_15_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_5_lut_LC_15_20_3 (
            .in0(_gnd_net_),
            .in1(N__54611),
            .in2(N__47926),
            .in3(N__47896),
            .lcout(n2898),
            .ltout(),
            .carryin(n12413),
            .carryout(n12414),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_15_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_15_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_6_lut_LC_15_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47893),
            .in3(N__47857),
            .lcout(n2897),
            .ltout(),
            .carryin(n12414),
            .carryout(n12415),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_15_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_15_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_7_lut_LC_15_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47854),
            .in3(N__47818),
            .lcout(n2896),
            .ltout(),
            .carryin(n12415),
            .carryout(n12416),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_15_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_15_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_15_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_8_lut_LC_15_20_6 (
            .in0(_gnd_net_),
            .in1(N__54613),
            .in2(N__47815),
            .in3(N__47785),
            .lcout(n2895),
            .ltout(),
            .carryin(n12416),
            .carryout(n12417),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_15_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_15_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_15_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_9_lut_LC_15_20_7 (
            .in0(_gnd_net_),
            .in1(N__54612),
            .in2(N__47781),
            .in3(N__47740),
            .lcout(n2894),
            .ltout(),
            .carryin(n12417),
            .carryout(n12418),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_15_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_15_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_15_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_10_lut_LC_15_21_0 (
            .in0(_gnd_net_),
            .in1(N__55233),
            .in2(N__47737),
            .in3(N__47698),
            .lcout(n2893),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(n12419),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_15_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_15_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_15_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_11_lut_LC_15_21_1 (
            .in0(_gnd_net_),
            .in1(N__54614),
            .in2(N__48304),
            .in3(N__48280),
            .lcout(n2892),
            .ltout(),
            .carryin(n12419),
            .carryout(n12420),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_15_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_15_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_15_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_12_lut_LC_15_21_2 (
            .in0(_gnd_net_),
            .in1(N__55234),
            .in2(N__48277),
            .in3(N__48238),
            .lcout(n2891),
            .ltout(),
            .carryin(n12420),
            .carryout(n12421),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_15_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_15_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_15_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_13_lut_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(N__54615),
            .in2(N__48235),
            .in3(N__48193),
            .lcout(n2890),
            .ltout(),
            .carryin(n12421),
            .carryout(n12422),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_15_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_15_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_14_lut_LC_15_21_4 (
            .in0(_gnd_net_),
            .in1(N__55235),
            .in2(N__48190),
            .in3(N__48145),
            .lcout(n2889),
            .ltout(),
            .carryin(n12422),
            .carryout(n12423),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_15_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_15_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_15_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_15_lut_LC_15_21_5 (
            .in0(_gnd_net_),
            .in1(N__54616),
            .in2(N__48142),
            .in3(N__48103),
            .lcout(n2888),
            .ltout(),
            .carryin(n12423),
            .carryout(n12424),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_15_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_15_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_15_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_16_lut_LC_15_21_6 (
            .in0(_gnd_net_),
            .in1(N__55236),
            .in2(N__48099),
            .in3(N__48052),
            .lcout(n2887),
            .ltout(),
            .carryin(n12424),
            .carryout(n12425),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_15_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_15_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_15_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_17_lut_LC_15_21_7 (
            .in0(_gnd_net_),
            .in1(N__54617),
            .in2(N__48049),
            .in3(N__48010),
            .lcout(n2886),
            .ltout(),
            .carryin(n12425),
            .carryout(n12426),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_15_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_15_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_18_lut_LC_15_22_0 (
            .in0(_gnd_net_),
            .in1(N__48007),
            .in2(N__54980),
            .in3(N__48592),
            .lcout(n2885),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(n12427),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_15_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_15_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_19_lut_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(N__48589),
            .in2(N__54984),
            .in3(N__48556),
            .lcout(n2884),
            .ltout(),
            .carryin(n12427),
            .carryout(n12428),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_15_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_15_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_20_lut_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(N__48552),
            .in2(N__54981),
            .in3(N__48508),
            .lcout(n2883),
            .ltout(),
            .carryin(n12428),
            .carryout(n12429),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_15_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_15_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_15_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_21_lut_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(N__48505),
            .in2(N__54985),
            .in3(N__48472),
            .lcout(n2882),
            .ltout(),
            .carryin(n12429),
            .carryout(n12430),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_15_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_15_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_22_lut_LC_15_22_4 (
            .in0(_gnd_net_),
            .in1(N__48465),
            .in2(N__54982),
            .in3(N__48433),
            .lcout(n2881),
            .ltout(),
            .carryin(n12430),
            .carryout(n12431),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_15_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_15_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_15_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_23_lut_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(N__48430),
            .in2(N__54986),
            .in3(N__48388),
            .lcout(n2880),
            .ltout(),
            .carryin(n12431),
            .carryout(n12432),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_15_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_15_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_24_lut_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(N__48385),
            .in2(N__54983),
            .in3(N__48340),
            .lcout(n2879),
            .ltout(),
            .carryin(n12432),
            .carryout(n12433),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_15_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_15_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_15_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_25_lut_LC_15_22_7 (
            .in0(_gnd_net_),
            .in1(N__48337),
            .in2(N__54987),
            .in3(N__48307),
            .lcout(n2878),
            .ltout(),
            .carryin(n12433),
            .carryout(n12434),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_15_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_15_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_15_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_26_lut_LC_15_23_0 (
            .in0(_gnd_net_),
            .in1(N__48907),
            .in2(N__54992),
            .in3(N__48868),
            .lcout(n2877),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(n12435),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_15_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_15_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_15_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_27_lut_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(N__48865),
            .in2(N__54993),
            .in3(N__48811),
            .lcout(n2876),
            .ltout(),
            .carryin(n12435),
            .carryout(n12436),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_15_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_15_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_15_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_28_lut_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(N__54668),
            .in2(N__48805),
            .in3(N__48808),
            .lcout(n2875),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1907_3_lut_LC_15_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1907_3_lut_LC_15_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1907_3_lut_LC_15_23_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1907_3_lut_LC_15_23_4 (
            .in0(N__48804),
            .in1(_gnd_net_),
            .in2(N__48775),
            .in3(N__49372),
            .lcout(n2907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_128_LC_15_24_1.C_ON=1'b0;
    defparam i1_4_lut_adj_128_LC_15_24_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_128_LC_15_24_1.LUT_INIT=16'b1111111110111000;
    LogicCell40 i1_4_lut_adj_128_LC_15_24_1 (
            .in0(N__48742),
            .in1(N__49616),
            .in2(N__48718),
            .in3(N__48706),
            .lcout(),
            .ltout(n13822_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_130_LC_15_24_2.C_ON=1'b0;
    defparam i1_4_lut_adj_130_LC_15_24_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_130_LC_15_24_2.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_130_LC_15_24_2 (
            .in0(N__49617),
            .in1(N__48700),
            .in2(N__48685),
            .in3(N__48681),
            .lcout(),
            .ltout(n13834_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_134_LC_15_24_3.C_ON=1'b0;
    defparam i1_4_lut_adj_134_LC_15_24_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_134_LC_15_24_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_134_LC_15_24_3 (
            .in0(N__48661),
            .in1(N__49477),
            .in2(N__48655),
            .in3(N__49672),
            .lcout(n13842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_15_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_15_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_15_24_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2193_3_lut_LC_15_24_5 (
            .in0(_gnd_net_),
            .in1(N__48643),
            .in2(N__48616),
            .in3(N__49613),
            .lcout(),
            .ltout(n27_adj_709_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_129_LC_15_24_6.C_ON=1'b0;
    defparam i1_4_lut_adj_129_LC_15_24_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_129_LC_15_24_6.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_129_LC_15_24_6 (
            .in0(N__49615),
            .in1(N__49705),
            .in2(N__49693),
            .in3(N__49690),
            .lcout(n13830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2196_3_lut_LC_15_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2196_3_lut_LC_15_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2196_3_lut_LC_15_24_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2196_3_lut_LC_15_24_7 (
            .in0(_gnd_net_),
            .in1(N__49666),
            .in2(N__49657),
            .in3(N__49614),
            .lcout(n21_adj_706),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_15_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_15_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_15_25_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2046_3_lut_LC_15_25_0 (
            .in0(N__49471),
            .in1(_gnd_net_),
            .in2(N__49447),
            .in3(N__49077),
            .lcout(n3110),
            .ltout(n3110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_15_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_15_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_15_25_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i2113_3_lut_LC_15_25_1 (
            .in0(N__50097),
            .in1(_gnd_net_),
            .in2(N__49432),
            .in3(N__52153),
            .lcout(n3209),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_15_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_15_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_15_25_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2130_3_lut_LC_15_25_2 (
            .in0(_gnd_net_),
            .in1(N__50788),
            .in2(N__50824),
            .in3(N__50095),
            .lcout(n3226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12449_1_lut_LC_15_25_3.C_ON=1'b0;
    defparam i12449_1_lut_LC_15_25_3.SEQ_MODE=4'b0000;
    defparam i12449_1_lut_LC_15_25_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12449_1_lut_LC_15_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49373),
            .lcout(n14921),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_15_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_15_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_15_25_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2044_3_lut_LC_15_25_4 (
            .in0(_gnd_net_),
            .in1(N__49189),
            .in2(N__49162),
            .in3(N__49078),
            .lcout(n3108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i0_LC_15_25_5 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i0_LC_15_25_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i0_LC_15_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i0_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49153),
            .lcout(\quad_counter0.b_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_15_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_15_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_15_25_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2050_3_lut_LC_15_25_6 (
            .in0(_gnd_net_),
            .in1(N__49129),
            .in2(N__49096),
            .in3(N__49076),
            .lcout(n3114),
            .ltout(n3114_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_15_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_15_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_15_25_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i2117_3_lut_LC_15_25_7 (
            .in0(N__50096),
            .in1(_gnd_net_),
            .in2(N__49933),
            .in3(N__51649),
            .lcout(n3213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_158_LC_15_26_2.C_ON=1'b0;
    defparam i2_2_lut_adj_158_LC_15_26_2.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_158_LC_15_26_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_adj_158_LC_15_26_2 (
            .in0(_gnd_net_),
            .in1(N__51875),
            .in2(_gnd_net_),
            .in3(N__52406),
            .lcout(),
            .ltout(n7_adj_712_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_15_26_3.C_ON=1'b0;
    defparam i2_4_lut_LC_15_26_3.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_15_26_3.LUT_INIT=16'b1000100010000000;
    LogicCell40 i2_4_lut_LC_15_26_3 (
            .in0(N__52352),
            .in1(N__52325),
            .in2(N__49900),
            .in3(N__49897),
            .lcout(n13676),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_15_26_5.C_ON=1'b0;
    defparam i3_3_lut_LC_15_26_5.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_15_26_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 i3_3_lut_LC_15_26_5 (
            .in0(N__52376),
            .in1(N__52433),
            .in2(_gnd_net_),
            .in3(N__52466),
            .lcout(n8_adj_711),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_15_27_2 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_15_27_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.b_prev_I_0_63_2_lut_LC_15_27_2  (
            .in0(_gnd_net_),
            .in1(N__50316),
            .in2(_gnd_net_),
            .in3(N__50376),
            .lcout(\quad_counter0.direction_N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_15_27_3.C_ON=1'b0;
    defparam i4_4_lut_LC_15_27_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_15_27_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_LC_15_27_3 (
            .in0(N__52694),
            .in1(N__52244),
            .in2(N__52280),
            .in3(N__49723),
            .lcout(),
            .ltout(n10_adj_714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_159_LC_15_27_4.C_ON=1'b0;
    defparam i4_4_lut_adj_159_LC_15_27_4.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_159_LC_15_27_4.LUT_INIT=16'b1010101010101000;
    LogicCell40 i4_4_lut_adj_159_LC_15_27_4 (
            .in0(N__55352),
            .in1(N__52301),
            .in2(N__49717),
            .in3(N__52670),
            .lcout(),
            .ltout(n16_adj_702_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_15_27_5.C_ON=1'b0;
    defparam i10_4_lut_LC_15_27_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_15_27_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 i10_4_lut_LC_15_27_5 (
            .in0(N__52640),
            .in1(N__55295),
            .in2(N__49714),
            .in3(N__49711),
            .lcout(n22_adj_699),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_161_LC_15_27_7.C_ON=1'b0;
    defparam i7_4_lut_adj_161_LC_15_27_7.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_161_LC_15_27_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 i7_4_lut_adj_161_LC_15_27_7 (
            .in0(N__52493),
            .in1(N__55382),
            .in2(N__52586),
            .in3(N__52550),
            .lcout(n19_adj_701),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i1_LC_15_28_2 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i1_LC_15_28_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i1_LC_15_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i1_LC_15_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50469),
            .lcout(\quad_counter0.b_new_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56084),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i2_1_lut_LC_15_28_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_15_28_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_15_28_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i2_1_lut_LC_15_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50154),
            .lcout(n24_adj_590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i4_1_lut_LC_15_28_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_15_28_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_15_28_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i4_1_lut_LC_15_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50190),
            .lcout(n22_adj_588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_15_28_5.C_ON=1'b0;
    defparam i9_4_lut_LC_15_28_5.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_15_28_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 i9_4_lut_LC_15_28_5 (
            .in0(N__55325),
            .in1(N__52526),
            .in2(N__52621),
            .in3(N__55268),
            .lcout(),
            .ltout(n21_adj_700_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12460_4_lut_LC_15_28_6.C_ON=1'b0;
    defparam i12460_4_lut_LC_15_28_6.SEQ_MODE=4'b0000;
    defparam i12460_4_lut_LC_15_28_6.LUT_INIT=16'b0000100010001000;
    LogicCell40 i12460_4_lut_LC_15_28_6 (
            .in0(N__52913),
            .in1(N__52865),
            .in2(N__50164),
            .in3(N__50161),
            .lcout(n4890),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i1_LC_15_28_7.C_ON=1'b0;
    defparam pwm_setpoint_i1_LC_15_28_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i1_LC_15_28_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 pwm_setpoint_i1_LC_15_28_7 (
            .in0(N__50155),
            .in1(N__50137),
            .in2(_gnd_net_),
            .in3(N__55644),
            .lcout(pwm_setpoint_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56084),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12421_4_lut_LC_15_29_0 .C_ON=1'b0;
    defparam \quad_counter0.i12421_4_lut_LC_15_29_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12421_4_lut_LC_15_29_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \quad_counter0.i12421_4_lut_LC_15_29_0  (
            .in0(N__50333),
            .in1(N__50483),
            .in2(N__50317),
            .in3(N__50465),
            .lcout(\quad_counter0.a_prev_N_537 ),
            .ltout(\quad_counter0.a_prev_N_537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_52_LC_15_29_1 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_52_LC_15_29_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_prev_52_LC_15_29_1 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \quad_counter0.b_prev_52_LC_15_29_1  (
            .in0(N__50484),
            .in1(N__50372),
            .in2(N__50122),
            .in3(N__50449),
            .lcout(b_prev),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56088),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_15_29_2 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_15_29_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_15_29_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.b_prev_I_0_65_2_lut_LC_15_29_2  (
            .in0(_gnd_net_),
            .in1(N__50482),
            .in2(_gnd_net_),
            .in3(N__50371),
            .lcout(),
            .ltout(\quad_counter0.direction_N_534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_15_29_3 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_15_29_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_15_29_3 .LUT_INIT=16'b1111011000000000;
    LogicCell40 \quad_counter0.debounce_cnt_I_0_4_lut_LC_15_29_3  (
            .in0(N__50309),
            .in1(N__50493),
            .in2(N__50506),
            .in3(N__50447),
            .lcout(direction_N_531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_prev_51_LC_15_29_4 .C_ON=1'b0;
    defparam \quad_counter0.a_prev_51_LC_15_29_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_prev_51_LC_15_29_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \quad_counter0.a_prev_51_LC_15_29_4  (
            .in0(N__50448),
            .in1(N__50503),
            .in2(N__50497),
            .in3(N__50310),
            .lcout(\quad_counter0.a_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56088),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_50_LC_15_29_7 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_50_LC_15_29_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.debounce_cnt_50_LC_15_29_7 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \quad_counter0.debounce_cnt_50_LC_15_29_7  (
            .in0(N__50485),
            .in1(N__50314),
            .in2(N__50470),
            .in3(N__50334),
            .lcout(\quad_counter0.debounce_cnt ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56088),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.direction_57_LC_15_30_1 .C_ON=1'b0;
    defparam \quad_counter0.direction_57_LC_15_30_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.direction_57_LC_15_30_1 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \quad_counter0.direction_57_LC_15_30_1  (
            .in0(N__50393),
            .in1(N__50315),
            .in2(N__50377),
            .in3(N__50347),
            .lcout(n1185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56092),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i1_LC_15_30_5 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i1_LC_15_30_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i1_LC_15_30_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.a_new_i1_LC_15_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50341),
            .lcout(a_new_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56092),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i20_1_lut_LC_15_30_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_15_30_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_15_30_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i20_1_lut_LC_15_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50277),
            .lcout(n6_adj_572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i19_1_lut_LC_15_31_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_15_31_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_15_31_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i19_1_lut_LC_15_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50250),
            .lcout(n7_adj_573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sweep_counter_631_632__i1_LC_16_17_0.C_ON=1'b1;
    defparam sweep_counter_631_632__i1_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i1_LC_16_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i1_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__50221),
            .in2(_gnd_net_),
            .in3(N__50209),
            .lcout(sweep_counter_0),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(n12606),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i2_LC_16_17_1.C_ON=1'b1;
    defparam sweep_counter_631_632__i2_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i2_LC_16_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i2_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(N__50650),
            .in2(_gnd_net_),
            .in3(N__50638),
            .lcout(sweep_counter_1),
            .ltout(),
            .carryin(n12606),
            .carryout(n12607),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i3_LC_16_17_2.C_ON=1'b1;
    defparam sweep_counter_631_632__i3_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i3_LC_16_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i3_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(N__50634),
            .in2(_gnd_net_),
            .in3(N__50620),
            .lcout(sweep_counter_2),
            .ltout(),
            .carryin(n12607),
            .carryout(n12608),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i4_LC_16_17_3.C_ON=1'b1;
    defparam sweep_counter_631_632__i4_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i4_LC_16_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i4_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(N__50617),
            .in2(_gnd_net_),
            .in3(N__50605),
            .lcout(sweep_counter_3),
            .ltout(),
            .carryin(n12608),
            .carryout(n12609),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i5_LC_16_17_4.C_ON=1'b1;
    defparam sweep_counter_631_632__i5_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i5_LC_16_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i5_LC_16_17_4 (
            .in0(_gnd_net_),
            .in1(N__50602),
            .in2(_gnd_net_),
            .in3(N__50590),
            .lcout(sweep_counter_4),
            .ltout(),
            .carryin(n12609),
            .carryout(n12610),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i6_LC_16_17_5.C_ON=1'b1;
    defparam sweep_counter_631_632__i6_LC_16_17_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i6_LC_16_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i6_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(N__50587),
            .in2(_gnd_net_),
            .in3(N__50575),
            .lcout(sweep_counter_5),
            .ltout(),
            .carryin(n12610),
            .carryout(n12611),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i7_LC_16_17_6.C_ON=1'b1;
    defparam sweep_counter_631_632__i7_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i7_LC_16_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i7_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(N__50571),
            .in2(_gnd_net_),
            .in3(N__50554),
            .lcout(sweep_counter_6),
            .ltout(),
            .carryin(n12611),
            .carryout(n12612),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i8_LC_16_17_7.C_ON=1'b1;
    defparam sweep_counter_631_632__i8_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i8_LC_16_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i8_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(N__50551),
            .in2(_gnd_net_),
            .in3(N__50539),
            .lcout(sweep_counter_7),
            .ltout(),
            .carryin(n12612),
            .carryout(n12613),
            .clk(N__56050),
            .ce(),
            .sr(N__52882));
    defparam sweep_counter_631_632__i9_LC_16_18_0.C_ON=1'b1;
    defparam sweep_counter_631_632__i9_LC_16_18_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i9_LC_16_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i9_LC_16_18_0 (
            .in0(_gnd_net_),
            .in1(N__50536),
            .in2(_gnd_net_),
            .in3(N__50524),
            .lcout(sweep_counter_8),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(n12614),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i10_LC_16_18_1.C_ON=1'b1;
    defparam sweep_counter_631_632__i10_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i10_LC_16_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i10_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(N__50521),
            .in2(_gnd_net_),
            .in3(N__50509),
            .lcout(sweep_counter_9),
            .ltout(),
            .carryin(n12614),
            .carryout(n12615),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i11_LC_16_18_2.C_ON=1'b1;
    defparam sweep_counter_631_632__i11_LC_16_18_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i11_LC_16_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i11_LC_16_18_2 (
            .in0(_gnd_net_),
            .in1(N__50776),
            .in2(_gnd_net_),
            .in3(N__50764),
            .lcout(sweep_counter_10),
            .ltout(),
            .carryin(n12615),
            .carryout(n12616),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i12_LC_16_18_3.C_ON=1'b1;
    defparam sweep_counter_631_632__i12_LC_16_18_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i12_LC_16_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i12_LC_16_18_3 (
            .in0(_gnd_net_),
            .in1(N__50761),
            .in2(_gnd_net_),
            .in3(N__50749),
            .lcout(sweep_counter_11),
            .ltout(),
            .carryin(n12616),
            .carryout(n12617),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i13_LC_16_18_4.C_ON=1'b1;
    defparam sweep_counter_631_632__i13_LC_16_18_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i13_LC_16_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i13_LC_16_18_4 (
            .in0(_gnd_net_),
            .in1(N__50746),
            .in2(_gnd_net_),
            .in3(N__50734),
            .lcout(sweep_counter_12),
            .ltout(),
            .carryin(n12617),
            .carryout(n12618),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i14_LC_16_18_5.C_ON=1'b1;
    defparam sweep_counter_631_632__i14_LC_16_18_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i14_LC_16_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i14_LC_16_18_5 (
            .in0(_gnd_net_),
            .in1(N__50731),
            .in2(_gnd_net_),
            .in3(N__50719),
            .lcout(sweep_counter_13),
            .ltout(),
            .carryin(n12618),
            .carryout(n12619),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i15_LC_16_18_6.C_ON=1'b1;
    defparam sweep_counter_631_632__i15_LC_16_18_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i15_LC_16_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i15_LC_16_18_6 (
            .in0(_gnd_net_),
            .in1(N__50715),
            .in2(_gnd_net_),
            .in3(N__50701),
            .lcout(sweep_counter_14),
            .ltout(),
            .carryin(n12619),
            .carryout(n12620),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i16_LC_16_18_7.C_ON=1'b1;
    defparam sweep_counter_631_632__i16_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i16_LC_16_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i16_LC_16_18_7 (
            .in0(_gnd_net_),
            .in1(N__50697),
            .in2(_gnd_net_),
            .in3(N__50683),
            .lcout(sweep_counter_15),
            .ltout(),
            .carryin(n12620),
            .carryout(n12621),
            .clk(N__56052),
            .ce(),
            .sr(N__52869));
    defparam sweep_counter_631_632__i17_LC_16_19_0.C_ON=1'b1;
    defparam sweep_counter_631_632__i17_LC_16_19_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i17_LC_16_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i17_LC_16_19_0 (
            .in0(_gnd_net_),
            .in1(N__50680),
            .in2(_gnd_net_),
            .in3(N__50668),
            .lcout(sweep_counter_16),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(n12622),
            .clk(N__56056),
            .ce(),
            .sr(N__52883));
    defparam sweep_counter_631_632__i18_LC_16_19_1.C_ON=1'b0;
    defparam sweep_counter_631_632__i18_LC_16_19_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_631_632__i18_LC_16_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_631_632__i18_LC_16_19_1 (
            .in0(_gnd_net_),
            .in1(N__50662),
            .in2(_gnd_net_),
            .in3(N__50665),
            .lcout(sweep_counter_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56056),
            .ce(),
            .sr(N__52883));
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_16_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_16_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_2_lut_LC_16_22_0 (
            .in0(_gnd_net_),
            .in1(N__51180),
            .in2(_gnd_net_),
            .in3(N__51121),
            .lcout(n3201),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(n12492),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_16_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_16_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_3_lut_LC_16_22_1 (
            .in0(_gnd_net_),
            .in1(N__54343),
            .in2(N__51118),
            .in3(N__51079),
            .lcout(n3200),
            .ltout(),
            .carryin(n12492),
            .carryout(n12493),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_16_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_16_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_16_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_4_lut_LC_16_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51076),
            .in3(N__51022),
            .lcout(n3199),
            .ltout(),
            .carryin(n12493),
            .carryout(n12494),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_16_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_16_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_16_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_5_lut_LC_16_22_3 (
            .in0(_gnd_net_),
            .in1(N__54344),
            .in2(N__51019),
            .in3(N__50986),
            .lcout(n3198),
            .ltout(),
            .carryin(n12494),
            .carryout(n12495),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_16_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_16_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_16_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_6_lut_LC_16_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50983),
            .in3(N__50932),
            .lcout(n3197),
            .ltout(),
            .carryin(n12495),
            .carryout(n12496),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_16_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_16_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_16_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_7_lut_LC_16_22_5 (
            .in0(_gnd_net_),
            .in1(N__50924),
            .in2(_gnd_net_),
            .in3(N__50881),
            .lcout(n3196),
            .ltout(),
            .carryin(n12496),
            .carryout(n12497),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_16_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_16_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_16_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_8_lut_LC_16_22_6 (
            .in0(_gnd_net_),
            .in1(N__54346),
            .in2(N__50878),
            .in3(N__50827),
            .lcout(n3195),
            .ltout(),
            .carryin(n12497),
            .carryout(n12498),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_16_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_16_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_16_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_9_lut_LC_16_22_7 (
            .in0(_gnd_net_),
            .in1(N__54345),
            .in2(N__50820),
            .in3(N__50779),
            .lcout(n3194),
            .ltout(),
            .carryin(n12498),
            .carryout(n12499),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_16_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_16_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_16_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_10_lut_LC_16_23_0 (
            .in0(_gnd_net_),
            .in1(N__54784),
            .in2(N__51555),
            .in3(N__51502),
            .lcout(n3193),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(n12500),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_16_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_16_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_16_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_11_lut_LC_16_23_1 (
            .in0(_gnd_net_),
            .in1(N__51499),
            .in2(N__55076),
            .in3(N__51451),
            .lcout(n3192),
            .ltout(),
            .carryin(n12500),
            .carryout(n12501),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_16_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_16_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_16_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_12_lut_LC_16_23_2 (
            .in0(_gnd_net_),
            .in1(N__51448),
            .in2(N__55122),
            .in3(N__51409),
            .lcout(n3191),
            .ltout(),
            .carryin(n12501),
            .carryout(n12502),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_16_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_16_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_16_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_13_lut_LC_16_23_3 (
            .in0(_gnd_net_),
            .in1(N__51405),
            .in2(N__55077),
            .in3(N__51352),
            .lcout(n3190),
            .ltout(),
            .carryin(n12502),
            .carryout(n12503),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_16_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_16_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_16_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_14_lut_LC_16_23_4 (
            .in0(_gnd_net_),
            .in1(N__51349),
            .in2(N__55123),
            .in3(N__51313),
            .lcout(n3189),
            .ltout(),
            .carryin(n12503),
            .carryout(n12504),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_16_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_16_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_16_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_15_lut_LC_16_23_5 (
            .in0(_gnd_net_),
            .in1(N__51309),
            .in2(N__55078),
            .in3(N__51277),
            .lcout(n3188),
            .ltout(),
            .carryin(n12504),
            .carryout(n12505),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_16_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_16_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_16_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_16_lut_LC_16_23_6 (
            .in0(_gnd_net_),
            .in1(N__51274),
            .in2(N__55124),
            .in3(N__51226),
            .lcout(n3187),
            .ltout(),
            .carryin(n12505),
            .carryout(n12506),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_16_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_16_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_16_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_17_lut_LC_16_23_7 (
            .in0(_gnd_net_),
            .in1(N__51223),
            .in2(N__55079),
            .in3(N__51184),
            .lcout(n3186),
            .ltout(),
            .carryin(n12506),
            .carryout(n12507),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_16_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_16_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_16_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_18_lut_LC_16_24_0 (
            .in0(_gnd_net_),
            .in1(N__51856),
            .in2(N__55080),
            .in3(N__51808),
            .lcout(n3185),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(n12508),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_16_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_16_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_16_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_19_lut_LC_16_24_1 (
            .in0(_gnd_net_),
            .in1(N__51804),
            .in2(N__55125),
            .in3(N__51760),
            .lcout(n3184),
            .ltout(),
            .carryin(n12508),
            .carryout(n12509),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_16_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_16_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_16_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_20_lut_LC_16_24_2 (
            .in0(_gnd_net_),
            .in1(N__51757),
            .in2(N__55081),
            .in3(N__51718),
            .lcout(n3183),
            .ltout(),
            .carryin(n12509),
            .carryout(n12510),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_16_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_16_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_16_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_21_lut_LC_16_24_3 (
            .in0(_gnd_net_),
            .in1(N__51711),
            .in2(N__55126),
            .in3(N__51673),
            .lcout(n3182),
            .ltout(),
            .carryin(n12510),
            .carryout(n12511),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_16_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_16_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_16_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_22_lut_LC_16_24_4 (
            .in0(_gnd_net_),
            .in1(N__51663),
            .in2(N__55082),
            .in3(N__51643),
            .lcout(n3181),
            .ltout(),
            .carryin(n12511),
            .carryout(n12512),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_16_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_16_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_16_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_23_lut_LC_16_24_5 (
            .in0(_gnd_net_),
            .in1(N__51640),
            .in2(N__55127),
            .in3(N__51595),
            .lcout(n3180),
            .ltout(),
            .carryin(n12512),
            .carryout(n12513),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_16_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_16_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_16_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_24_lut_LC_16_24_6 (
            .in0(_gnd_net_),
            .in1(N__51592),
            .in2(N__55083),
            .in3(N__51559),
            .lcout(n3179),
            .ltout(),
            .carryin(n12513),
            .carryout(n12514),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_16_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_16_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_16_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_25_lut_LC_16_24_7 (
            .in0(_gnd_net_),
            .in1(N__52225),
            .in2(N__55128),
            .in3(N__52177),
            .lcout(n3178),
            .ltout(),
            .carryin(n12514),
            .carryout(n12515),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_16_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_16_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_16_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_26_lut_LC_16_25_0 (
            .in0(_gnd_net_),
            .in1(N__52167),
            .in2(N__55129),
            .in3(N__52147),
            .lcout(n3177),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(n12516),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_16_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_16_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_16_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_27_lut_LC_16_25_1 (
            .in0(_gnd_net_),
            .in1(N__52144),
            .in2(N__55084),
            .in3(N__52096),
            .lcout(n3176),
            .ltout(),
            .carryin(n12516),
            .carryout(n12517),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_16_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_16_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_16_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_28_lut_LC_16_25_2 (
            .in0(_gnd_net_),
            .in1(N__52077),
            .in2(N__55130),
            .in3(N__52048),
            .lcout(n3175),
            .ltout(),
            .carryin(n12517),
            .carryout(n12518),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_16_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_16_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_16_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_29_lut_LC_16_25_3 (
            .in0(_gnd_net_),
            .in1(N__52045),
            .in2(N__55085),
            .in3(N__52003),
            .lcout(n3174),
            .ltout(),
            .carryin(n12518),
            .carryout(n12519),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_16_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_16_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_16_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_30_lut_LC_16_25_4 (
            .in0(_gnd_net_),
            .in1(N__52000),
            .in2(N__55131),
            .in3(N__51955),
            .lcout(n3173),
            .ltout(),
            .carryin(n12519),
            .carryout(n12520),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_16_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_16_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_16_25_5.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_2106_31_lut_LC_16_25_5 (
            .in0(N__54815),
            .in1(N__51952),
            .in2(N__51937),
            .in3(N__51913),
            .lcout(n3204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_630__i0_LC_16_26_0.C_ON=1'b1;
    defparam encoder0_position_target_630__i0_LC_16_26_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i0_LC_16_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i0_LC_16_26_0 (
            .in0(_gnd_net_),
            .in1(N__51879),
            .in2(_gnd_net_),
            .in3(N__51859),
            .lcout(encoder0_position_target_0),
            .ltout(),
            .carryin(bfn_16_26_0_),
            .carryout(n12663),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i1_LC_16_26_1.C_ON=1'b1;
    defparam encoder0_position_target_630__i1_LC_16_26_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i1_LC_16_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i1_LC_16_26_1 (
            .in0(_gnd_net_),
            .in1(N__52470),
            .in2(N__55086),
            .in3(N__52450),
            .lcout(encoder0_position_target_1),
            .ltout(),
            .carryin(n12663),
            .carryout(n12664),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i2_LC_16_26_2.C_ON=1'b1;
    defparam encoder0_position_target_630__i2_LC_16_26_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i2_LC_16_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i2_LC_16_26_2 (
            .in0(_gnd_net_),
            .in1(N__54819),
            .in2(N__52443),
            .in3(N__52417),
            .lcout(encoder0_position_target_2),
            .ltout(),
            .carryin(n12664),
            .carryout(n12665),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i3_LC_16_26_3.C_ON=1'b1;
    defparam encoder0_position_target_630__i3_LC_16_26_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i3_LC_16_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i3_LC_16_26_3 (
            .in0(_gnd_net_),
            .in1(N__52410),
            .in2(N__55087),
            .in3(N__52390),
            .lcout(encoder0_position_target_3),
            .ltout(),
            .carryin(n12665),
            .carryout(n12666),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i4_LC_16_26_4.C_ON=1'b1;
    defparam encoder0_position_target_630__i4_LC_16_26_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i4_LC_16_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i4_LC_16_26_4 (
            .in0(_gnd_net_),
            .in1(N__54823),
            .in2(N__52386),
            .in3(N__52360),
            .lcout(encoder0_position_target_4),
            .ltout(),
            .carryin(n12666),
            .carryout(n12667),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i5_LC_16_26_5.C_ON=1'b1;
    defparam encoder0_position_target_630__i5_LC_16_26_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i5_LC_16_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i5_LC_16_26_5 (
            .in0(_gnd_net_),
            .in1(N__52356),
            .in2(N__55088),
            .in3(N__52336),
            .lcout(encoder0_position_target_5),
            .ltout(),
            .carryin(n12667),
            .carryout(n12668),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i6_LC_16_26_6.C_ON=1'b1;
    defparam encoder0_position_target_630__i6_LC_16_26_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i6_LC_16_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i6_LC_16_26_6 (
            .in0(_gnd_net_),
            .in1(N__54827),
            .in2(N__52333),
            .in3(N__52309),
            .lcout(encoder0_position_target_6),
            .ltout(),
            .carryin(n12668),
            .carryout(n12669),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i7_LC_16_26_7.C_ON=1'b1;
    defparam encoder0_position_target_630__i7_LC_16_26_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i7_LC_16_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i7_LC_16_26_7 (
            .in0(_gnd_net_),
            .in1(N__52305),
            .in2(N__55089),
            .in3(N__52285),
            .lcout(encoder0_position_target_7),
            .ltout(),
            .carryin(n12669),
            .carryout(n12670),
            .clk(N__56080),
            .ce(N__52896),
            .sr(N__52827));
    defparam encoder0_position_target_630__i8_LC_16_27_0.C_ON=1'b1;
    defparam encoder0_position_target_630__i8_LC_16_27_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i8_LC_16_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i8_LC_16_27_0 (
            .in0(_gnd_net_),
            .in1(N__55102),
            .in2(N__52282),
            .in3(N__52255),
            .lcout(encoder0_position_target_8),
            .ltout(),
            .carryin(bfn_16_27_0_),
            .carryout(n12671),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i9_LC_16_27_1.C_ON=1'b1;
    defparam encoder0_position_target_630__i9_LC_16_27_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i9_LC_16_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i9_LC_16_27_1 (
            .in0(_gnd_net_),
            .in1(N__52248),
            .in2(N__55213),
            .in3(N__52228),
            .lcout(encoder0_position_target_9),
            .ltout(),
            .carryin(n12671),
            .carryout(n12672),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i10_LC_16_27_2.C_ON=1'b1;
    defparam encoder0_position_target_630__i10_LC_16_27_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i10_LC_16_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i10_LC_16_27_2 (
            .in0(_gnd_net_),
            .in1(N__55090),
            .in2(N__52702),
            .in3(N__52678),
            .lcout(encoder0_position_target_10),
            .ltout(),
            .carryin(n12672),
            .carryout(n12673),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i11_LC_16_27_3.C_ON=1'b1;
    defparam encoder0_position_target_630__i11_LC_16_27_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i11_LC_16_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i11_LC_16_27_3 (
            .in0(_gnd_net_),
            .in1(N__52674),
            .in2(N__55210),
            .in3(N__52654),
            .lcout(encoder0_position_target_11),
            .ltout(),
            .carryin(n12673),
            .carryout(n12674),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i12_LC_16_27_4.C_ON=1'b1;
    defparam encoder0_position_target_630__i12_LC_16_27_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i12_LC_16_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i12_LC_16_27_4 (
            .in0(_gnd_net_),
            .in1(N__55094),
            .in2(N__52650),
            .in3(N__52624),
            .lcout(encoder0_position_target_12),
            .ltout(),
            .carryin(n12674),
            .carryout(n12675),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i13_LC_16_27_5.C_ON=1'b1;
    defparam encoder0_position_target_630__i13_LC_16_27_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i13_LC_16_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i13_LC_16_27_5 (
            .in0(_gnd_net_),
            .in1(N__52616),
            .in2(N__55211),
            .in3(N__52594),
            .lcout(encoder0_position_target_13),
            .ltout(),
            .carryin(n12675),
            .carryout(n12676),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i14_LC_16_27_6.C_ON=1'b1;
    defparam encoder0_position_target_630__i14_LC_16_27_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i14_LC_16_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i14_LC_16_27_6 (
            .in0(_gnd_net_),
            .in1(N__55098),
            .in2(N__52590),
            .in3(N__52561),
            .lcout(encoder0_position_target_14),
            .ltout(),
            .carryin(n12676),
            .carryout(n12677),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i15_LC_16_27_7.C_ON=1'b1;
    defparam encoder0_position_target_630__i15_LC_16_27_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i15_LC_16_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i15_LC_16_27_7 (
            .in0(_gnd_net_),
            .in1(N__52554),
            .in2(N__55212),
            .in3(N__52534),
            .lcout(encoder0_position_target_15),
            .ltout(),
            .carryin(n12677),
            .carryout(n12678),
            .clk(N__56085),
            .ce(N__52897),
            .sr(N__52828));
    defparam encoder0_position_target_630__i16_LC_16_28_0.C_ON=1'b1;
    defparam encoder0_position_target_630__i16_LC_16_28_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i16_LC_16_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i16_LC_16_28_0 (
            .in0(_gnd_net_),
            .in1(N__52530),
            .in2(N__55214),
            .in3(N__52510),
            .lcout(encoder0_position_target_16),
            .ltout(),
            .carryin(bfn_16_28_0_),
            .carryout(n12679),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i17_LC_16_28_1.C_ON=1'b1;
    defparam encoder0_position_target_630__i17_LC_16_28_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i17_LC_16_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i17_LC_16_28_1 (
            .in0(_gnd_net_),
            .in1(N__55109),
            .in2(N__52503),
            .in3(N__52477),
            .lcout(encoder0_position_target_17),
            .ltout(),
            .carryin(n12679),
            .carryout(n12680),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i18_LC_16_28_2.C_ON=1'b1;
    defparam encoder0_position_target_630__i18_LC_16_28_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i18_LC_16_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i18_LC_16_28_2 (
            .in0(_gnd_net_),
            .in1(N__55392),
            .in2(N__55215),
            .in3(N__55369),
            .lcout(encoder0_position_target_18),
            .ltout(),
            .carryin(n12680),
            .carryout(n12681),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i19_LC_16_28_3.C_ON=1'b1;
    defparam encoder0_position_target_630__i19_LC_16_28_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i19_LC_16_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i19_LC_16_28_3 (
            .in0(_gnd_net_),
            .in1(N__55113),
            .in2(N__55362),
            .in3(N__55336),
            .lcout(encoder0_position_target_19),
            .ltout(),
            .carryin(n12681),
            .carryout(n12682),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i20_LC_16_28_4.C_ON=1'b1;
    defparam encoder0_position_target_630__i20_LC_16_28_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i20_LC_16_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i20_LC_16_28_4 (
            .in0(_gnd_net_),
            .in1(N__55329),
            .in2(N__55216),
            .in3(N__55309),
            .lcout(encoder0_position_target_20),
            .ltout(),
            .carryin(n12682),
            .carryout(n12683),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i21_LC_16_28_5.C_ON=1'b1;
    defparam encoder0_position_target_630__i21_LC_16_28_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i21_LC_16_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i21_LC_16_28_5 (
            .in0(_gnd_net_),
            .in1(N__55117),
            .in2(N__55305),
            .in3(N__55279),
            .lcout(encoder0_position_target_21),
            .ltout(),
            .carryin(n12683),
            .carryout(n12684),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i22_LC_16_28_6.C_ON=1'b1;
    defparam encoder0_position_target_630__i22_LC_16_28_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i22_LC_16_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_630__i22_LC_16_28_6 (
            .in0(_gnd_net_),
            .in1(N__55272),
            .in2(N__55217),
            .in3(N__55252),
            .lcout(encoder0_position_target_22),
            .ltout(),
            .carryin(n12684),
            .carryout(n12685),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam encoder0_position_target_630__i23_LC_16_28_7.C_ON=1'b0;
    defparam encoder0_position_target_630__i23_LC_16_28_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_630__i23_LC_16_28_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_target_630__i23_LC_16_28_7 (
            .in0(N__52917),
            .in1(N__55121),
            .in2(_gnd_net_),
            .in3(N__52921),
            .lcout(encoder0_position_target_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56089),
            .ce(N__52881),
            .sr(N__52823));
    defparam pwm_setpoint_i9_LC_16_29_0.C_ON=1'b0;
    defparam pwm_setpoint_i9_LC_16_29_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i9_LC_16_29_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i9_LC_16_29_0 (
            .in0(N__55706),
            .in1(N__52801),
            .in2(_gnd_net_),
            .in3(N__52792),
            .lcout(pwm_setpoint_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i9_1_lut_LC_16_29_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_16_29_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_16_29_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i9_1_lut_LC_16_29_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52731),
            .lcout(n17_adj_583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i1_LC_16_29_6.C_ON=1'b0;
    defparam commutation_state_prev_i1_LC_16_29_6.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i1_LC_16_29_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 commutation_state_prev_i1_LC_16_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56382),
            .lcout(commutation_state_prev_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam dir_151_LC_16_30_4.C_ON=1'b0;
    defparam dir_151_LC_16_30_4.SEQ_MODE=4'b1000;
    defparam dir_151_LC_16_30_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 dir_151_LC_16_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55707),
            .lcout(dir),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56094),
            .ce(),
            .sr(_gnd_net_));
    defparam i2137_1_lut_LC_17_27_0.C_ON=1'b0;
    defparam i2137_1_lut_LC_17_27_0.SEQ_MODE=4'b0000;
    defparam i2137_1_lut_LC_17_27_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i2137_1_lut_LC_17_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55695),
            .lcout(pwm_setpoint_23__N_195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_inv_0_i7_1_lut_LC_17_27_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_inv_0_i7_1_lut_LC_17_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_inv_0_i7_1_lut_LC_17_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_inv_0_i7_1_lut_LC_17_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55546),
            .lcout(n19_adj_551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3168_2_lut_LC_17_30_1.C_ON=1'b0;
    defparam i3168_2_lut_LC_17_30_1.SEQ_MODE=4'b0000;
    defparam i3168_2_lut_LC_17_30_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i3168_2_lut_LC_17_30_1 (
            .in0(_gnd_net_),
            .in1(N__55887),
            .in2(_gnd_net_),
            .in3(N__55516),
            .lcout(n4886),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12416_4_lut_LC_17_31_0.C_ON=1'b0;
    defparam i12416_4_lut_LC_17_31_0.SEQ_MODE=4'b0000;
    defparam i12416_4_lut_LC_17_31_0.LUT_INIT=16'b1101111100010011;
    LogicCell40 i12416_4_lut_LC_17_31_0 (
            .in0(N__56374),
            .in1(N__55515),
            .in2(N__56180),
            .in3(N__55471),
            .lcout(n4842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GLC_165_LC_17_31_7.C_ON=1'b0;
    defparam GLC_165_LC_17_31_7.SEQ_MODE=4'b1000;
    defparam GLC_165_LC_17_31_7.LUT_INIT=16'b0101110000101100;
    LogicCell40 GLC_165_LC_17_31_7 (
            .in0(N__56301),
            .in1(N__56165),
            .in2(N__56434),
            .in3(N__56375),
            .lcout(INLC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56095),
            .ce(N__55900),
            .sr(N__55855));
    defparam GLA_161_LC_18_31_7.C_ON=1'b0;
    defparam GLA_161_LC_18_31_7.SEQ_MODE=4'b1000;
    defparam GLA_161_LC_18_31_7.LUT_INIT=16'b1001100000000011;
    LogicCell40 GLA_161_LC_18_31_7 (
            .in0(N__56296),
            .in1(N__56376),
            .in2(N__56194),
            .in3(N__56437),
            .lcout(INLA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56096),
            .ce(N__55901),
            .sr(N__55859));
    defparam GHB_162_LC_19_30_0.C_ON=1'b0;
    defparam GHB_162_LC_19_30_0.SEQ_MODE=4'b1000;
    defparam GHB_162_LC_19_30_0.LUT_INIT=16'b1100110000100001;
    LogicCell40 GHB_162_LC_19_30_0 (
            .in0(N__56294),
            .in1(N__56389),
            .in2(N__56196),
            .in3(N__56429),
            .lcout(GHB),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56097),
            .ce(N__55912),
            .sr(N__55864));
    defparam GHC_164_LC_19_30_4.C_ON=1'b0;
    defparam GHC_164_LC_19_30_4.SEQ_MODE=4'b1000;
    defparam GHC_164_LC_19_30_4.LUT_INIT=16'b1111000001000110;
    LogicCell40 GHC_164_LC_19_30_4 (
            .in0(N__56295),
            .in1(N__56390),
            .in2(N__56197),
            .in3(N__56430),
            .lcout(GHC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56097),
            .ce(N__55912),
            .sr(N__55864));
    defparam GLB_163_LC_19_31_3.C_ON=1'b0;
    defparam GLB_163_LC_19_31_3.SEQ_MODE=4'b1000;
    defparam GLB_163_LC_19_31_3.LUT_INIT=16'b0110001000100110;
    LogicCell40 GLB_163_LC_19_31_3 (
            .in0(N__56391),
            .in1(N__56436),
            .in2(N__56195),
            .in3(N__56300),
            .lcout(INLB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56098),
            .ce(N__55908),
            .sr(N__55860));
    defparam GHA_160_LC_19_31_6.C_ON=1'b0;
    defparam GHA_160_LC_19_31_6.SEQ_MODE=4'b1000;
    defparam GHA_160_LC_19_31_6.LUT_INIT=16'b0100000101100010;
    LogicCell40 GHA_160_LC_19_31_6 (
            .in0(N__56435),
            .in1(N__56392),
            .in2(N__56302),
            .in3(N__56187),
            .lcout(GHA),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56098),
            .ce(N__55908),
            .sr(N__55860));
    defparam i9555_2_lut_LC_19_32_6.C_ON=1'b0;
    defparam i9555_2_lut_LC_19_32_6.SEQ_MODE=4'b0000;
    defparam i9555_2_lut_LC_19_32_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9555_2_lut_LC_19_32_6 (
            .in0(N__55816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55771),
            .lcout(INHA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9489_2_lut_LC_20_30_0.C_ON=1'b0;
    defparam i9489_2_lut_LC_20_30_0.SEQ_MODE=4'b0000;
    defparam i9489_2_lut_LC_20_30_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9489_2_lut_LC_20_30_0 (
            .in0(N__55767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55795),
            .lcout(INHC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9488_2_lut_LC_20_30_7.C_ON=1'b0;
    defparam i9488_2_lut_LC_20_30_7.SEQ_MODE=4'b0000;
    defparam i9488_2_lut_LC_20_30_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9488_2_lut_LC_20_30_7 (
            .in0(N__55777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55766),
            .lcout(INHB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
