// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Mar  9 10:47:44 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, n861, 
        GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    
    wire n52116, n52115, n51636;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n60859, n52114;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n52113, n51635, data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(363[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(371[15:20])
    
    wire pwm_setpoint_23__N_255, n209, n211, n52112, n60700, n26490, 
        n249, n250, n251, n252, n253, n254, n255, n256, n257, 
        n258, n259, n260, n261, n262, n263, n264, n265, n266, 
        n267, n268, n269, n270, n51634, n296, n10, n10_adj_5842, 
        n9, n8, n330, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345, n7;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n356, n70963, n70957, n70951, n70945, n379, n59065, n6196, 
        n418, n419, n420, n421, n422, n423, n424, n425, n426, 
        n427, n428, n429, n430, n431, n432, n433, n434, n435, 
        n436, n437, n438, n439, n440, n441, n67742, n51633;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n29784, n51321, n25959;
    wire [7:0]commutation_state_7__N_256;
    
    wire n51632, commutation_state_7__N_264;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n28507, GHA_N_468, GLA_N_485, GHB_N_490, GLB_N_499, GHC_N_504, 
        GLC_N_513, dti_N_517, RX_N_2;
    wire [31:0]motor_state_23__N_115;
    wire [31:0]encoder0_position_scaled_23__N_319;
    wire [32:0]encoder0_position_scaled_23__N_43;
    
    wire encoder1_position_scaled_23__N_351;
    wire [31:0]encoder1_position_scaled_23__N_67;
    wire [23:0]displacement_23__N_91;
    
    wire n52111, n2275, n833, n832, n831, n830, n829, n828, 
        n7903, n7904, n7905, n7906, n7907, n7908, n8_adj_5843, 
        n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
        n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
        n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
        n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
        read_N_522, n1642, n52110, n52109, n51631, n52108, n24, 
        n69639, n19, n17, n16, n15, n13, n11, n9_adj_5844, n8_adj_5845, 
        n7_adj_5846, n6, n5, n4, n2092, n2234;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[11:16])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n60713, n5439, n5438, n6_adj_5847, n5437, n5436, n5435, 
        n5434, n5433, n15_adj_5848, n23298, n52107, n5431, n5430, 
        n5429, n5428, n5427, n51630, n5426, n44625, n5425, n5424, 
        n5423, n5422, n49984, n51792, n51629, n51628, n40, n51791, 
        n52106, n3, n4_adj_5849, n5_adj_5850, n6_adj_5851, n7_adj_5852, 
        n8_adj_5853, n9_adj_5854, n10_adj_5855, n11_adj_5856, n12, 
        n13_adj_5857, n14, n15_adj_5858, n16_adj_5859, n17_adj_5860, 
        n18, n19_adj_5861, n20, n21, n22, n23, n24_adj_5862, n2, 
        n51790, n14_adj_5863, n15_adj_5864, n16_adj_5865, n17_adj_5866, 
        n18_adj_5867, n19_adj_5868, n20_adj_5869, n21_adj_5870, n22_adj_5871, 
        n23_adj_5872, n24_adj_5873, n25, n6_adj_5874, n37022, n52105, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active, n52104, n5_adj_5875, n51789;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n4_adj_5876, n3_adj_5877, 
        n51788, n51787, n3305, n51627, n2_adj_5878, n52103, n51626, 
        n52102, n51391, n3358, n52101, n63662, n52100, n52099, 
        n51390, n51320, n52098, n43, n51625, n51624, n51623, n51389, 
        n51622, n58976, n58975, n58974, n58973, n58972, n58971, 
        n58970, n58969, n58968, n58967, n58966, n58965, n58964, 
        n58963, n58962, n58961, n58960, n58959, n58826, n58958, 
        n58957, n58956, n58955, n58954, n58953, n58952, n58951, 
        n58950, n58949, n58948, n58947, n58946, n58945, n58944, 
        n58943, n58942, n58941, n58940, n58939, n58938, n58937, 
        n58936, n58935, n58934, n58933, n58932, n58931, n58930, 
        n58929, n58928, n58927, n58926, n58827, n58925, n58924, 
        n58923, n58922, n58921, n58920, n58919, n58918, n58917, 
        n58916, n58915, n58914, n58913, n58912, n58911, n58910, 
        n58909, n58908, n58907, n58906, n58905, n58904, n58903, 
        n58902, n58901, n58900, n58830, n58833, n58834, n58835, 
        n58836, n58837, n58842, n58844, n58848, n58849, n58850, 
        n58845, n58851, n58852, n58847, n58853, n58854, n58855, 
        n58856, n58857, n58858, n58859, n58828, n58860, n58861, 
        n58862, n58863, n58864, n58865, n58866, n29319, n29318, 
        n29317, n58867, n58868, n58869, n58870, n58871, n29311, 
        n58872, n58873, n58874, n58875, n58876, n58877, n58878, 
        n58879, n58839, n58880, n58838, n58882, n58883, n58884, 
        n58832, n58831, n58886, n58887, n58888, n58889, n58890, 
        n58891, n58892, n58893, n58894, n29283, n58896, n29256, 
        n29255, n29254, n58825, n29251, n58897, n58898, n58829, 
        n63656, n14_adj_5879, n13_adj_5880, n12_adj_5881, n63650, 
        n51786, n51785, n63644, n51621, n51784, n52097, n51783, 
        n51782, n63642, n51620, n51619, n51618, n51617, n52096, 
        n52095, n51616, n51615, n51388, n51387, n52094, n52093, 
        n51614, n51613, n51612, n52092, n51611, n51610, n52091, 
        n51609, n51386, n52090, n51608, n52089, n51607, n51385, 
        n52088, n52087, n52086, n52085, n51767, n52084, n51766, 
        n51337, n52083, n51384, n62, n52082, n51765, n52081, n51383, 
        n51764, n52080, n51763, n51762, n52079, n51382, n51761, 
        n51760, n51759, n63628, n52078, n52077, n51336, n51381, 
        n51758, n63626, n52076, n52075, n52074, n51335, n52073, 
        n51380, n51379, n43962, n51378, n52072, n51319, n52071, 
        n63624, n51377, n52070, n51376, n53140, n53139, n53138, 
        n43842, n63618, n63614, n5421, n63606, n70939, n70933, 
        n11_adj_5882, n5257, n63600, n63598, n70125, n63892, n67674, 
        n51375, n5254, n5246, n61411, n60053, n63566, n63562, 
        n26087, n63556, n63554, n60009, n59994, n63540, n53137, 
        n63534, n6_adj_5883, \FRAME_MATCHER.i_31__N_2638 , n59975, n26, 
        n19_adj_5884, n17_adj_5885, n16_adj_5886, n15_adj_5887, n69353, 
        n13_adj_5888, n11_adj_5889, n9_adj_5890, n8_adj_5891, n7_adj_5892, 
        n6_adj_5893, n5_adj_5894, n4_adj_5895, n59971, n44799, n30260, 
        n30257, n30256, n30255, n30254, n30253, n30252, n30250, 
        n30249, n30248, n30247, n30246, n30245, n30244, n30243, 
        n30242, n30241, n30240, n30239, n30238, n30237, n30236, 
        n30235, n30234, n30233, n30232, n30231, n44797, n44695, 
        n30228, n44795, n58881, n30225, n30222, n30219, n30216, 
        n44787, n30208, n30207, n30130, n30129, n30128, n30127, 
        n30126, n30125, n30124, n30123, n30121, n57536, n44781, 
        n44779, n30090, n30075, n30074, n30073, n30072, n30068, 
        n30067, n30066, n44777, n30062, n30061, n30060, n30059, 
        n30058, n30057, n30054, n44775, n30049, n30047, n44773, 
        n30042, n30041, n30035, n30034, n63528, n30031, n30028, 
        n30025, n30024, n30023, n44771, n30016, n30015, n30014, 
        n30013, n30012, n30010, n44767, n30003, n29995, n44765, 
        n29992, n29989, n29986, n29983, n29980, n29977, n53136, 
        n29968, n29964, n53135, n29961, n29958, n63526, n29952, 
        n29949, n58226, n58228, n58230, n29921, n29912, n29909, 
        n44831, n44827, n44823, n29867, n29861, n32, n24_adj_5896, 
        n17_adj_5897, n15_adj_5898, n14_adj_5899, n13_adj_5900, n11_adj_5901, 
        n53134, n4_adj_5902, n67659, n9_adj_5903, n70372, n7_adj_5904, 
        n6_adj_5905, n5_adj_5906, n4_adj_5907, n53133, n51738, n31166, 
        n51737, n31164, n63512, n8_adj_5908, n31163, n31162, n58824, 
        n51736, n51735, n15_adj_5909, n51734, n4_adj_5910, n63506, 
        n4_adj_5911, n31082, n31075, n31074, n25984, n63504, n11_adj_5912, 
        n11_adj_5913, n63498, n6_adj_5914, n63490, n44803, n6_adj_5915, 
        n30855, n30854, n15_adj_5916, n652, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n30850, n60079, n30847, n63484, n53132, n30842, n30841, 
        n25_adj_5917, n24_adj_5918, n23_adj_5919, n22_adj_5920, n21_adj_5921, 
        n20_adj_5922, n19_adj_5923, n18_adj_5924, n17_adj_5925, n16_adj_5926, 
        n58352, n136, n149, n155, n181, n188, n219;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3844 ;
    
    wire n379_adj_5927, n70927, n405, n30828, n30827, n30826, n11_adj_5928, 
        n30825, n30824, n30823, n30822, n30821, n30820, n30819, 
        n30818, n30817, n30816, n30815, n30814, n30813, n30812, 
        n30811, n30810, n30809, n30808, n30807, n30806, n30805, 
        n30804, n30803, n30802, n30801;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, n30800, n30799, n30798, n30797, position_31__N_3956, 
        n625, n623, n622, n621, n51733, n51732, n53131, n63478, 
        n5420, n5419, n5418, n5417, n5416, n5415, n5414, n5413, 
        n5412, n5411, n5409, n15_adj_5929, n30796, n30795, n30794, 
        n30793, n30792, n30791, n30790, n25840;
    wire [1:0]a_new_adj_6125;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5931, position_31__N_3956_adj_5932, n53130, n63476, 
        n53129, n519, n518, n59887, n516, n53128, n59885, n59883, 
        n59881, n59878, n30773, n30772, n30771, n15_adj_5933, n30770, 
        n63470, n30769, n30768, n53127, n63466, n30767, n30766;
    wire [7:0]data_adj_6138;   // verilog/eeprom.v(23[12:16])
    
    wire ready_prev, n30765, rw;
    wire [7:0]state_adj_6139;   // verilog/eeprom.v(27[11:16])
    wire [7:0]state_7__N_4045;
    
    wire n30763, n63462, n30761, n30760, n8_adj_5936, n30759, n30758, 
        n30757, n30756, n30755, n30754, n33, n32_adj_5937, n31, 
        n30, n54986, n58274, n29, n28, n70921, n30753, n30752, 
        n30751, n30750, n30749, n27, n7082, n26_adj_5938, n25_adj_5939, 
        n24_adj_5940, n23_adj_5941, n22_adj_5942, n30744, n5456, n5454, 
        n5453, n5452, n21_adj_5943, n20_adj_5944, n19_adj_5945, n18_adj_5946, 
        n17_adj_5947, n16_adj_5948, n30742, n15_adj_5949, n14_adj_5950, 
        n13_adj_5951, n12_adj_5952, n11_adj_5953, n10_adj_5954, n9_adj_5955, 
        n8_adj_5956, n7_adj_5957, n6_adj_5958, n5_adj_5959, n4_adj_5960, 
        n3_adj_5961, n2_adj_5962, n30710, n30707, n30706, n30705, 
        n30703, n30702, n53126, n5451, clk_out;
    wire [15:0]data_adj_6147;   // verilog/tli4970.v(27[14:18])
    
    wire n63450;
    wire [7:0]state_adj_6149;   // verilog/tli4970.v(29[13:18])
    
    wire n30693, n30690, n63446, n30677, n30674, n30672, n53125, 
        n5450, n5449, n5448, n5447, n5446, n5445, n5444, n5443, 
        n5442, n5441, n5440, state_7__N_4446, n30669, n63440, n30664, 
        n8_adj_5973, n63430, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n51731, n63428, n30639, n30638, n63422, n44815;
    wire [24:0]o_Rx_DV_N_3617;
    
    wire n70915, n30616;
    wire [2:0]r_SM_Main_adj_6161;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_6162;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_6163;   // verilog/uart_tx.v(34[16:27])
    
    wire n34987, n51730, n58899, n23164, n44755, n30587;
    wire [7:0]state_adj_6170;   // verilog/i2c_controller.v(33[12:17])
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire enable_slow_N_4340, n53124;
    wire [7:0]state_7__N_4237;
    
    wire n30566, n44805, n30562, n53123, n1, n52047, n6878;
    wire [7:0]state_7__N_4253;
    
    wire n30558, n30554, n30550, n30539, n37023, n53122, n29_adj_5988, 
        n58296, n52046, n896, n897, n898, n899, n900, n901, 
        n51, n42182, n60, n64453, n42166, n927, n928, n929, 
        n930, n931, n932, n933, n934, n935, n936, n937, n938, 
        n939, n940, n941, n942, n943, n944, n945, n946, n947, 
        n948, n949, n950, n951, n952, n953, n954, n955, n956, 
        n957, n960, n70897, n995, n996, n997, n998, n999, n1000, 
        n1001, n27_adj_5989, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1059, n23_adj_5990, n60745, n1093, 
        n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
        n53121, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
        n1132, n1133, n52045, n52044, n52043, n52866, n1158, n52865, 
        n69235, n52042, n52041, n52864, n52040, n52039, n53120, 
        n53119, n52863, n1193, n1194, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n52862, n52038, n52037, n52036, n52035, 
        n52861, n53118, n52034, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1233, n52860, n52033, n52859, 
        n52032, n53117, n53116, n52858, n1257, n52857, n52856, 
        n52031, n52030, n53115, n53114, n52855, n52854, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
        n1301, n53113, n52853, n53112, n53111, n53110, n52852, 
        n52851, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
        n1330, n1331, n1332, n1333, n52850, n52849, n52848, n1356, 
        n52847, n52846, n52845, n52844, n52843, n52842, n52841, 
        n52840, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
        n1397, n1398, n1399, n1400, n1401, n52839, n52838, n52837, 
        n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
        n1430, n1431, n1432, n1433, n52836, n1455, n1490, n1491, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531_adj_5991, n1532_adj_5992, 
        n1533_adj_5993, n1554_adj_5994, n51374, n51334, n70891, n1589, 
        n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
        n1598, n1599, n1600, n1601, n52008, n52007, n52387, n52386, 
        n52385, n52006, n52384, n1620, n1621, n1622, n1623, n1624, 
        n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
        n1633, n52005, n52383, n52382, n52381, n52380, n1653, 
        n52004, n52003, n52379, n52002, n52001, n52378, n52377, 
        n52000, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
        n1695, n1696, n1697, n1698, n1699, n1700, n1701, n51999, 
        n52376, n52375, n51717, n52374, n51998, n51997, n52373, 
        n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n52372, 
        n52371, n51716, n51333, n52370, n52369, n51996, n51715, 
        n51995, n52368, n52367, n1752, n51994, n51993, n51714, 
        n52366, n52365, n51373, n52364, n51992, n1787, n1788, 
        n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
        n1797, n1798, n1799, n1800, n1801, n52363, n52362, n52361, 
        n52360, n51713, n52359, n1818, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n51712, n52358, n1851, n52357, n52356, 
        n52355, n52354, n52353, n52352, n52351, n1886, n1887, 
        n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
        n1896, n1897, n1898, n1899, n1900, n1901, n52350, n52349, 
        n52348, n51711, n52347, n51710, n1917, n1918, n1919, n1920, 
        n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
        n1929, n1930, n1931, n1932, n1933, n52346, n52345, n52344, 
        n52343, n51412, n1950, n52342, n52341, n51971, n52340, 
        n51372, n51332, n51411, n51410, n51409, n52339, n70885, 
        n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
        n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
        n2001, n51408, n51371, n52338, n51970, n51370, n51969, 
        n52337, n52336, n2016, n2017, n2018, n2019, n2020, n2021, 
        n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n51318, n51369, n52335, n51968, 
        n51967, n52334, n52333, n2049, n52332, n51966, n51965, 
        n52331, n52330, n51964, n52329, n52328, n52327, n52326, 
        n51963, n52325, n2084, n2085, n2086, n2087, n2088, n2089, 
        n2090, n2091, n2092_adj_5995, n2093, n2094, n2095, n2096, 
        n2097, n2098, n2099, n2100, n2101, n52324, n51407, n52323, 
        n52322, n51406, n51962, n51961, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n52321, 
        n51960, n52320, n51959, n52319, n70464, n2148, n52318, 
        n51958, n51957, n52317, n51956, n51405, n51404, n52316, 
        n52315, n52314, n2182, n2183, n2184, n2185, n2186, n2187, 
        n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
        n2196, n2197, n2198, n2199, n2200, n2201, n52313, n52312, 
        n52311, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
        n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
        n2229, n2230, n2231, n2232, n2233, n52310, n52309, n2247, 
        n52308, n52307, n52306, n52305, n52304, n52303, n52302, 
        n52301, n51403, n2282, n2283, n2284, n2285, n2286, n2287, 
        n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
        n2296, n2297, n2298, n2299, n2300, n2301, n52300, n2313, 
        n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, 
        n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
        n2330, n2331, n2332, n2333, n52299, n52298, n52297, n51402, 
        n52296, n52295, n2346, n52294, n51317, n52293, n52292, 
        n52291, n51401, n2381, n2382, n2383, n2384, n2385, n2386, 
        n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
        n2395, n2396, n2397, n2398, n2399, n2400, n2401, n52290, 
        n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
        n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
        n2428, n2429, n2430, n2431, n2432, n2433, n52289, n52288, 
        n52287, n52286, n2445, n52285, n52284, n52283, n52282, 
        n52281, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
        n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
        n2495, n2496, n2497, n2498, n2499, n2500, n2501, n52280, 
        n52279, n52278, n2511, n2512, n2513, n2514, n2515, n2516, 
        n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
        n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
        n2533, n52277, n52276, n2544, n51400, n52275, n52274, 
        n52273, n51368, n52272, n52271, n51927, n52270, n52269, 
        n51926, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
        n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
        n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
        n51925, n51399, n51367, n52268, n52267, n2610, n2611, 
        n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
        n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
        n2628, n2629, n2630, n2631, n2632, n2633, n51924, n51923, 
        n2643, n51398, n52266, n51922, n52265, n52264, n52263, 
        n51921, n51920, n51366, n52262, n52261, n52260, n51693, 
        n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
        n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
        n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
        n2701, n51919, n52259, n52258, n51918, n2709, n2710, n2711, 
        n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
        n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
        n2728, n2729, n2730, n2731, n2732, n2733, n51692, n44006, 
        n2742, n52257, n2777, n2778, n2779, n2780, n2781, n2782, 
        n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
        n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
        n2799, n2800, n2801, n2808, n2809, n2810, n2811, n2812, 
        n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
        n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
        n2829, n2830, n2831, n2832, n2833, n70294, n2841, n2875, 
        n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
        n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
        n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
        n2900, n2901, n2907, n2908, n2909, n2910, n2911, n2912, 
        n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
        n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2929, n2930, n2931, n2932, n2933, n70182, n2940, n51917, 
        n43986, n51397, n51916, n52256, n2975, n2976, n2977, n2978, 
        n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
        n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
        n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3006, 
        n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
        n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
        n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
        n3031, n3032, n3033, n3039, n68222, n40932, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3138, 
        n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
        n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
        n3197, n3198, n3199, n3200, n3201, n3204, n3205, n3206, 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3233, n70130, n3237, n3271, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
        n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, 
        n3299, n3300, n3301, n58895, n61238, n51915, n52255, n52254, 
        n24_adj_5996, n62_adj_5997, n51914, n60932, n63356, n63350, 
        n25863, n63344, n64452, n51913, n28324, n28320, n70582, 
        n69347, n52253, n44807, n63334, n52252, n44717, n51396, 
        n52251, n44719, n30515, n30512, n30509, n63328, n63326, 
        n68130, n28182, n30499, n52250, n51365, n30495, n30492, 
        n51395, n52249, n51394, n52248, n28127, n52247, n51364, 
        n63318, n30489, n68124, n58524, n28109, n52246, n51363, 
        n52245, n68122, n28100, n30485, n52244, n52243, n12_adj_5998, 
        n52242, n52241, n52240, n51691, n63312, n52239, n52238, 
        n51690, n52237, n51689, n52236, n52235, n52234, n63308, 
        n52233, n30482, n52232, n28059, n52231, n51688, n11_adj_5999, 
        n37, n4_adj_6000, n69181, n30479, n63302, n30475, n28033, 
        n4_adj_6001, n6_adj_6002, n8_adj_6003, n9_adj_6004, n11_adj_6005, 
        n13_adj_6006, n15_adj_6007, n4_adj_6008, n63298, n52230, n51687, 
        n51686, n52229, n51685, n63292, n20576, n52228, n52227, 
        n20577, n52226, n20625, n52225, n52224, n52223, n52222, 
        n52221, n61039, n71059, n51684, n51393, n63278, n52220, 
        n52219, n51683, n63272, n20626, n52218, n52217, n51682, 
        n51681, n69346, n52216, n63264, n52215, n63258, n51680, 
        n52214, n63250, n52213, n63248, n52212, n63244, n63238, 
        n70642, n52211, n63232, n110, n70864, n59138, n52210, 
        n52209, n38, n56, n63222, n25605, n63216, n63210, n28_adj_6009, 
        n63204, n63198, n63194, n63192, n23230, n63180, n63178, 
        n25977, n6_adj_6010, n63176, n63174, n70861, n63172, n52208, 
        n52207, n63170, n63168, n63166, n63164, n63162, n63160, 
        n51679, n52206, n52205, n63156, n51678, n51894, n63154, 
        n51362, n63150, n70089, n51893, n52204, n63142, n63140, 
        n63138, n63136, n63134, n51892, n51891, n63132, n63126, 
        n63120, n70629, n52203, n63116, n4_adj_6011, n6_adj_6012, 
        n8_adj_6013, n9_adj_6014, n51890, n51677, n51392, n52202, 
        n51889, n52201, n52200, n38_adj_6015, n39, n40_adj_6016, 
        n41, n42, n43_adj_6017, n44, n45, n29833, n51331, n11999, 
        n51888, n52199, n51676, n52198, n51887, n51361, n71047, 
        n52197, n52196, n63104, n51886, n63794, n63098, n29536, 
        n63092, n69827, n63086, n63080, n29464, n58846, n59004, 
        n59003, n59002, n59001, n59000, n58999, n58998, n58997, 
        n58996, n58843, n58995, n58994, n58993, n58992, n58991, 
        n58990, n58989, n58988, n58987, n58986, n58841, n58840, 
        n58985, n58984, n70290, n59086, n59079, n28801, n28791, 
        n28780, n28778, n28774, n28772, n28770, n28768, n28733, 
        n29221, n28725, n28723, n28719, n28717, n63074, n67833, 
        n26902, n63068, n51885, n51360, n52195, n52194, n51884, 
        n51883, n63062, n52193, n52192, n52191, n51882, n51881, 
        n67821, n51316, n67819, n52190, n60788, n30469, n63056, 
        n51359, n51358, n51357, n69352, n57856, n52189, n30466, 
        n30465, n52188, n51356, n52187, n71041, n63050, n51330, 
        n4_adj_6018, n63048, n60705, n63046, n67789, n64056, n52186, 
        n62060, n51355, n44869, n30413, n30409, n30406, n30403, 
        n30399, n52185, n51354, n63034, n51329, n51328, n44859, 
        n30387, n44857, n30381, n44855, n30378, n52184, n58983, 
        n51353, n63028, n30375, n44851, n30371, n30368, n30365, 
        n30361, n30352, n30348, n63022, n58982, n29813, n67770, 
        n67768, n30342, n44839, n30338, n25966, n52183, n60777, 
        n63012, n29791, n52182, n52181, n52180, n52179, n63006, 
        n51665, n52178, n52177, n51664, n52176, n52175, n63000, 
        n52174, n51663, n51662, n52173, n52172, n51661, n2_adj_6019, 
        n3_adj_6020, n4_adj_6021, n5_adj_6022, n6_adj_6023, n7_adj_6024, 
        n8_adj_6025, n9_adj_6026, n10_adj_6027, n11_adj_6028, n12_adj_6029, 
        n13_adj_6030, n14_adj_6031, n15_adj_6032, n16_adj_6033, n17_adj_6034, 
        n18_adj_6035, n19_adj_6036, n20_adj_6037, n21_adj_6038, n22_adj_6039, 
        n23_adj_6040, n24_adj_6041, n25_adj_6042, n26_adj_6043, n27_adj_6044, 
        n28_adj_6045, n29_adj_6046, n30_adj_6047, n31_adj_6048, n32_adj_6049, 
        n33_adj_6050, n52171, n51660, n51352, n51351, n51273, n52170, 
        n51659, n52169, n52168, n51327, n51658, n51326, n51350, 
        n52167, n52166, n52631, n52165, n67130, n52164, n52163, 
        n51349, n51657, n52162, n52630, n51855, n52161, n52629, 
        n52628, n51854, n51853, n52160, n52627, n52626, n51852, 
        n52625, n51851, n52159, n51656, n52158, n59879, n52157, 
        n51655, n51850, n5_adj_6051, n51849, n52156, n6_adj_6052, 
        n52155, n51848, n51654, n51847, n52154, n51348, n52153, 
        n4_adj_6053, n51846, n51347, n51845, n52152, n51315, n51844, 
        n51843, n52151, n51346, n51345, n52150, n51653, n51652, 
        n52149, n52148, n51651, n52147, n51650, n67126, n67746, 
        n52146, n52145, n52144, n51649, n51648, n52143, n52142, 
        n52141, n51647, n52140, n51344, n71035, n51343, n52139, 
        n52138, n52137, n51826, n52136, n51646, n51325, n52135, 
        n51825, n51324, n52134, n52133, n51824, n51823, n52132, 
        n51822, n51821, n51820, n51342, n51819, n51645, n52131, 
        n52130, n51818, n51817, n51816, n51815, n51644, n51643, 
        n52129, n52128, n3_adj_6054, n52127, n51323, n52126, n51642, 
        n52125, n51341, n34970, n51322, n9_adj_6055, n51641, n51640, 
        n51639, n52124, n52123, n52122, n13_adj_6056, n17_adj_6057, 
        n23_adj_6058, n25_adj_6059, n27_adj_6060, n33_adj_6061, n37_adj_6062, 
        n41_adj_6063, n69906, n70570, n67082, n67080, n29783, n62864, 
        n52121, n7_adj_6064, n51340, n52120, n58885, n67072, n67070, 
        n62846, n71029, n67067, n69236, n51638, n70055, n64451, 
        n58981, n58980, n58979, n51339, n51314, n52119, n70259, 
        n10_adj_6065, n51338, n52118, n58978, n54003, n62828, n25860, 
        n70548, n51637, n35592, n67059, n55126, n62812, n52117, 
        n25975, n70321, n25971, n58977, n62796, n71023, n70527, 
        n70489, n64193, n8_adj_6066, n7_adj_6067, n64052, n70229, 
        n6_adj_6068, n71017, n25956, n62780, n62764, n62748, n69848, 
        n69847, n69763, n69840, n69839, n69828, n67030, n5_adj_6069, 
        n69659, n59967, n17_adj_6070, n25_adj_6071, n24_adj_6072, 
        n69616, n57618, n71011, n63736, n14_adj_6073, n69615, n69523, 
        n13_adj_6074, n61445, n62100, n69637, n63730, n69351, n69350, 
        n63724, n61350, n59067, n6_adj_6075, n5_adj_6076, n70460, 
        n63718, n63714, n60797, n61284, n61279, n61267, n61264, 
        n15_adj_6077, n70178, n63704, n24_adj_6078, n63698, n20_adj_6079, 
        n62584, n62091, n61896, n62578, n60803, n78, n63692, n63688, 
        n60781, n63682, n63680, n63678, n14_adj_6080, n71005, n70433, 
        n60702, n68554, n14_adj_6081, n10_adj_6082, n4_adj_6083, n69755, 
        n67754, n58198, n58202, n58208, n58212, n58216, n61347, 
        n58220, n58224, n62253, n58234, n58238, n62248, n60718, 
        n58244, n58248, n58252, n60850, n58256, n58260, n58264, 
        n58268, n58272, n58278, n58282, n58286, n58290, n58294, 
        n15_adj_6084, n9_adj_6085, n14_adj_6086, n58340, n59593, n59011, 
        n8_adj_6087, n12_adj_6088, n58384, n58398, n61440, n69908, 
        n64201, n59499, n6_adj_6089, n71131, n70999, n66923, n70993, 
        n70401, n62096, n60768, n59093, n66915, n58604, n70599, 
        n66911, n58640, n70691, n60806, n6_adj_6090, n70987;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dir_206 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_255));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_208 (.Q(dti), .C(clk16MHz), .E(n28033), .D(dti_N_517));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5848));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_6_lut (.I0(GND_net), 
            .I1(n3030), .I2(GND_net), .I3(n52280), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_6_lut (.I0(GND_net), 
            .I1(n1730), .I2(GND_net), .I3(n51916), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[0]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_91[0]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4253[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.n29783(n29783), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .clk16MHz(clk16MHz), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .GND_net(GND_net), .n40932(n40932), .neopxl_color({neopxl_color}), 
            .timer({timer}), .n30237(n30237), .n30236(n30236), .n30235(n30235), 
            .n30234(n30234), .n30233(n30233), .n30232(n30232), .VCC_net(VCC_net), 
            .n30231(n30231), .\state[0] (state[0]), .\state[1] (state[1]), 
            .n43(n43), .n30014(n30014), .n30013(n30013), .n57856(n57856), 
            .start(start), .n29784(n29784), .NEOPXL_c(NEOPXL_c), .LED_c(LED_c), 
            .n78(n78)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_7_lut (.I0(GND_net), 
            .I1(n929), .I2(GND_net), .I3(n51691), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_5_lut (.I0(GND_net), 
            .I1(n2731), .I2(VCC_net), .I3(n52201), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_6 (.CI(n52280), 
            .I0(n3030), .I1(GND_net), .CO(n52281));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_32 (.CI(n52363), 
            .I0(n3205), .I1(VCC_net), .CO(n52364));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_3_lut (.I0(GND_net), 
            .I1(n2233), .I2(VCC_net), .I3(n52089), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_3 (.CI(n52089), 
            .I0(n2233), .I1(VCC_net), .CO(n52090));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_31_lut (.I0(GND_net), 
            .I1(n3206), .I2(VCC_net), .I3(n52362), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5853));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5852));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_1_lut (.I0(current[15]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5851));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n5257), .I1(r_SM_Main_adj_6161[0]), .I2(GND_net), 
            .I3(GND_net), .O(n62578));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut (.I0(n29_adj_5988), .I1(n23_adj_5990), .I2(o_Rx_DV_N_3617[12]), 
            .I3(n62578), .O(n62584));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mux_1123_i1_4_lut (.I0(n66911), .I1(duty[0]), .I2(n296), .I3(n356), 
            .O(n5456));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam mux_1123_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1043_3_lut (.I0(n1528), 
            .I1(n1595), .I2(n1554_adj_5994), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut (.I0(n11999), .I1(n418), .I2(current[15]), 
            .I3(duty[23]), .O(n71059));
    defparam n11999_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71059_bdd_3_lut (.I0(n71059), .I1(duty[23]), .I2(n249), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam n71059_bdd_3_lut.LUT_INIT = 16'h9898;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1110_3_lut (.I0(n1627), 
            .I1(n1694), .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i8_3_lut (.I0(encoder0_position_scaled_23__N_319[7]), 
            .I1(n26_adj_5938), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1864_3_lut (.I0(n2733), 
            .I1(n2800), .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n1929), .I1(n44779), .I2(n1930), .I3(n1931), 
            .O(n60745));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2133_3_lut (.I0(n3130), 
            .I1(n3197), .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1037_3_lut (.I0(n1522), 
            .I1(n1589), .I2(n1554_adj_5994), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1748 (.I0(n296), .I1(duty[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_6055));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_2_lut_adj_1748.LUT_INIT = 16'h2222;
    SB_LUT4 i30224_2_lut (.I0(duty[2]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5454));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30224_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1177_3_lut (.I0(n1726), 
            .I1(n1793), .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n1925), .I1(n1926), .I2(n1928), .I3(n1927), 
            .O(n63022));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5850));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30223_2_lut (.I0(duty[3]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5453));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30223_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1244_3_lut (.I0(n1825), 
            .I1(n1892), .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1104_3_lut (.I0(n1621), 
            .I1(n1688), .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5849));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30222_2_lut (.I0(duty[4]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5452));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30222_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1171_3_lut (.I0(n1720), 
            .I1(n1787), .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_282_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_115[4]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5879));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_31 (.CI(n52362), 
            .I0(n3206), .I1(VCC_net), .CO(n52363));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_30_lut (.I0(GND_net), 
            .I1(n3207), .I2(VCC_net), .I3(n52361), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_115[5]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i30221_2_lut (.I0(duty[5]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5451));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30221_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1238_3_lut (.I0(n1819), 
            .I1(n1886), .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_6 (.CI(n51916), 
            .I0(n1730), .I1(GND_net), .CO(n51917));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1305_3_lut (.I0(n1918), 
            .I1(n1985), .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1372_3_lut (.I0(n2017), 
            .I1(n2084), .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1787_3_lut (.I0(n2624), 
            .I1(n2691), .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1439_3_lut (.I0(n2116), 
            .I1(n2183), .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_7 (.CI(n51691), 
            .I0(n929), .I1(GND_net), .CO(n51692));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1506_3_lut (.I0(n2215), 
            .I1(n2282), .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_5_lut (.I0(GND_net), 
            .I1(n1731), .I2(VCC_net), .I3(n51915), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11999_bdd_4_lut_54819 (.I0(n11999), .I1(n419), .I2(current[15]), 
            .I3(duty[23]), .O(n71047));
    defparam n11999_bdd_4_lut_54819.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_5_lut (.I0(GND_net), 
            .I1(n3031), .I2(VCC_net), .I3(n52279), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1573_3_lut (.I0(n2314), 
            .I1(n2381), .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_5 (.CI(n51915), 
            .I0(n1731), .I1(VCC_net), .CO(n51916));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1640_3_lut (.I0(n2413), 
            .I1(n2480), .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1854_3_lut (.I0(n2723), 
            .I1(n2790), .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_5 (.CI(n52201), 
            .I0(n2731), .I1(VCC_net), .CO(n52202));
    SB_LUT4 n71047_bdd_4_lut (.I0(n71047), .I1(duty[22]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam n71047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_6_lut (.I0(GND_net), 
            .I1(n930), .I2(GND_net), .I3(n51690), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_5 (.CI(n52279), 
            .I0(n3031), .I1(VCC_net), .CO(n52280));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1311_3_lut (.I0(n1924), 
            .I1(n1991), .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1707_3_lut (.I0(n2512), 
            .I1(n2579), .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54809 (.I0(n11999), .I1(n420), .I2(current[15]), 
            .I3(duty[23]), .O(n71041));
    defparam n11999_bdd_4_lut_54809.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_6 (.CI(n51690), 
            .I0(n930), .I1(GND_net), .CO(n51691));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_4_lut (.I0(GND_net), 
            .I1(n2732), .I2(GND_net), .I3(n52200), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_2_lut (.I0(GND_net), 
            .I1(n947), .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_5_lut (.I0(GND_net), 
            .I1(n931), .I2(VCC_net), .I3(n51689), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_2 (.CI(VCC_net), 
            .I0(n947), .I1(GND_net), .CO(n52089));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1378_3_lut (.I0(n2023), 
            .I1(n2090), .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_4 (.CI(n52200), 
            .I0(n2732), .I1(GND_net), .CO(n52201));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1774_3_lut (.I0(n2611), 
            .I1(n2678), .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30220_2_lut (.I0(duty[6]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5450));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30220_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_4_lut (.I0(GND_net), 
            .I1(n1732), .I2(GND_net), .I3(n51914), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_21_lut (.I0(GND_net), 
            .I1(n2115), .I2(VCC_net), .I3(n52088), .O(n2182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_4 (.CI(n51914), 
            .I0(n1732), .I1(GND_net), .CO(n51915));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_3_lut (.I0(GND_net), 
            .I1(n1733), .I2(VCC_net), .I3(n51913), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1841_3_lut (.I0(n2710), 
            .I1(n2777), .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_30 (.CI(n52361), 
            .I0(n3207), .I1(VCC_net), .CO(n52362));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_20_lut (.I0(GND_net), 
            .I1(n2116), .I2(VCC_net), .I3(n52087), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_5 (.CI(n51689), 
            .I0(n931), .I1(VCC_net), .CO(n51690));
    SB_LUT4 i43760_3_lut (.I0(n4_adj_5960), .I1(n7905), .I2(n59878), .I3(GND_net), 
            .O(n59881));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43760_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_20 (.CI(n52087), 
            .I0(n2116), .I1(VCC_net), .CO(n52088));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_3 (.CI(n51913), 
            .I0(n1733), .I1(VCC_net), .CO(n51914));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_19_lut (.I0(GND_net), 
            .I1(n2117), .I2(VCC_net), .I3(n52086), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_2_lut (.I0(GND_net), 
            .I1(n942), .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_4_lut (.I0(GND_net), 
            .I1(n3032), .I2(GND_net), .I3(n52278), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51631_2_lut (.I0(n43), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n67082));   // verilog/neopixel.v(34[12] 116[6])
    defparam i51631_2_lut.LUT_INIT = 16'h2222;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 i43761_3_lut (.I0(encoder0_position_scaled_23__N_319[29]), .I1(n59881), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43761_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_2 (.CI(VCC_net), 
            .I0(n942), .I1(GND_net), .CO(n51913));
    SB_LUT4 i20_4_lut (.I0(n67082), .I1(n67080), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n57856));   // verilog/neopixel.v(34[12] 116[6])
    defparam i20_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_29_lut (.I0(GND_net), 
            .I1(n3208), .I2(VCC_net), .I3(n52360), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_19 (.CI(n52086), 
            .I0(n2117), .I1(VCC_net), .CO(n52087));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_4_lut (.I0(GND_net), 
            .I1(n932), .I2(GND_net), .I3(n51688), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_4 (.CI(n51688), 
            .I0(n932), .I1(GND_net), .CO(n51689));
    SB_LUT4 i54289_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70464));
    defparam i54289_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_3_lut (.I0(GND_net), 
            .I1(n933), .I2(VCC_net), .I3(n51687), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_3_lut (.I0(GND_net), 
            .I1(n2733), .I2(VCC_net), .I3(n52199), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_18_lut (.I0(GND_net), 
            .I1(n2118), .I2(VCC_net), .I3(n52085), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_18 (.CI(n52085), 
            .I0(n2118), .I1(VCC_net), .CO(n52086));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_4 (.CI(n52278), 
            .I0(n3032), .I1(GND_net), .CO(n52279));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_3 (.CI(n51687), 
            .I0(n933), .I1(VCC_net), .CO(n51688));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_29 (.CI(n52360), 
            .I0(n3208), .I1(VCC_net), .CO(n52361));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_17_lut (.I0(GND_net), 
            .I1(n2119), .I2(VCC_net), .I3(n52084), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_28_lut (.I0(GND_net), 
            .I1(n3209), .I2(VCC_net), .I3(n52359), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_28 (.CI(n52359), 
            .I0(n3209), .I1(VCC_net), .CO(n52360));
    SB_CARRY add_174_30 (.CI(n51385), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n51386));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1096_1_lut (.I0(n296), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n5246));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1096_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_174_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n51384), .O(n1535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71041_bdd_4_lut (.I0(n71041), .I1(duty[21]), .I2(n249), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam n71041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30219_2_lut (.I0(duty[7]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5449));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30219_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_174_29 (.CI(n51384), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n51385));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1445_3_lut (.I0(n2122), 
            .I1(n2189), .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54804 (.I0(n11999), .I1(n421), .I2(current[15]), 
            .I3(duty[23]), .O(n71035));
    defparam n11999_bdd_4_lut_54804.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_27_lut (.I0(GND_net), 
            .I1(n3210), .I2(VCC_net), .I3(n52358), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_2_lut (.I0(GND_net), 
            .I1(n934), .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_27 (.CI(n52358), 
            .I0(n3210), .I1(VCC_net), .CO(n52359));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71035_bdd_4_lut (.I0(n71035), .I1(duty[20]), .I2(n250), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam n71035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5880));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_3_lut (.I0(GND_net), 
            .I1(n3033), .I2(VCC_net), .I3(n52277), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_3 (.CI(n52199), 
            .I0(n2733), .I1(VCC_net), .CO(n52200));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_17 (.CI(n52084), 
            .I0(n2119), .I1(VCC_net), .CO(n52085));
    SB_LUT4 add_264_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n51324), .O(encoder1_position_scaled_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30218_2_lut (.I0(duty[8]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5448));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30218_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_2 (.CI(VCC_net), 
            .I0(n934), .I1(GND_net), .CO(n51687));
    SB_CARRY add_262_17 (.CI(n51351), .I0(duty[18]), .I1(n70691), .CO(n51352));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_8_lut (.I0(n861), 
            .I1(n828), .I2(VCC_net), .I3(n51686), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5881));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15800_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n23164), .I3(GND_net), .O(n30207));   // verilog/coms.v(130[12] 305[6])
    defparam i15800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30217_2_lut (.I0(duty[9]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5447));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30217_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1512_3_lut (.I0(n2221), 
            .I1(n2288), .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54799 (.I0(n11999), .I1(n422), .I2(current[15]), 
            .I3(duty[23]), .O(n71029));
    defparam n11999_bdd_4_lut_54799.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_16_lut (.I0(GND_net), 
            .I1(n2120), .I2(VCC_net), .I3(n52083), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_16 (.CI(n52083), 
            .I0(n2120), .I1(VCC_net), .CO(n52084));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_3 (.CI(n52277), 
            .I0(n3033), .I1(VCC_net), .CO(n52278));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_2_lut (.I0(GND_net), 
            .I1(n952), .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_15_lut (.I0(GND_net), 
            .I1(n2121), .I2(VCC_net), .I3(n52082), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_2 (.CI(VCC_net), 
            .I0(n952), .I1(GND_net), .CO(n52199));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_15 (.CI(n52082), 
            .I0(n2121), .I1(VCC_net), .CO(n52083));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_14_lut (.I0(GND_net), 
            .I1(n2122), .I2(VCC_net), .I3(n52081), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_14 (.CI(n52081), 
            .I0(n2122), .I1(VCC_net), .CO(n52082));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_2_lut (.I0(GND_net), 
            .I1(n955), .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_26_lut (.I0(GND_net), 
            .I1(n3211), .I2(VCC_net), .I3(n52357), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_7_lut (.I0(GND_net), 
            .I1(n829), .I2(GND_net), .I3(n51685), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_26 (.CI(n52357), 
            .I0(n3211), .I1(VCC_net), .CO(n52358));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_25_lut (.I0(GND_net), 
            .I1(n3212), .I2(VCC_net), .I3(n52356), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_115[6]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_282_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_115[7]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i30216_2_lut (.I0(duty[10]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5446));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30216_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_13_lut (.I0(GND_net), 
            .I1(n2123), .I2(VCC_net), .I3(n52080), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_7 (.CI(n51685), 
            .I0(n829), .I1(GND_net), .CO(n51686));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_26_lut (.I0(GND_net), 
            .I1(n2610), .I2(VCC_net), .I3(n52198), .O(n2677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n51316), .O(encoder1_position_scaled_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_13 (.CI(n52080), 
            .I0(n2123), .I1(VCC_net), .CO(n52081));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_25_lut (.I0(GND_net), 
            .I1(n2611), .I2(VCC_net), .I3(n52197), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_16_lut (.I0(current[15]), .I1(duty[17]), .I2(n70691), 
            .I3(n51350), .O(n256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_16_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_6_lut (.I0(GND_net), 
            .I1(n830), .I2(GND_net), .I3(n51684), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_25 (.CI(n52356), 
            .I0(n3212), .I1(VCC_net), .CO(n52357));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_24_lut (.I0(GND_net), 
            .I1(n3213), .I2(VCC_net), .I3(n52355), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_6 (.CI(n51684), 
            .I0(n830), .I1(GND_net), .CO(n51685));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_24 (.CI(n52355), 
            .I0(n3213), .I1(VCC_net), .CO(n52356));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_23_lut (.I0(GND_net), 
            .I1(n3214), .I2(VCC_net), .I3(n52354), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_12_lut (.I0(GND_net), 
            .I1(n2124), .I2(VCC_net), .I3(n52079), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_25 (.CI(n52197), 
            .I0(n2611), .I1(VCC_net), .CO(n52198));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_23 (.CI(n52354), 
            .I0(n3214), .I1(VCC_net), .CO(n52355));
    SB_CARRY add_264_13 (.CI(n51324), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n51325));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_5_lut (.I0(GND_net), 
            .I1(n831), .I2(VCC_net), .I3(n51683), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_5 (.CI(n51683), 
            .I0(n831), .I1(VCC_net), .CO(n51684));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_22_lut (.I0(GND_net), 
            .I1(n3215), .I2(VCC_net), .I3(n52353), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_4_lut (.I0(GND_net), 
            .I1(n832), .I2(GND_net), .I3(n51682), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_12 (.CI(n52079), 
            .I0(n2124), .I1(VCC_net), .CO(n52080));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_22 (.CI(n52353), 
            .I0(n3215), .I1(VCC_net), .CO(n52354));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_2 (.CI(VCC_net), 
            .I0(n955), .I1(GND_net), .CO(n52277));
    SB_LUT4 i15801_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n59079), 
            .I3(GND_net), .O(n30208));   // verilog/coms.v(130[12] 305[6])
    defparam i15801_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_4 (.CI(n51682), 
            .I0(n832), .I1(GND_net), .CO(n51683));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_24_lut (.I0(GND_net), 
            .I1(n2612), .I2(VCC_net), .I3(n52196), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i837_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_24 (.CI(n52196), 
            .I0(n2612), .I1(VCC_net), .CO(n52197));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_11_lut (.I0(GND_net), 
            .I1(n2125), .I2(VCC_net), .I3(n52078), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n51383), .O(n1536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_29_lut (.I0(n70178), 
            .I1(n2907), .I2(VCC_net), .I3(n52276), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_21_lut (.I0(GND_net), 
            .I1(n3216), .I2(VCC_net), .I3(n52352), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_115[8]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i9_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_11 (.CI(n52078), 
            .I0(n2125), .I1(VCC_net), .CO(n52079));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2132_3_lut (.I0(n3129), 
            .I1(n3196), .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_3_lut (.I0(GND_net), 
            .I1(n833), .I2(VCC_net), .I3(n51681), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_28 (.CI(n51383), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n51384));
    SB_LUT4 add_174_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n51382), .O(n1537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_10_lut (.I0(GND_net), 
            .I1(n2126), .I2(VCC_net), .I3(n52077), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_21 (.CI(n52352), 
            .I0(n3216), .I1(VCC_net), .CO(n52353));
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n1921), .I1(n60745), .I2(n1923), .I3(n1924), 
            .O(n63334));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_CARRY add_174_27 (.CI(n51382), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n51383));
    SB_LUT4 add_174_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n51381), .O(n1538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_262_16 (.CI(n51350), .I0(duty[17]), .I1(n70691), .CO(n51351));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i904_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_3 (.CI(n51681), 
            .I0(n833), .I1(VCC_net), .CO(n51682));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_565_2_lut (.I0(GND_net), 
            .I1(n519), .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_10 (.CI(n52077), 
            .I0(n2126), .I1(VCC_net), .CO(n52078));
    SB_LUT4 add_262_15_lut (.I0(current[15]), .I1(duty[16]), .I2(n70691), 
            .I3(n51349), .O(n257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_15_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_20_lut (.I0(GND_net), 
            .I1(n3217), .I2(VCC_net), .I3(n52351), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_565_2 (.CI(VCC_net), 
            .I0(n519), .I1(GND_net), .CO(n51681));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1579_3_lut (.I0(n2320), 
            .I1(n2387), .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n1918), .I1(n1920), .I2(n1922), .I3(n63022), 
            .O(n63028));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_CARRY add_174_26 (.CI(n51381), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n51382));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_28_lut (.I0(GND_net), 
            .I1(n2908), .I2(VCC_net), .I3(n52275), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_28 (.CI(n52275), 
            .I0(n2908), .I1(VCC_net), .CO(n52276));
    SB_LUT4 add_174_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n51380), .O(n1539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_23_lut (.I0(GND_net), 
            .I1(n2613), .I2(VCC_net), .I3(n52195), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_25 (.CI(n51380), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n51381));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_9_lut (.I0(GND_net), 
            .I1(n2127), .I2(VCC_net), .I3(n52076), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_9 (.CI(n52076), 
            .I0(n2127), .I1(VCC_net), .CO(n52077));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_20 (.CI(n52351), 
            .I0(n3217), .I1(VCC_net), .CO(n52352));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_8_lut (.I0(GND_net), 
            .I1(n2128), .I2(VCC_net), .I3(n52075), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_23 (.CI(n52195), 
            .I0(n2613), .I1(VCC_net), .CO(n52196));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_22_lut (.I0(GND_net), 
            .I1(n2614), .I2(VCC_net), .I3(n52194), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2528_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n51680), 
            .O(n7903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2528_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n51679), 
            .O(n7904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n51379), .O(n1540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_24 (.CI(n51379), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n51380));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_22 (.CI(n52194), 
            .I0(n2614), .I1(VCC_net), .CO(n52195));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_19_lut (.I0(GND_net), 
            .I1(n3218), .I2(VCC_net), .I3(n52350), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_8 (.CI(n52075), 
            .I0(n2128), .I1(VCC_net), .CO(n52076));
    SB_LUT4 add_174_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n51378), .O(n1541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71029_bdd_4_lut (.I0(n71029), .I1(duty[19]), .I2(n251), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[19]));
    defparam n71029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_7_lut (.I0(GND_net), 
            .I1(n2129), .I2(GND_net), .I3(n52074), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2528_6 (.CI(n51679), .I0(n622), .I1(GND_net), .CO(n51680));
    SB_LUT4 add_2528_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n51678), 
            .O(n7905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_7 (.CI(n52074), 
            .I0(n2129), .I1(GND_net), .CO(n52075));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1038_3_lut (.I0(n1523), 
            .I1(n1590), .I2(n1554_adj_5994), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_6_lut (.I0(GND_net), 
            .I1(n2130), .I2(GND_net), .I3(n52073), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2528_5 (.CI(n51678), .I0(n623), .I1(VCC_net), .CO(n51679));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_19 (.CI(n52350), 
            .I0(n3218), .I1(VCC_net), .CO(n52351));
    SB_CARRY add_174_23 (.CI(n51378), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n51379));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_21_lut (.I0(GND_net), 
            .I1(n2615), .I2(VCC_net), .I3(n52193), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_6 (.CI(n52073), 
            .I0(n2130), .I1(GND_net), .CO(n52074));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1646_3_lut (.I0(n2419), 
            .I1(n2486), .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_5_lut (.I0(GND_net), 
            .I1(n2131), .I2(VCC_net), .I3(n52072), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n51377), .O(n1542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_21 (.CI(n52193), 
            .I0(n2615), .I1(VCC_net), .CO(n52194));
    SB_CARRY add_262_15 (.CI(n51349), .I0(duty[16]), .I1(n70691), .CO(n51350));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_5 (.CI(n52072), 
            .I0(n2131), .I1(VCC_net), .CO(n52073));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1713_3_lut (.I0(n2518), 
            .I1(n2585), .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_4_lut (.I0(GND_net), 
            .I1(n2132), .I2(GND_net), .I3(n52071), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2528_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n51677), 
            .O(n7906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2528_4 (.CI(n51677), .I0(n516), .I1(GND_net), .CO(n51678));
    SB_CARRY add_174_22 (.CI(n51377), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n51378));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_16_lut (.I0(n70527), 
            .I1(n1620), .I2(VCC_net), .I3(n51894), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2528_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n51676), 
            .O(n7907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n51376), .O(n1543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30215_2_lut (.I0(duty[11]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5445));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30215_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY add_2528_3 (.CI(n51676), .I0(n625), .I1(VCC_net), .CO(n51677));
    SB_LUT4 add_2528_2_lut (.I0(GND_net), .I1(n518), .I2(GND_net), .I3(VCC_net), 
            .O(n7908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2528_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_4 (.CI(n52071), 
            .I0(n2132), .I1(GND_net), .CO(n52072));
    SB_CARRY add_2528_2 (.CI(VCC_net), .I0(n518), .I1(GND_net), .CO(n51676));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1105_3_lut (.I0(n1622), 
            .I1(n1689), .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1172_3_lut (.I0(n1721), 
            .I1(n1788), .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_15_lut (.I0(GND_net), 
            .I1(n1621), .I2(VCC_net), .I3(n51893), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_14_lut (.I0(current[15]), .I1(duty[15]), .I2(n70691), 
            .I3(n51348), .O(n258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_14_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_15 (.CI(n51893), 
            .I0(n1621), .I1(VCC_net), .CO(n51894));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_18_lut (.I0(GND_net), 
            .I1(n3219), .I2(VCC_net), .I3(n52349), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_20_lut (.I0(GND_net), 
            .I1(n2616), .I2(VCC_net), .I3(n52192), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_20 (.CI(n52192), 
            .I0(n2616), .I1(VCC_net), .CO(n52193));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_27_lut (.I0(GND_net), 
            .I1(n2909), .I2(VCC_net), .I3(n52274), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_3_lut (.I0(GND_net), 
            .I1(n2133), .I2(VCC_net), .I3(n52070), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_19_lut (.I0(GND_net), 
            .I1(n2617), .I2(VCC_net), .I3(n52191), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_14_lut (.I0(GND_net), 
            .I1(n1622), .I2(VCC_net), .I3(n51892), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_27 (.CI(n52274), 
            .I0(n2909), .I1(VCC_net), .CO(n52275));
    SB_LUT4 i54146_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70321));
    defparam i54146_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_14 (.CI(n51892), 
            .I0(n1622), .I1(VCC_net), .CO(n51893));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_13_lut (.I0(GND_net), 
            .I1(n1623), .I2(VCC_net), .I3(n51891), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_13 (.CI(n51891), 
            .I0(n1623), .I1(VCC_net), .CO(n51892));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_3 (.CI(n52070), 
            .I0(n2133), .I1(VCC_net), .CO(n52071));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_12_lut (.I0(GND_net), 
            .I1(n1624), .I2(VCC_net), .I3(n51890), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_12 (.CI(n51890), 
            .I0(n1624), .I1(VCC_net), .CO(n51891));
    SB_CARRY add_174_21 (.CI(n51376), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n51377));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_11_lut (.I0(GND_net), 
            .I1(n1625), .I2(VCC_net), .I3(n51889), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_11 (.CI(n51889), 
            .I0(n1625), .I1(VCC_net), .CO(n51890));
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [7]), .I1(n44625), .I2(n28768), 
            .I3(rx_data[7]), .O(n58340));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_174_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n51375), .O(n1544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_20_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_10_lut (.I0(GND_net), 
            .I1(n1626), .I2(VCC_net), .I3(n51888), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1436_2_lut (.I0(GND_net), 
            .I1(n946), .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_19 (.CI(n52191), 
            .I0(n2617), .I1(VCC_net), .CO(n52192));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_10 (.CI(n51888), 
            .I0(n1626), .I1(VCC_net), .CO(n51889));
    SB_CARRY add_174_20 (.CI(n51375), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n51376));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1436_2 (.CI(VCC_net), 
            .I0(n946), .I1(GND_net), .CO(n52070));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_9_lut (.I0(GND_net), 
            .I1(n1627), .I2(VCC_net), .I3(n51887), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_9 (.CI(n51887), 
            .I0(n1627), .I1(VCC_net), .CO(n51888));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_18_lut (.I0(GND_net), 
            .I1(n2618), .I2(VCC_net), .I3(n52190), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_8_lut (.I0(GND_net), 
            .I1(n1628), .I2(VCC_net), .I3(n51886), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_8 (.CI(n51886), 
            .I0(n1628), .I1(VCC_net), .CO(n51887));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_7_lut (.I0(GND_net), 
            .I1(n1629), .I2(GND_net), .I3(n51885), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1239_3_lut (.I0(n1820), 
            .I1(n1887), .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_18 (.CI(n52349), 
            .I0(n3219), .I1(VCC_net), .CO(n52350));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_6050));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53955_1_lut (.I0(n44815), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70130));
    defparam i53955_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2194_3_lut (.I0(n3223), 
            .I1(n3290), .I2(n3237), .I3(GND_net), .O(n25_adj_6059));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2193_3_lut (.I0(n3222), 
            .I1(n3289), .I2(n3237), .I3(GND_net), .O(n27_adj_6060));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2200_3_lut (.I0(n3229), 
            .I1(n3296), .I2(n3237), .I3(GND_net), .O(n13_adj_6056));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2198_3_lut (.I0(n3227), 
            .I1(n3294), .I2(n3237), .I3(GND_net), .O(n17_adj_6057));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2195_3_lut (.I0(n3224), 
            .I1(n3291), .I2(n3237), .I3(GND_net), .O(n23_adj_6058));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n3220), .I1(n25_adj_6059), .I2(n3287), 
            .I3(n3237), .O(n63132));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n3226), .I1(n13_adj_6056), .I2(n3293), 
            .I3(n3237), .O(n63134));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n3221), .I1(n17_adj_6057), .I2(n3288), 
            .I3(n3237), .O(n63136));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n3225), .I1(n23_adj_6058), .I2(n3292), 
            .I3(n3237), .O(n63140));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2190_3_lut (.I0(n3219), 
            .I1(n3286), .I2(n3237), .I3(GND_net), .O(n33_adj_6061));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n3228), .I1(n27_adj_6060), .I2(n3295), 
            .I3(n3237), .O(n63138));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_17_lut (.I0(GND_net), 
            .I1(n3220), .I2(VCC_net), .I3(n52348), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n3218), .I1(n33_adj_6061), .I2(n3285), 
            .I3(n3237), .O(n63142));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2188_3_lut (.I0(n3217), 
            .I1(n3284), .I2(n3237), .I3(GND_net), .O(n37_adj_6062));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n63140), .I1(n63136), .I2(n63134), 
            .I3(n63132), .O(n63150));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n63150), .I1(n37_adj_6062), .I2(n63142), 
            .I3(n63138), .O(n63154));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i30417_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n44717));
    defparam i30417_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i30419_4_lut (.I0(n44717), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n44719));
    defparam i30419_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n67030), .I2(n3237), .I3(n3230), 
            .O(n5_adj_6051));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n3216), .I1(n63154), .I2(n3283), .I3(n3237), 
            .O(n63156));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'heefc;
    SB_LUT4 i30503_4_lut (.I0(n44719), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n44807));
    defparam i30503_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2186_3_lut (.I0(n3215), 
            .I1(n3282), .I2(n3237), .I3(GND_net), .O(n41_adj_6063));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n41_adj_6063), .I1(n44807), .I2(n63156), 
            .I3(n5_adj_6051), .O(n63160));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n3214), .I1(n63160), .I2(n3281), .I3(n3237), 
            .O(n63162));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n3213), .I1(n63162), .I2(n3280), .I3(n3237), 
            .O(n63164));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n3212), .I1(n63164), .I2(n3279), .I3(n3237), 
            .O(n63166));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'heefc;
    SB_LUT4 i15596_3_lut (.I0(\data_in_frame[0] [7]), .I1(rx_data[7]), .I2(n60009), 
            .I3(GND_net), .O(n30003));   // verilog/coms.v(130[12] 305[6])
    defparam i15596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n3211), .I1(n63166), .I2(n3278), .I3(n3237), 
            .O(n63168));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n3210), .I1(n63168), .I2(n3277), .I3(n3237), 
            .O(n63170));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'heefc;
    SB_LUT4 i51382_4_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n60), .I2(\FRAME_MATCHER.i [3]), 
            .I3(n59967), .O(n67059));   // verilog/coms.v(94[13:20])
    defparam i51382_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 n11999_bdd_4_lut_54794 (.I0(n11999), .I1(n423), .I2(current[15]), 
            .I3(duty[23]), .O(n71023));
    defparam n11999_bdd_4_lut_54794.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1306_3_lut (.I0(n1919), 
            .I1(n1986), .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n3209), .I1(n63170), .I2(n3276), .I3(n3237), 
            .O(n63172));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n3208), .I1(n63172), .I2(n3275), .I3(n3237), 
            .O(n63174));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n3207), .I1(n63174), .I2(n3274), .I3(n3237), 
            .O(n63176));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1373_3_lut (.I0(n2018), 
            .I1(n2085), .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n3206), .I1(n63176), .I2(n3273), .I3(n3237), 
            .O(n63178));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n3205), .I1(n63178), .I2(n3272), .I3(n3237), 
            .O(n63180));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'heefc;
    SB_LUT4 i53958_4_lut (.I0(n63180), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n44815));
    defparam i53958_4_lut.LUT_INIT = 16'h1105;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position_scaled_23__N_319[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_6049));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54310_4_lut (.I0(n63028), .I1(n1917), .I2(n63334), .I3(n1919), 
            .O(n1950));
    defparam i54310_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i27854_4_lut (.I0(n67059), .I1(n51), .I2(rx_data[2]), .I3(\data_in_frame[23] [2]), 
            .O(n42182));   // verilog/coms.v(94[13:20])
    defparam i27854_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27855_3_lut (.I0(n42182), .I1(\data_in_frame[23] [2]), .I2(reset), 
            .I3(GND_net), .O(n30465));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position_scaled_23__N_319[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_6048));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position_scaled_23__N_319[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_6047));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position_scaled_23__N_319[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_6046));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position_scaled_23__N_319[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_6045));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53950_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70125));
    defparam i53950_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut (.I0(n3220), .I1(n3218), .I2(n3225), .I3(GND_net), 
            .O(n63714));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n3224), .I1(n3228), .I2(n3227), .I3(n3223), 
            .O(n63644));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1440_3_lut (.I0(n2117), 
            .I1(n2184), .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1773 (.I0(n3222), .I1(n3217), .I2(n3226), .I3(GND_net), 
            .O(n63642));
    defparam i1_3_lut_adj_1773.LUT_INIT = 16'hfefe;
    SB_LUT4 i15588_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n60009), 
            .I3(GND_net), .O(n29995));   // verilog/coms.v(130[12] 305[6])
    defparam i15588_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_17 (.CI(n52348), 
            .I0(n3220), .I1(VCC_net), .CO(n52349));
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n3214), .I1(n3215), .I2(n63642), .I3(n63644), 
            .O(n63650));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n3210), .I1(n3211), .I2(n3213), .I3(n63650), 
            .O(n63656));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i30501_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n44805));
    defparam i30501_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n3216), .I1(n63714), .I2(n3221), .I3(n3219), 
            .O(n63718));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1507_3_lut (.I0(n2216), 
            .I1(n2283), .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15585_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n60009), 
            .I3(GND_net), .O(n29992));   // verilog/coms.v(130[12] 305[6])
    defparam i15585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n3229), .I1(n44805), .I2(n3230), .I3(n3231), 
            .O(n60850));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n63656), 
            .O(n63662));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i15582_3_lut (.I0(\data_in_frame[0] [4]), .I1(rx_data[4]), .I2(n60009), 
            .I3(GND_net), .O(n29989));   // verilog/coms.v(130[12] 305[6])
    defparam i15582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n3205), .I1(n3212), .I2(n60850), .I3(n63718), 
            .O(n63724));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 i53954_4_lut (.I0(n3206), .I1(n63724), .I2(n63662), .I3(n3204), 
            .O(n3237));
    defparam i53954_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position_scaled_23__N_319[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_6044));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position_scaled_23__N_319[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_6043));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position_scaled_23__N_319[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_6042));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position_scaled_23__N_319[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_6041));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53914_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70089));
    defparam i53914_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position_scaled_23__N_319[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_6040));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15579_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n60009), 
            .I3(GND_net), .O(n29986));   // verilog/coms.v(130[12] 305[6])
    defparam i15579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_2_lut (.I0(n188), .I1(n136), .I2(GND_net), .I3(GND_net), 
            .O(n37));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1574_3_lut (.I0(n2315), 
            .I1(n2382), .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position_scaled_23__N_319[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_6039));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position_scaled_23__N_319[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_6038));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position_scaled_23__N_319[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_6037));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_26_lut (.I0(GND_net), 
            .I1(n2910), .I2(VCC_net), .I3(n52273), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position_scaled_23__N_319[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_6036));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position_scaled_23__N_319[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_6035));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_26 (.CI(n52273), 
            .I0(n2910), .I1(VCC_net), .CO(n52274));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1641_3_lut (.I0(n2414), 
            .I1(n2481), .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1780 (.I0(n37023), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_1780.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position_scaled_23__N_319[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_6034));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15576_3_lut (.I0(\data_in_frame[0] [2]), .I1(rx_data[2]), .I2(n60009), 
            .I3(GND_net), .O(n29983));   // verilog/coms.v(130[12] 305[6])
    defparam i15576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position_scaled_23__N_319[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_6033));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_18 (.CI(n52190), 
            .I0(n2618), .I1(VCC_net), .CO(n52191));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position_scaled_23__N_319[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_6032));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53880_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70055));
    defparam i53880_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position_scaled_23__N_319[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_6031));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position_scaled_23__N_319[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_6030));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position_scaled_23__N_319[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_6029));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_7 (.CI(n51885), 
            .I0(n1629), .I1(GND_net), .CO(n51886));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1708_3_lut (.I0(n2513), 
            .I1(n2580), .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position_scaled_23__N_319[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_6028));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position_scaled_23__N_319[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_6027));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position_scaled_23__N_319[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_6026));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position_scaled_23__N_319[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_6025));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position_scaled_23__N_319[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_6024));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position_scaled_23__N_319[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_6023));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_6_lut (.I0(GND_net), 
            .I1(n1630), .I2(GND_net), .I3(n51884), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position_scaled_23__N_319[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_6022));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_17_lut (.I0(GND_net), 
            .I1(n2619), .I2(VCC_net), .I3(n52189), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position_scaled_23__N_319[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_6021));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position_scaled_23__N_319[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_6020));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54003_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70178));
    defparam i54003_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1775_3_lut (.I0(n2612), 
            .I1(n2679), .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54115_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70290));
    defparam i54115_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30214_2_lut (.I0(duty[12]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5444));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30214_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_6 (.CI(n51884), 
            .I0(n1630), .I1(GND_net), .CO(n51885));
    SB_LUT4 i1_2_lut_adj_1781 (.I0(\PID_CONTROLLER.integral_23__N_3844 [12]), 
            .I1(Ki[1]), .I2(GND_net), .I3(GND_net), .O(n110));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1248_3_lut (.I0(n1829), 
            .I1(n1896), .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21219_3_lut (.I0(n60009), .I1(rx_data[1]), .I2(\data_in_frame[0] [1]), 
            .I3(GND_net), .O(n30539));   // verilog/coms.v(94[13:20])
    defparam i21219_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_17 (.CI(n52189), 
            .I0(n2619), .I1(VCC_net), .CO(n52190));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1842_3_lut (.I0(n2711), 
            .I1(n2778), .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_5_lut (.I0(GND_net), 
            .I1(n1631), .I2(VCC_net), .I3(n51883), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_5 (.CI(n51883), 
            .I0(n1631), .I1(VCC_net), .CO(n51884));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1909_3_lut (.I0(n2810), 
            .I1(n2877), .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_25_lut (.I0(GND_net), 
            .I1(n2911), .I2(VCC_net), .I3(n52272), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[22] [7]), .I1(n28723), .I2(n28770), 
            .I3(rx_data[7]), .O(n58198));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_4_lut (.I0(GND_net), 
            .I1(n1632), .I2(GND_net), .I3(n51882), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_16_lut (.I0(GND_net), 
            .I1(n3221), .I2(VCC_net), .I3(n52347), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_4 (.CI(n51882), 
            .I0(n1632), .I1(GND_net), .CO(n51883));
    SB_LUT4 i15561_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n28770), .I3(GND_net), .O(n29968));   // verilog/coms.v(130[12] 305[6])
    defparam i15561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15557_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n28770), .I3(GND_net), .O(n29964));   // verilog/coms.v(130[12] 305[6])
    defparam i15557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15554_3_lut (.I0(\data_in_frame[22] [4]), .I1(rx_data[4]), 
            .I2(n28770), .I3(GND_net), .O(n29961));   // verilog/coms.v(130[12] 305[6])
    defparam i15554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_174_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n51374), .O(n1545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15551_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n28770), .I3(GND_net), .O(n29958));   // verilog/coms.v(130[12] 305[6])
    defparam i15551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1907_3_lut (.I0(n2808), 
            .I1(n2875), .I2(n2841), .I3(GND_net), .O(n2907));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1782 (.I0(\data_in_frame[22] [2]), .I1(n28723), 
            .I2(n28770), .I3(rx_data[2]), .O(n58202));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1782.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_3_lut (.I0(GND_net), 
            .I1(n1633), .I2(VCC_net), .I3(n51881), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1908_3_lut (.I0(n2809), 
            .I1(n2876), .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15545_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n28770), .I3(GND_net), .O(n29952));   // verilog/coms.v(130[12] 305[6])
    defparam i15545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(duty[2]), .I1(duty[23]), .I2(duty[1]), .I3(duty[0]), 
            .O(n211));   // verilog/TinyFPGA_B.v(111[25:31])
    defparam i14_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_16_lut (.I0(GND_net), 
            .I1(n2620), .I2(VCC_net), .I3(n52188), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15542_3_lut (.I0(\data_in_frame[22] [0]), .I1(rx_data[0]), 
            .I2(n28770), .I3(GND_net), .O(n29949));   // verilog/coms.v(130[12] 305[6])
    defparam i15542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1783 (.I0(\data_in_frame[21] [7]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[7]), .O(n58208));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1783.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i15_3_lut (.I0(encoder0_position_scaled_23__N_319[14]), 
            .I1(n19_adj_5945), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30213_2_lut (.I0(duty[13]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5443));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30213_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_3 (.CI(n51881), 
            .I0(n1633), .I1(VCC_net), .CO(n51882));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_16 (.CI(n52188), 
            .I0(n2620), .I1(VCC_net), .CO(n52189));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_25 (.CI(n52272), 
            .I0(n2911), .I1(VCC_net), .CO(n52273));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_24_lut (.I0(GND_net), 
            .I1(n2912), .I2(VCC_net), .I3(n52271), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1784 (.I0(\data_in_frame[21] [6]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[6]), .O(n58212));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1784.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_16 (.CI(n52347), 
            .I0(n3221), .I1(VCC_net), .CO(n52348));
    SB_LUT4 i54084_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70259));
    defparam i54084_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_1785 (.I0(\data_in_frame[21] [5]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[5]), .O(n58216));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1785.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_15_lut (.I0(GND_net), 
            .I1(n3222), .I2(VCC_net), .I3(n52346), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71023_bdd_4_lut (.I0(n71023), .I1(duty[18]), .I2(n252), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[18]));
    defparam n71023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1786 (.I0(\data_in_frame[21] [4]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[4]), .O(n58220));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1786.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1780_3_lut (.I0(n2617), 
            .I1(n2684), .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54789 (.I0(n11999), .I1(n424), .I2(current[15]), 
            .I3(duty[23]), .O(n71017));
    defparam n11999_bdd_4_lut_54789.LUT_INIT = 16'he4aa;
    SB_LUT4 i37005_3_lut_4_lut (.I0(n37023), .I1(Ki[3]), .I2(n4_adj_6053), 
            .I3(n20625), .O(n6_adj_6052));
    defparam i37005_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i12_4_lut_adj_1787 (.I0(\data_in_frame[21] [3]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[3]), .O(n58224));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1787.LUT_INIT = 16'h3a0a;
    SB_LUT4 i54314_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70489));
    defparam i54314_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54226_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70401));
    defparam i54226_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1847_3_lut (.I0(n2716), 
            .I1(n2783), .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1788 (.I0(n2028), .I1(n2026), .I2(n2025), .I3(GND_net), 
            .O(n63476));
    defparam i1_3_lut_adj_1788.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1789 (.I0(\data_in_frame[21] [2]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[2]), .O(n58226));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1789.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54197_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70372));
    defparam i54197_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_174_19 (.CI(n51374), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n51375));
    SB_LUT4 n71017_bdd_4_lut (.I0(n71017), .I1(duty[17]), .I2(n253), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[17]));
    defparam n71017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1790 (.I0(\data_in_frame[21] [1]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[1]), .O(n58228));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1790.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_3_lut_4_lut (.I0(n37023), .I1(Ki[3]), .I2(n4_adj_6053), 
            .I3(n20625), .O(n20576));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i1_2_lut_adj_1791 (.I0(n42166), .I1(n8_adj_5936), .I2(GND_net), 
            .I3(GND_net), .O(n28772));
    defparam i1_2_lut_adj_1791.LUT_INIT = 16'h2222;
    SB_LUT4 mux_282_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1792 (.I0(\PID_CONTROLLER.integral_23__N_3844 [12]), 
            .I1(Ki[0]), .I2(GND_net), .I3(GND_net), .O(n38));
    defparam i1_2_lut_adj_1792.LUT_INIT = 16'h8888;
    SB_LUT4 mux_277_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_115[9]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_174_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n51373), .O(n1546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2113_3_lut (.I0(n3110), 
            .I1(n3177), .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1793 (.I0(\data_in_frame[21] [0]), .I1(n28733), 
            .I2(n28772), .I3(rx_data[0]), .O(n58230));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1793.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_15 (.CI(n52346), 
            .I0(n3222), .I1(VCC_net), .CO(n52347));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1101_2_lut (.I0(GND_net), 
            .I1(n941), .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_15_lut (.I0(GND_net), 
            .I1(n2621), .I2(VCC_net), .I3(n52187), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_18 (.CI(n51373), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n51374));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_15 (.CI(n52187), 
            .I0(n2621), .I1(VCC_net), .CO(n52188));
    SB_LUT4 i12_4_lut_adj_1794 (.I0(\data_in_frame[20] [7]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[7]), .O(n58234));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1794.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_24 (.CI(n52271), 
            .I0(n2912), .I1(VCC_net), .CO(n52272));
    SB_LUT4 i54007_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70182));
    defparam i54007_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_6073));   // verilog/TinyFPGA_B.v(389[12:17])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_6074));   // verilog/TinyFPGA_B.v(389[12:17])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1438_3_lut (.I0(n2115), 
            .I1(n2182), .I2(n2148), .I3(GND_net), .O(n2214));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54054_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70229));
    defparam i54054_1_lut.LUT_INIT = 16'h5555;
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_14_lut (.I0(GND_net), 
            .I1(n3223), .I2(VCC_net), .I3(n52345), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_23_lut (.I0(GND_net), 
            .I1(n2913), .I2(VCC_net), .I3(n52270), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1848_3_lut (.I0(n2717), 
            .I1(n2784), .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54784 (.I0(n11999), .I1(n425), .I2(current[15]), 
            .I3(duty[23]), .O(n71011));
    defparam n11999_bdd_4_lut_54784.LUT_INIT = 16'he4aa;
    SB_LUT4 n71011_bdd_4_lut (.I0(n71011), .I1(duty[16]), .I2(n254), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[16]));
    defparam n71011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1915_3_lut (.I0(n2816), 
            .I1(n2883), .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54779 (.I0(n11999), .I1(n426), .I2(current[15]), 
            .I3(duty[23]), .O(n71005));
    defparam n11999_bdd_4_lut_54779.LUT_INIT = 16'he4aa;
    SB_LUT4 n71005_bdd_4_lut (.I0(n71005), .I1(duty[15]), .I2(n255), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[15]));
    defparam n71005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1914_3_lut (.I0(n2815), 
            .I1(n2882), .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54774 (.I0(n11999), .I1(n427), .I2(current[15]), 
            .I3(duty[23]), .O(n70999));
    defparam n11999_bdd_4_lut_54774.LUT_INIT = 16'he4aa;
    SB_LUT4 n70999_bdd_4_lut (.I0(n70999), .I1(duty[14]), .I2(n256), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[14]));
    defparam n70999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1913_3_lut (.I0(n2814), 
            .I1(n2881), .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54769 (.I0(n11999), .I1(n428), .I2(current[15]), 
            .I3(duty[23]), .O(n70993));
    defparam n11999_bdd_4_lut_54769.LUT_INIT = 16'he4aa;
    SB_LUT4 n70993_bdd_4_lut (.I0(n70993), .I1(duty[13]), .I2(n257), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[13]));
    defparam n70993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i22_3_lut (.I0(encoder0_position_scaled_23__N_319[21]), 
            .I1(n12_adj_5952), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n937));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11999_bdd_4_lut_54764 (.I0(n11999), .I1(n429), .I2(current[15]), 
            .I3(duty[23]), .O(n70987));
    defparam n11999_bdd_4_lut_54764.LUT_INIT = 16'he4aa;
    SB_LUT4 n70987_bdd_4_lut (.I0(n70987), .I1(duty[12]), .I2(n258), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[12]));
    defparam n70987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531_adj_5991));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i979_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1101_2 (.CI(VCC_net), 
            .I0(n941), .I1(GND_net), .CO(n51881));
    SB_LUT4 add_174_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n51372), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29548_4_lut (.I0(n13_adj_6074), .I1(baudrate[0]), .I2(n14_adj_6073), 
            .I3(n25975), .O(n43842));
    defparam i29548_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_14_lut (.I0(GND_net), 
            .I1(n2622), .I2(VCC_net), .I3(n52186), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_17 (.CI(n51372), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n51373));
    SB_CARRY add_262_14 (.CI(n51348), .I0(duty[15]), .I1(n70691), .CO(n51349));
    SB_LUT4 add_174_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n51371), .O(n1548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_14 (.CI(n52186), 
            .I0(n2622), .I1(VCC_net), .CO(n52187));
    SB_LUT4 i12_4_lut_adj_1795 (.I0(\data_in_frame[20] [5]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[5]), .O(n58238));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1795.LUT_INIT = 16'h3a0a;
    SB_CARRY add_174_16 (.CI(n51371), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n51372));
    SB_LUT4 add_262_13_lut (.I0(current[11]), .I1(duty[14]), .I2(n70691), 
            .I3(n51347), .O(n259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_13_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_262_13 (.CI(n51347), .I0(duty[14]), .I1(n70691), .CO(n51348));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_13_lut (.I0(GND_net), 
            .I1(n2623), .I2(VCC_net), .I3(n52185), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30212_2_lut (.I0(duty[14]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5442));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30212_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1796 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_6008));
    defparam i1_2_lut_adj_1796.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_14 (.CI(n52345), 
            .I0(n3223), .I1(VCC_net), .CO(n52346));
    SB_LUT4 add_174_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n51370), .O(n1549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_15 (.CI(n51370), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n51371));
    SB_LUT4 add_174_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n51369), .O(n1550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_12_lut (.I0(current[10]), .I1(duty[13]), .I2(n70691), 
            .I3(n51346), .O(n260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_12_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1046_3_lut (.I0(n1531_adj_5991), 
            .I1(n1598), .I2(n1554_adj_5994), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_264_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n51323), .O(encoder1_position_scaled_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_13_lut (.I0(GND_net), 
            .I1(n3224), .I2(VCC_net), .I3(n52344), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5878), .I3(n51665), .O(displacement_23__N_91[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_23 (.CI(n52270), 
            .I0(n2913), .I1(VCC_net), .CO(n52271));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5877), .I3(n51664), .O(displacement_23__N_91[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_6008), .I2(delay_counter[10]), 
            .I3(n25840), .O(n61896));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_4_lut_adj_1797 (.I0(n37023), .I1(Ki[2]), .I2(n51273), 
            .I3(n20626), .O(n20577));
    defparam i1_3_lut_4_lut_adj_1797.LUT_INIT = 16'h8778;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n51664), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5877), .CO(n51665));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5876), .I3(n51663), .O(displacement_23__N_91[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_13 (.CI(n52344), 
            .I0(n3224), .I1(VCC_net), .CO(n52345));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_22_lut (.I0(GND_net), 
            .I1(n2914), .I2(VCC_net), .I3(n52269), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_12_lut (.I0(GND_net), 
            .I1(n3225), .I2(VCC_net), .I3(n52343), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_14 (.CI(n51369), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n51370));
    SB_LUT4 add_174_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n51368), .O(n1551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_13 (.CI(n51368), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n51369));
    SB_LUT4 i2_4_lut_adj_1798 (.I0(n61896), .I1(n25860), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n62100));
    defparam i2_4_lut_adj_1798.LUT_INIT = 16'hffec;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n51663), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5876), .CO(n51664));
    SB_LUT4 add_174_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n51367), .O(n1552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_13 (.CI(n52185), 
            .I0(n2623), .I1(VCC_net), .CO(n52186));
    SB_CARRY add_262_12 (.CI(n51346), .I0(duty[13]), .I1(n70691), .CO(n51347));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5875), .I3(n51662), .O(displacement_23__N_91[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n51662), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5875), .CO(n51663));
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_6066));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY add_264_5 (.CI(n51316), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n51317));
    SB_LUT4 i2_4_lut_adj_1799 (.I0(delay_counter[22]), .I1(n62100), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_6067));
    defparam i2_4_lut_adj_1799.LUT_INIT = 16'ha8a0;
    SB_LUT4 add_262_11_lut (.I0(current[9]), .I1(duty[12]), .I2(n70691), 
            .I3(n51345), .O(n261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_11_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i29722_4_lut (.I0(n7_adj_6067), .I1(delay_counter[31]), .I2(n25863), 
            .I3(n8_adj_6066), .O(n1642));   // verilog/TinyFPGA_B.v(391[14:38])
    defparam i29722_4_lut.LUT_INIT = 16'h3230;
    SB_CARRY add_264_12 (.CI(n51323), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n51324));
    SB_CARRY add_262_11 (.CI(n51345), .I0(duty[12]), .I1(n70691), .CO(n51346));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1388_3_lut (.I0(n2033), 
            .I1(n2100), .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1455_3_lut (.I0(n2132), 
            .I1(n2199), .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1522_3_lut (.I0(n2231), 
            .I1(n2298), .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1589_3_lut (.I0(n2330), 
            .I1(n2397), .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1656_3_lut (.I0(n2429), 
            .I1(n2496), .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1723_3_lut (.I0(n2528), 
            .I1(n2595), .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1790_3_lut (.I0(n2627), 
            .I1(n2694), .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1857_3_lut (.I0(n2726), 
            .I1(n2793), .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1041_3_lut (.I0(n1526), 
            .I1(n1593), .I2(n1554_adj_5994), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1108_3_lut (.I0(n1625), 
            .I1(n1692), .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1175_3_lut (.I0(n1724), 
            .I1(n1791), .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1242_3_lut (.I0(n1823), 
            .I1(n1890), .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1309_3_lut (.I0(n1922), 
            .I1(n1989), .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1376_3_lut (.I0(n2021), 
            .I1(n2088), .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1443_3_lut (.I0(n2120), 
            .I1(n2187), .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1510_3_lut (.I0(n2219), 
            .I1(n2286), .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1577_3_lut (.I0(n2318), 
            .I1(n2385), .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1644_3_lut (.I0(n2417), 
            .I1(n2484), .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1711_3_lut (.I0(n2516), 
            .I1(n2583), .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_12_lut (.I0(GND_net), 
            .I1(n2624), .I2(VCC_net), .I3(n52184), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5874), .I3(n51661), .O(displacement_23__N_91[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5862));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54285_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70460));
    defparam i54285_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_174_12 (.CI(n51367), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n51368));
    SB_LUT4 i12_4_lut_adj_1800 (.I0(\data_in_frame[20] [2]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[2]), .O(n58244));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1800.LUT_INIT = 16'h3a0a;
    SB_LUT4 i36997_3_lut_4_lut (.I0(n37023), .I1(Ki[2]), .I2(n51273), 
            .I3(n20626), .O(n4_adj_6053));
    defparam i36997_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n51661), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5874), .CO(n51662));
    SB_LUT4 add_174_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n51366), .O(n1553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1801 (.I0(\data_in_frame[20] [1]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[1]), .O(n58248));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1801.LUT_INIT = 16'h3a0a;
    SB_LUT4 n11999_bdd_4_lut_54759 (.I0(n11999), .I1(n430), .I2(current[11]), 
            .I3(duty[23]), .O(n70963));
    defparam n11999_bdd_4_lut_54759.LUT_INIT = 16'he4aa;
    SB_LUT4 add_262_10_lut (.I0(current[8]), .I1(duty[11]), .I2(n70691), 
            .I3(n51344), .O(n262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_10_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_262_10 (.CI(n51344), .I0(duty[11]), .I1(n70691), .CO(n51345));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_12 (.CI(n52184), 
            .I0(n2624), .I1(VCC_net), .CO(n52185));
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n25860));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 dti_counter_2046_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n52631), .O(n38_adj_6015)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR dti_counter_2046__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n28182), 
            .D(n44), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i5_4_lut_adj_1802 (.I0(delay_counter[27]), .I1(delay_counter[26]), 
            .I2(delay_counter[24]), .I3(delay_counter[28]), .O(n12_adj_5998));
    defparam i5_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1803 (.I0(delay_counter[29]), .I1(n12_adj_5998), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25863));
    defparam i6_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i26_3_lut (.I0(encoder0_position_scaled_23__N_319[25]), 
            .I1(n8_adj_5956), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i573_3_lut (.I0(n519), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2112_3_lut (.I0(n3109), 
            .I1(n3176), .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_12 (.CI(n52343), 
            .I0(n3225), .I1(VCC_net), .CO(n52344));
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_6086));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_DFFESR dti_counter_2046__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n28182), 
            .D(n43_adj_6017), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2046__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n28182), 
            .D(n42), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1113_3_lut (.I0(n1630), 
            .I1(n1697), .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2046_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n52630), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7), .I3(n51660), .O(displacement_23__N_91[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2046_add_4_8 (.CI(n52630), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n52631));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_22 (.CI(n52269), 
            .I0(n2914), .I1(VCC_net), .CO(n52270));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_11_lut (.I0(GND_net), 
            .I1(n2625), .I2(VCC_net), .I3(n52183), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n51660), .I0(encoder0_position_scaled[18]), 
            .I1(n7), .CO(n51661));
    SB_LUT4 dti_counter_2046_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n52629), .O(n40_adj_6016)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_11 (.CI(n51366), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n51367));
    SB_CARRY dti_counter_2046_add_4_7 (.CI(n52629), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n52630));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_11_lut (.I0(GND_net), 
            .I1(n3226), .I2(VCC_net), .I3(n52342), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n51365), .O(n1554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_10 (.CI(n51365), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n51366));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8), .I3(n51659), .O(displacement_23__N_91[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n51659), .I0(encoder0_position_scaled[17]), 
            .I1(n8), .CO(n51660));
    SB_LUT4 i1_2_lut_adj_1804 (.I0(n42166), .I1(n8_adj_5973), .I2(GND_net), 
            .I3(GND_net), .O(n28774));
    defparam i1_2_lut_adj_1804.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1805 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_6084));
    defparam i6_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_11 (.CI(n52183), 
            .I0(n2625), .I1(VCC_net), .CO(n52184));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9), .I3(n51658), .O(displacement_23__N_91[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n15_adj_6084), .I1(delay_counter[2]), .I2(n14_adj_6086), 
            .I3(delay_counter[6]), .O(n25840));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n70963_bdd_4_lut (.I0(n70963), .I1(duty[11]), .I2(n259), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[11]));
    defparam n70963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_10_lut (.I0(GND_net), 
            .I1(n2626), .I2(VCC_net), .I3(n52182), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n51658), .I0(encoder0_position_scaled[16]), 
            .I1(n9), .CO(n51659));
    SB_LUT4 add_174_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n51364), .O(n1555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_9 (.CI(n51364), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n51365));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_21_lut (.I0(GND_net), 
            .I1(n2915), .I2(VCC_net), .I3(n52268), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4958_4_lut (.I0(n25840), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5996));
    defparam i4958_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1180_3_lut (.I0(n1729), 
            .I1(n1796), .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR dti_counter_2046__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n28182), 
            .D(n41), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i2_4_lut_adj_1806 (.I0(n24_adj_5996), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n60932));
    defparam i2_4_lut_adj_1806.LUT_INIT = 16'hc800;
    SB_LUT4 i12_4_lut_adj_1807 (.I0(\data_in_frame[20] [0]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[0]), .O(n58252));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1807.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_21 (.CI(n52268), 
            .I0(n2915), .I1(VCC_net), .CO(n52269));
    SB_LUT4 dti_counter_2046_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n52628), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_10 (.CI(n52182), 
            .I0(n2626), .I1(VCC_net), .CO(n52183));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1778_3_lut (.I0(n2615), 
            .I1(n2682), .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_11 (.CI(n52342), 
            .I0(n3226), .I1(VCC_net), .CO(n52343));
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_9_lut (.I0(GND_net), 
            .I1(n2627), .I2(VCC_net), .I3(n52181), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_10_lut (.I0(GND_net), 
            .I1(n3227), .I2(VCC_net), .I3(n52341), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(delay_counter[22]), .I1(delay_counter[21]), 
            .I2(n25863), .I3(delay_counter[23]), .O(n4_adj_6018));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_20_lut (.I0(GND_net), 
            .I1(n2916), .I2(VCC_net), .I3(n52267), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1809 (.I0(n60932), .I1(delay_counter[18]), .I2(n25860), 
            .I3(GND_net), .O(n62096));
    defparam i2_3_lut_adj_1809.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_9 (.CI(n52181), 
            .I0(n2627), .I1(VCC_net), .CO(n52182));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_10 (.CI(n52341), 
            .I0(n3227), .I1(VCC_net), .CO(n52342));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_8_lut (.I0(GND_net), 
            .I1(n2628), .I2(VCC_net), .I3(n52180), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n51363), .O(n1556)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5842), .I3(n51657), .O(displacement_23__N_91[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_8 (.CI(n52180), 
            .I0(n2628), .I1(VCC_net), .CO(n52181));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n51657), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5842), .CO(n51658));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5882), .I3(n51656), .O(displacement_23__N_91[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_7_lut (.I0(GND_net), 
            .I1(n2629), .I2(GND_net), .I3(n52179), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2046_add_4_6 (.CI(n52628), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n52629));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_7 (.CI(n52179), 
            .I0(n2629), .I1(GND_net), .CO(n52180));
    SB_LUT4 i43762_3_lut (.I0(n5_adj_5959), .I1(n7906), .I2(n59878), .I3(GND_net), 
            .O(n59883));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2046_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n52627), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16180_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n23164), .I3(GND_net), .O(n30587));   // verilog/coms.v(130[12] 305[6])
    defparam i16180_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n17_adj_6070));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1247_3_lut (.I0(n1828), 
            .I1(n1895), .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_20 (.CI(n52267), 
            .I0(n2916), .I1(VCC_net), .CO(n52268));
    SB_LUT4 i2_4_lut_adj_1810 (.I0(n62096), .I1(n4_adj_6018), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n62_adj_5997));
    defparam i2_4_lut_adj_1810.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_9_lut (.I0(GND_net), 
            .I1(n3228), .I2(VCC_net), .I3(n52340), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_19_lut (.I0(GND_net), 
            .I1(n2917), .I2(VCC_net), .I3(n52266), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11999_bdd_4_lut_54739 (.I0(n11999), .I1(n431), .I2(current[10]), 
            .I3(duty[23]), .O(n70957));
    defparam n11999_bdd_4_lut_54739.LUT_INIT = 16'he4aa;
    SB_LUT4 n70957_bdd_4_lut (.I0(n70957), .I1(duty[10]), .I2(n260), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[10]));
    defparam n70957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1314_3_lut (.I0(n1927), 
            .I1(n1994), .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_6_lut (.I0(GND_net), 
            .I1(n2630), .I2(GND_net), .I3(n52178), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_8 (.CI(n51363), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n51364));
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY dti_counter_2046_add_4_5 (.CI(n52627), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n52628));
    SB_LUT4 add_262_9_lut (.I0(current[7]), .I1(duty[10]), .I2(n70691), 
            .I3(n51343), .O(n263)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_174_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n51362), .O(n1557)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_7 (.CI(n51362), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n51363));
    SB_LUT4 add_174_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n51361), .O(n1558)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_6 (.CI(n51361), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n51362));
    SB_LUT4 add_174_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n51360), .O(n1559)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54258_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70433));
    defparam i54258_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_19 (.CI(n52266), 
            .I0(n2917), .I1(VCC_net), .CO(n52267));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_18_lut (.I0(GND_net), 
            .I1(n2918), .I2(VCC_net), .I3(n52265), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_5 (.CI(n51360), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n51361));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n51656), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5882), .CO(n51657));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_18 (.CI(n52265), 
            .I0(n2918), .I1(VCC_net), .CO(n52266));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_17_lut (.I0(GND_net), 
            .I1(n2919), .I2(VCC_net), .I3(n52264), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n51359), .O(n1560)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11999_bdd_4_lut_54734 (.I0(n11999), .I1(n432), .I2(current[9]), 
            .I3(duty[23]), .O(n70951));
    defparam n11999_bdd_4_lut_54734.LUT_INIT = 16'he4aa;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 dti_counter_2046_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n52626), .O(n43_adj_6017)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5861));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5881), .I3(n51655), .O(displacement_23__N_91[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_4 (.CI(n51359), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n51360));
    SB_LUT4 i43763_3_lut (.I0(encoder0_position_scaled_23__N_319[28]), .I1(n59883), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n70951_bdd_4_lut (.I0(n70951), .I1(duty[9]), .I2(n261), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n70951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY dti_counter_2046_add_4_4 (.CI(n52626), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n52627));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n51655), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5881), .CO(n51656));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_262_9 (.CI(n51343), .I0(duty[10]), .I1(n70691), .CO(n51344));
    SB_LUT4 i16159_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n59086), .I3(GND_net), .O(n30566));   // verilog/coms.v(130[12] 305[6])
    defparam i16159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2046_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n52625), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29721_2_lut (.I0(n62_adj_5997), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_522));   // verilog/TinyFPGA_B.v(377[12:35])
    defparam i29721_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i623_2_lut (.I0(n1642), .I1(n43842), .I2(GND_net), .I3(GND_net), 
            .O(n3305));   // verilog/TinyFPGA_B.v(395[18] 397[12])
    defparam i623_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_351));   // verilog/TinyFPGA_B.v(325[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_17 (.CI(n52264), 
            .I0(n2919), .I1(VCC_net), .CO(n52265));
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16155_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n59086), .I3(GND_net), .O(n30562));   // verilog/coms.v(130[12] 305[6])
    defparam i16155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15377_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n78), .I3(GND_net), .O(n29784));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5860));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16667_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [1]), 
            .O(n31074));   // verilog/coms.v(130[12] 305[6])
    defparam i16667_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16151_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n59086), .I3(GND_net), .O(n30558));   // verilog/coms.v(130[12] 305[6])
    defparam i16151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48036_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64201));
    defparam i48036_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54119_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70294));
    defparam i54119_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_9 (.CI(n52340), 
            .I0(n3228), .I1(VCC_net), .CO(n52341));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5880), .I3(n51654), .O(displacement_23__N_91[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54481_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7082), .I2(n64201), 
            .I3(n25_adj_6071), .O(n17_adj_6070));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i54481_4_lut.LUT_INIT = 16'h88ba;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_6 (.CI(n52178), 
            .I0(n2630), .I1(GND_net), .CO(n52179));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1381_3_lut (.I0(n2026), 
            .I1(n2093), .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16147_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n59086), .I3(GND_net), .O(n30554));   // verilog/coms.v(130[12] 305[6])
    defparam i16147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1811 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[16] [7]), .I3(GND_net), .O(n59138));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1811.LUT_INIT = 16'h9696;
    SB_LUT4 i16143_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n59086), .I3(GND_net), .O(n30550));   // verilog/coms.v(130[12] 305[6])
    defparam i16143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1812 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_264));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_3_lut_adj_1812.LUT_INIT = 16'h0202;
    SB_LUT4 i4_4_lut (.I0(n7_adj_6064), .I1(\data_in_frame[12] [3]), .I2(n54986), 
            .I3(n59499), .O(n25605));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_6090));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1813 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_256[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1813.LUT_INIT = 16'h1414;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_adj_1814 (.I0(\data_in_frame[14] [5]), .I1(n26902), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5847));
    defparam i1_2_lut_adj_1814.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1815 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [4]), 
            .I2(n54986), .I3(n6_adj_5847), .O(n61411));
    defparam i4_4_lut_adj_1815.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1816 (.I0(n2023), .I1(n2027), .I2(n2024), .I3(GND_net), 
            .O(n63478));
    defparam i1_3_lut_adj_1816.LUT_INIT = 16'hfefe;
    SB_LUT4 i16755_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [0]), 
            .O(n31162));   // verilog/coms.v(130[12] 305[6])
    defparam i16755_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1448_3_lut (.I0(n2125), 
            .I1(n2192), .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30395_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n44695));
    defparam i30395_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1515_3_lut (.I0(n2224), 
            .I1(n2291), .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n2021), .I1(n2022), .I2(n63478), .I3(n63476), 
            .O(n63484));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 n11999_bdd_4_lut_54729 (.I0(n11999), .I1(n433), .I2(current[8]), 
            .I3(duty[23]), .O(n70945));
    defparam n11999_bdd_4_lut_54729.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1582_3_lut (.I0(n2323), 
            .I1(n2390), .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1649_3_lut (.I0(n2422), 
            .I1(n2489), .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n2029), .I1(n44695), .I2(n2030), .I3(n2031), 
            .O(n60781));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'ha080;
    SB_CARRY dti_counter_2046_add_4_3 (.CI(n52625), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n52626));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n51654), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5880), .CO(n51655));
    SB_LUT4 dti_counter_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_5_lut (.I0(GND_net), 
            .I1(n2631), .I2(VCC_net), .I3(n52177), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5879), .I3(n51653), .O(displacement_23__N_91[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_16_lut (.I0(GND_net), 
            .I1(n2920), .I2(VCC_net), .I3(n52263), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1716_3_lut (.I0(n2521), 
            .I1(n2588), .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1783_3_lut (.I0(n2620), 
            .I1(n2687), .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n52625));
    SB_LUT4 i54407_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70582));
    defparam i54407_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5882));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n2019), .I1(n60781), .I2(n2020), .I3(n63484), 
            .O(n63490));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i15809_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n59079), 
            .I3(GND_net), .O(n30216));   // verilog/coms.v(130[12] 305[6])
    defparam i15809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5859));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n51653), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5879), .CO(n51654));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_8_lut (.I0(GND_net), 
            .I1(n3229), .I2(GND_net), .I3(n52339), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_16 (.CI(n52263), 
            .I0(n2920), .I1(VCC_net), .CO(n52264));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_5 (.CI(n52177), 
            .I0(n2631), .I1(VCC_net), .CO(n52178));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5848), .I3(n51652), .O(displacement_23__N_91[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_174_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n51358), .O(n1561)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_15_lut (.I0(GND_net), 
            .I1(n2921), .I2(VCC_net), .I3(n52262), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16668_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [2]), 
            .O(n31075));   // verilog/coms.v(130[12] 305[6])
    defparam i16668_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5858));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_4_lut (.I0(GND_net), 
            .I1(n2632), .I2(GND_net), .I3(n52176), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5842));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_115[10]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i11_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_15 (.CI(n52262), 
            .I0(n2921), .I1(VCC_net), .CO(n52263));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_20_lut (.I0(n70433), 
            .I1(n2016), .I2(VCC_net), .I3(n52047), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_174_3 (.CI(n51358), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n51359));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_4 (.CI(n52176), 
            .I0(n2632), .I1(GND_net), .CO(n52177));
    SB_LUT4 add_174_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1562)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_8_lut (.I0(current[6]), .I1(duty[9]), .I2(n70691), 
            .I3(n51342), .O(n264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_15_lut (.I0(n70548), 
            .I1(n1521), .I2(VCC_net), .I3(n51855), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_3_lut (.I0(GND_net), 
            .I1(n2633), .I2(VCC_net), .I3(n52175), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_3 (.CI(n52175), 
            .I0(n2633), .I1(VCC_net), .CO(n52176));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n51652), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5848), .CO(n51653));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_14_lut (.I0(GND_net), 
            .I1(n2922), .I2(VCC_net), .I3(n52261), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1773_3_lut (.I0(n2610), 
            .I1(n2677), .I2(n2643), .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16108_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n59975), .I3(GND_net), .O(n30515));   // verilog/coms.v(130[12] 305[6])
    defparam i16108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15812_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n59079), 
            .I3(GND_net), .O(n30219));   // verilog/coms.v(130[12] 305[6])
    defparam i15812_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16105_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n59975), .I3(GND_net), .O(n30512));   // verilog/coms.v(130[12] 305[6])
    defparam i16105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15815_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n59079), 
            .I3(GND_net), .O(n30222));   // verilog/coms.v(130[12] 305[6])
    defparam i15815_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_8 (.CI(n52339), 
            .I0(n3229), .I1(GND_net), .CO(n52340));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5926), .I3(n51651), .O(displacement_23__N_91[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16102_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n59975), .I3(GND_net), .O(n30509));   // verilog/coms.v(130[12] 305[6])
    defparam i16102_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_14 (.CI(n52261), 
            .I0(n2922), .I1(VCC_net), .CO(n52262));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_19_lut (.I0(GND_net), 
            .I1(n2017), .I2(VCC_net), .I3(n52046), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_13_lut (.I0(GND_net), 
            .I1(n2923), .I2(VCC_net), .I3(n52260), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_14_lut (.I0(GND_net), 
            .I1(n1522), .I2(VCC_net), .I3(n51854), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n51358));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1771_2_lut (.I0(GND_net), 
            .I1(n951), .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n51651), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5926), .CO(n51652));
    SB_LUT4 add_262_23_lut (.I0(current[15]), .I1(duty[23]), .I2(n70691), 
            .I3(n51357), .O(n249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_23_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2131_3_lut (.I0(n3128), 
            .I1(n3195), .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_7_lut (.I0(n3298), 
            .I1(n3230), .I2(GND_net), .I3(n52338), .O(n67030)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1771_2 (.CI(VCC_net), 
            .I0(n951), .I1(GND_net), .CO(n52175));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_19 (.CI(n52046), 
            .I0(n2017), .I1(VCC_net), .CO(n52047));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5925), .I3(n51650), .O(displacement_23__N_91[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_22_lut (.I0(current[15]), .I1(duty[23]), .I2(n70691), 
            .I3(n51356), .O(n250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_22_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_262_22 (.CI(n51356), .I0(duty[23]), .I1(n70691), .CO(n51357));
    SB_LUT4 i14808_2_lut (.I0(n28059), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14808_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53720_4_lut (.I0(commutation_state[1]), .I1(n23298), .I2(dti), 
            .I3(commutation_state[2]), .O(n28059));
    defparam i53720_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i53722_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[12] [4]), 
            .I2(n59975), .I3(GND_net), .O(n58398));   // verilog/coms.v(94[13:20])
    defparam i53722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53721_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[12] [3]), 
            .I2(n59975), .I3(GND_net), .O(n58384));   // verilog/coms.v(94[13:20])
    defparam i53721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16092_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n59975), .I3(GND_net), .O(n30499));   // verilog/coms.v(130[12] 305[6])
    defparam i16092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16088_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n59975), .I3(GND_net), .O(n30495));   // verilog/coms.v(130[12] 305[6])
    defparam i16088_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_14 (.CI(n51854), 
            .I0(n1522), .I1(VCC_net), .CO(n51855));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_18_lut (.I0(GND_net), 
            .I1(n2018), .I2(VCC_net), .I3(n52045), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_13 (.CI(n52260), 
            .I0(n2923), .I1(VCC_net), .CO(n52261));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_25_lut (.I0(n70372), 
            .I1(n2511), .I2(VCC_net), .I3(n52174), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_13_lut (.I0(GND_net), 
            .I1(n1523), .I2(VCC_net), .I3(n51853), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_13 (.CI(n51853), 
            .I0(n1523), .I1(VCC_net), .CO(n51854));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_24_lut (.I0(GND_net), 
            .I1(n2512), .I2(VCC_net), .I3(n52173), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_18 (.CI(n52045), 
            .I0(n2018), .I1(VCC_net), .CO(n52046));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_12_lut (.I0(GND_net), 
            .I1(n1524), .I2(VCC_net), .I3(n51852), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n51650), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5925), .CO(n51651));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_17_lut (.I0(GND_net), 
            .I1(n2019), .I2(VCC_net), .I3(n52044), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16085_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n59975), .I3(GND_net), .O(n30492));   // verilog/coms.v(130[12] 305[6])
    defparam i16085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5924), .I3(n51649), .O(displacement_23__N_91[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_12 (.CI(n51852), 
            .I0(n1524), .I1(VCC_net), .CO(n51853));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n51649), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5924), .CO(n51650));
    SB_LUT4 mux_277_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_115[11]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_11_lut (.I0(GND_net), 
            .I1(n1525), .I2(VCC_net), .I3(n51851), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5923), .I3(n51648), .O(displacement_23__N_91[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_24 (.CI(n52173), 
            .I0(n2512), .I1(VCC_net), .CO(n52174));
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5857));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1039_3_lut (.I0(n1524), 
            .I1(n1591), .I2(n1554_adj_5994), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_277_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_115[12]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_19_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16082_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n28791), .I3(GND_net), .O(n30489));   // verilog/coms.v(130[12] 305[6])
    defparam i16082_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16078_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n28791), .I3(GND_net), .O(n30485));   // verilog/coms.v(130[12] 305[6])
    defparam i16078_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_11 (.CI(n51851), 
            .I0(n1525), .I1(VCC_net), .CO(n51852));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n51648), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5923), .CO(n51649));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_17 (.CI(n52044), 
            .I0(n2019), .I1(VCC_net), .CO(n52045));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_23_lut (.I0(GND_net), 
            .I1(n2513), .I2(VCC_net), .I3(n52172), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_10_lut (.I0(GND_net), 
            .I1(n1526), .I2(VCC_net), .I3(n51850), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_10 (.CI(n51850), 
            .I0(n1526), .I1(VCC_net), .CO(n51851));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_9_lut (.I0(GND_net), 
            .I1(n1527), .I2(VCC_net), .I3(n51849), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_12_lut (.I0(GND_net), 
            .I1(n2924), .I2(VCC_net), .I3(n52259), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_16_lut (.I0(GND_net), 
            .I1(n2020), .I2(VCC_net), .I3(n52043), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5922), .I3(n51647), .O(displacement_23__N_91[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_9 (.CI(n51849), 
            .I0(n1527), .I1(VCC_net), .CO(n51850));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n51647), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5922), .CO(n51648));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_8_lut (.I0(GND_net), 
            .I1(n1528), .I2(VCC_net), .I3(n51848), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_23 (.CI(n52172), 
            .I0(n2513), .I1(VCC_net), .CO(n52173));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_8 (.CI(n51848), 
            .I0(n1528), .I1(VCC_net), .CO(n51849));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1106_3_lut (.I0(n1623), 
            .I1(n1690), .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16075_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n28791), .I3(GND_net), .O(n30482));   // verilog/coms.v(130[12] 305[6])
    defparam i16075_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_12 (.CI(n52259), 
            .I0(n2924), .I1(VCC_net), .CO(n52260));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_16 (.CI(n52043), 
            .I0(n2020), .I1(VCC_net), .CO(n52044));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1173_3_lut (.I0(n1722), 
            .I1(n1789), .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i27_3_lut (.I0(encoder0_position_scaled_23__N_319[26]), 
            .I1(n7_adj_5957), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5873));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5872));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_15_lut (.I0(GND_net), 
            .I1(n2021), .I2(VCC_net), .I3(n52042), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_11_lut (.I0(GND_net), 
            .I1(n2925), .I2(VCC_net), .I3(n52258), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_7 (.CI(n52338), 
            .I0(n3230), .I1(GND_net), .CO(n52339));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5921), .I3(n51646), .O(displacement_23__N_91[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n51646), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5921), .CO(n51647));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_7_lut (.I0(GND_net), 
            .I1(n1529), .I2(GND_net), .I3(n51847), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_22_lut (.I0(GND_net), 
            .I1(n2514), .I2(VCC_net), .I3(n52171), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_22 (.CI(n52171), 
            .I0(n2514), .I1(VCC_net), .CO(n52172));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_21_lut (.I0(GND_net), 
            .I1(n2515), .I2(VCC_net), .I3(n52170), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_15 (.CI(n52042), 
            .I0(n2021), .I1(VCC_net), .CO(n52043));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_14_lut (.I0(GND_net), 
            .I1(n2022), .I2(VCC_net), .I3(n52041), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_14 (.CI(n52041), 
            .I0(n2022), .I1(VCC_net), .CO(n52042));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_11 (.CI(n52258), 
            .I0(n2925), .I1(VCC_net), .CO(n52259));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_7 (.CI(n51847), 
            .I0(n1529), .I1(GND_net), .CO(n51848));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_6_lut (.I0(GND_net), 
            .I1(n1530), .I2(GND_net), .I3(n51846), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n70945_bdd_4_lut (.I0(n70945), .I1(duty[8]), .I2(n262), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n70945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_19_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5871));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_10_lut (.I0(GND_net), 
            .I1(n2926), .I2(VCC_net), .I3(n52257), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5870));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30211_2_lut (.I0(duty[15]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5441));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30211_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i16072_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n28791), .I3(GND_net), .O(n30479));   // verilog/coms.v(130[12] 305[6])
    defparam i16072_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5869));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5856));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5868));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16068_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n28791), .I3(GND_net), .O(n30475));   // verilog/coms.v(130[12] 305[6])
    defparam i16068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15818_3_lut (.I0(\data_in_frame[2] [4]), .I1(rx_data[4]), .I2(n59079), 
            .I3(GND_net), .O(n30225));   // verilog/coms.v(130[12] 305[6])
    defparam i15818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54424_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70599));
    defparam i54424_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_21 (.CI(n52170), 
            .I0(n2515), .I1(VCC_net), .CO(n52171));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_13_lut (.I0(GND_net), 
            .I1(n2023), .I2(VCC_net), .I3(n52040), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22669_3_lut (.I0(n28791), .I1(rx_data[2]), .I2(\data_in_frame[11] [2]), 
            .I3(GND_net), .O(n30616));   // verilog/coms.v(94[13:20])
    defparam i22669_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_13 (.CI(n52040), 
            .I0(n2023), .I1(VCC_net), .CO(n52041));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_20_lut (.I0(GND_net), 
            .I1(n2516), .I2(VCC_net), .I3(n52169), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_6 (.CI(n51846), 
            .I0(n1530), .I1(GND_net), .CO(n51847));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1240_3_lut (.I0(n1821), 
            .I1(n1888), .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_5_lut (.I0(GND_net), 
            .I1(n1531_adj_5991), .I2(VCC_net), .I3(n51845), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1863_3_lut (.I0(n2732), 
            .I1(n2799), .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_5 (.CI(n51845), 
            .I0(n1531_adj_5991), .I1(VCC_net), .CO(n51846));
    SB_LUT4 i16062_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n28791), .I3(GND_net), .O(n30469));   // verilog/coms.v(130[12] 305[6])
    defparam i16062_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_20 (.CI(n52169), 
            .I0(n2516), .I1(VCC_net), .CO(n52170));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_12_lut (.I0(GND_net), 
            .I1(n2024), .I2(VCC_net), .I3(n52039), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_6_lut (.I0(GND_net), 
            .I1(n3231), .I2(VCC_net), .I3(n52337), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_4_lut (.I0(GND_net), 
            .I1(n1532_adj_5992), .I2(GND_net), .I3(n51844), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5920), .I3(n51645), .O(displacement_23__N_91[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_10 (.CI(n52257), 
            .I0(n2926), .I1(VCC_net), .CO(n52258));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_9_lut (.I0(GND_net), 
            .I1(n2927), .I2(VCC_net), .I3(n52256), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_9 (.CI(n52256), 
            .I0(n2927), .I1(VCC_net), .CO(n52257));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_4 (.CI(n51844), 
            .I0(n1532_adj_5992), .I1(GND_net), .CO(n51845));
    SB_LUT4 add_262_21_lut (.I0(current[15]), .I1(duty[22]), .I2(n70691), 
            .I3(n51355), .O(n251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_21_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_6 (.CI(n52337), 
            .I0(n3231), .I1(VCC_net), .CO(n52338));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1307_3_lut (.I0(n1920), 
            .I1(n1987), .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1374_3_lut (.I0(n2019), 
            .I1(n2086), .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1441_3_lut (.I0(n2118), 
            .I1(n2185), .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1508_3_lut (.I0(n2217), 
            .I1(n2284), .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2130_3_lut (.I0(n3127), 
            .I1(n3194), .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_19_lut (.I0(GND_net), 
            .I1(n2517), .I2(VCC_net), .I3(n52168), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n51645), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5920), .CO(n51646));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_3_lut (.I0(GND_net), 
            .I1(n1533_adj_5993), .I2(VCC_net), .I3(n51843), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_12 (.CI(n52039), 
            .I0(n2024), .I1(VCC_net), .CO(n52040));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_5_lut (.I0(GND_net), 
            .I1(n3232), .I2(GND_net), .I3(n52336), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5919), .I3(n51644), .O(displacement_23__N_91[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_19 (.CI(n52168), 
            .I0(n2517), .I1(VCC_net), .CO(n52169));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1575_3_lut (.I0(n2316), 
            .I1(n2383), .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16059_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n28791), .I3(GND_net), .O(n30466));   // verilog/coms.v(130[12] 305[6])
    defparam i16059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_277_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_115[14]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_282_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_115[15]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_8_lut (.I0(GND_net), 
            .I1(n2928), .I2(VCC_net), .I3(n52255), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_3 (.CI(n51843), 
            .I0(n1533_adj_5993), .I1(VCC_net), .CO(n51844));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1034_2_lut (.I0(GND_net), 
            .I1(n940), .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n51644), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5919), .CO(n51645));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_5 (.CI(n52336), 
            .I0(n3232), .I1(GND_net), .CO(n52337));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_18_lut (.I0(GND_net), 
            .I1(n2518), .I2(VCC_net), .I3(n52167), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_18 (.CI(n52167), 
            .I0(n2518), .I1(VCC_net), .CO(n52168));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_8 (.CI(n52255), 
            .I0(n2928), .I1(VCC_net), .CO(n52256));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1034_2 (.CI(VCC_net), 
            .I0(n940), .I1(GND_net), .CO(n51843));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_11_lut (.I0(GND_net), 
            .I1(n2025), .I2(VCC_net), .I3(n52038), .O(n2092_adj_5995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1642_3_lut (.I0(n2415), 
            .I1(n2482), .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54352_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70527));
    defparam i54352_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_262_21 (.CI(n51355), .I0(duty[22]), .I1(n70691), .CO(n51356));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_11 (.CI(n52038), 
            .I0(n2025), .I1(VCC_net), .CO(n52039));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_10_lut (.I0(GND_net), 
            .I1(n2026), .I2(VCC_net), .I3(n52037), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5918), .I3(n51643), .O(displacement_23__N_91[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_20_lut (.I0(current[15]), .I1(duty[21]), .I2(n70691), 
            .I3(n51354), .O(n252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_20_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_7_lut (.I0(GND_net), 
            .I1(n2929), .I2(GND_net), .I3(n52254), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_7 (.CI(n52254), 
            .I0(n2929), .I1(GND_net), .CO(n52255));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_4_lut (.I0(GND_net), 
            .I1(n3233), .I2(VCC_net), .I3(n52335), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_17_lut (.I0(GND_net), 
            .I1(n2519), .I2(VCC_net), .I3(n52166), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_10 (.CI(n52037), 
            .I0(n2026), .I1(VCC_net), .CO(n52038));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n51643), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5918), .CO(n51644));
    SB_LUT4 i15821_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n59079), 
            .I3(GND_net), .O(n30228));   // verilog/coms.v(130[12] 305[6])
    defparam i15821_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15824_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n78), .I3(GND_net), .O(n30231));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15824_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_17 (.CI(n52166), 
            .I0(n2519), .I1(VCC_net), .CO(n52167));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5917), .I3(VCC_net), .O(displacement_23__N_91[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_9_lut (.I0(GND_net), 
            .I1(n2027), .I2(VCC_net), .I3(n52036), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5917), .CO(n51643));
    SB_CARRY add_262_20 (.CI(n51354), .I0(duty[21]), .I1(n70691), .CO(n51355));
    SB_LUT4 unary_minus_19_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5867));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1709_3_lut (.I0(n2514), 
            .I1(n2581), .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54373_1_lut (.I0(n1554_adj_5994), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n70548));
    defparam i54373_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1125_25_lut (.I0(GND_net), .I1(n5409), .I2(n5433), .I3(n51642), 
            .O(n418)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5855));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_9 (.CI(n52036), 
            .I0(n2027), .I1(VCC_net), .CO(n52037));
    SB_LUT4 unary_minus_19_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5866));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1776_3_lut (.I0(n2613), 
            .I1(n2680), .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54395_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70570));
    defparam i54395_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_1125_24_lut (.I0(GND_net), .I1(n5409), .I2(n5434), .I3(n51641), 
            .O(n419)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_19_lut (.I0(current[15]), .I1(duty[20]), .I2(n70691), 
            .I3(n51353), .O(n253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_19_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_16_lut (.I0(GND_net), 
            .I1(n2520), .I2(VCC_net), .I3(n52165), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_16 (.CI(n52165), 
            .I0(n2520), .I1(VCC_net), .CO(n52166));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_8_lut (.I0(GND_net), 
            .I1(n2028), .I2(VCC_net), .I3(n52035), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_8 (.CI(n52035), 
            .I0(n2028), .I1(VCC_net), .CO(n52036));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_4 (.CI(n52335), 
            .I0(n3233), .I1(VCC_net), .CO(n52336));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_3_lut (.I0(GND_net), 
            .I1(n957), .I2(GND_net), .I3(n52334), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_6_lut (.I0(GND_net), 
            .I1(n2930), .I2(GND_net), .I3(n52253), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5865));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54454_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70629));
    defparam i54454_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_262_19 (.CI(n51353), .I0(duty[20]), .I1(n70691), .CO(n51354));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_7_lut (.I0(GND_net), 
            .I1(n2029), .I2(GND_net), .I3(n52034), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_6 (.CI(n52253), 
            .I0(n2930), .I1(GND_net), .CO(n52254));
    SB_CARRY add_1125_24 (.CI(n51641), .I0(n5409), .I1(n5434), .CO(n51642));
    SB_LUT4 add_262_18_lut (.I0(current[15]), .I1(duty[19]), .I2(n70691), 
            .I3(n51352), .O(n254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_18_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 unary_minus_19_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5864));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1843_3_lut (.I0(n2712), 
            .I1(n2779), .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5854));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_19_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5863));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_19_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_277_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_115[16]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_15_lut (.I0(GND_net), 
            .I1(n2521), .I2(VCC_net), .I3(n52164), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_15 (.CI(n52164), 
            .I0(n2521), .I1(VCC_net), .CO(n52165));
    SB_LUT4 add_1125_23_lut (.I0(GND_net), .I1(n5409), .I2(n5435), .I3(n51640), 
            .O(n420)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_262_18 (.CI(n51352), .I0(duty[19]), .I1(n70691), .CO(n51353));
    SB_LUT4 add_264_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n51322), .O(encoder1_position_scaled_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_14_lut (.I0(GND_net), 
            .I1(n2522), .I2(VCC_net), .I3(n52163), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_7 (.CI(n52034), 
            .I0(n2029), .I1(GND_net), .CO(n52035));
    SB_LUT4 i54467_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n70642));
    defparam i54467_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position_scaled_23__N_319[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_6019));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5874));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1125_23 (.CI(n51640), .I0(n5409), .I1(n5435), .CO(n51641));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_3 (.CI(n52334), 
            .I0(n957), .I1(GND_net), .CO(n52335));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_14 (.CI(n52163), 
            .I0(n2522), .I1(VCC_net), .CO(n52164));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1452_3_lut (.I0(n2129), 
            .I1(n2196), .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43764_3_lut (.I0(n6_adj_5958), .I1(n7907), .I2(n59878), .I3(GND_net), 
            .O(n59885));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1125_22_lut (.I0(GND_net), .I1(n5411), .I2(n5436), .I3(n51639), 
            .O(n421)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_5_lut (.I0(GND_net), 
            .I1(n2931), .I2(VCC_net), .I3(n52252), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2173_2 (.CI(VCC_net), 
            .I0(n652), .I1(VCC_net), .CO(n52334));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1519_3_lut (.I0(n2228), 
            .I1(n2295), .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i43765_3_lut (.I0(encoder0_position_scaled_23__N_319[27]), .I1(n59885), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1586_3_lut (.I0(n2327), 
            .I1(n2394), .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_6_lut (.I0(GND_net), 
            .I1(n2030), .I2(GND_net), .I3(n52033), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_31_lut (.I0(n70089), 
            .I1(n3105), .I2(VCC_net), .I3(n52333), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1125_22 (.CI(n51639), .I0(n5411), .I1(n5436), .CO(n51640));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_30_lut (.I0(GND_net), 
            .I1(n3106), .I2(VCC_net), .I3(n52332), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR dti_counter_2046__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n28182), 
            .D(n40_adj_6016), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1653_3_lut (.I0(n2426), 
            .I1(n2493), .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1720_3_lut (.I0(n2525), 
            .I1(n2592), .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_30 (.CI(n52332), 
            .I0(n3106), .I1(VCC_net), .CO(n52333));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_13_lut (.I0(GND_net), 
            .I1(n2523), .I2(VCC_net), .I3(n52162), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_6 (.CI(n52033), 
            .I0(n2030), .I1(GND_net), .CO(n52034));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_5_lut (.I0(GND_net), 
            .I1(n2031), .I2(VCC_net), .I3(n52032), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_5 (.CI(n52032), 
            .I0(n2031), .I1(VCC_net), .CO(n52033));
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFESR dti_counter_2046__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n28182), 
            .D(n39), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2046__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n28182), 
            .D(n38_adj_6015), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 add_1125_21_lut (.I0(GND_net), .I1(n5412), .I2(n5437), .I3(n51638), 
            .O(n422)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_21 (.CI(n51638), .I0(n5412), .I1(n5437), .CO(n51639));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5875));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15825_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n78), .I3(GND_net), .O(n30232));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15825_3_lut.LUT_INIT = 16'hacac;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_4_lut (.I0(GND_net), 
            .I1(n2032), .I2(GND_net), .I3(n52031), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_5 (.CI(n52252), 
            .I0(n2931), .I1(VCC_net), .CO(n52253));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_13 (.CI(n52162), 
            .I0(n2523), .I1(VCC_net), .CO(n52163));
    SB_LUT4 i15826_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n78), .I3(GND_net), .O(n30233));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2129_3_lut (.I0(n3126), 
            .I1(n3193), .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5876));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_12_lut (.I0(GND_net), 
            .I1(n2524), .I2(VCC_net), .I3(n52161), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5877));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_4_lut (.I0(GND_net), 
            .I1(n2932), .I2(GND_net), .I3(n52251), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_282_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_115[17]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i705_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i16006_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n59971), 
            .I3(GND_net), .O(n30413));   // verilog/coms.v(130[12] 305[6])
    defparam i16006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16002_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n59971), 
            .I3(GND_net), .O(n30409));   // verilog/coms.v(130[12] 305[6])
    defparam i16002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5878));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15999_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n59971), 
            .I3(GND_net), .O(n30406));   // verilog/coms.v(130[12] 305[6])
    defparam i15999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2128_3_lut (.I0(n3125), 
            .I1(n3192), .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16231_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n23164), .I3(GND_net), .O(n30638));   // verilog/coms.v(130[12] 305[6])
    defparam i16231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16232_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n23164), .I3(GND_net), .O(n30639));   // verilog/coms.v(130[12] 305[6])
    defparam i16232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_282_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_115[18]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15827_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n78), .I3(GND_net), .O(n30234));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15827_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15996_3_lut (.I0(\data_in_frame[8] [4]), .I1(rx_data[4]), .I2(n59971), 
            .I3(GND_net), .O(n30403));   // verilog/coms.v(130[12] 305[6])
    defparam i15996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_282_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_277_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_115[19]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i20_3_lut.LUT_INIT = 16'h3535;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i15828_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n78), .I3(GND_net), .O(n30235));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15828_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i15384_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n62864), 
            .I3(n27_adj_5989), .O(n29791));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15384_4_lut.LUT_INIT = 16'hccca;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2127_3_lut (.I0(n3124), 
            .I1(n3191), .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15992_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n59971), 
            .I3(GND_net), .O(n30399));   // verilog/coms.v(130[12] 305[6])
    defparam i15992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15829_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n78), .I3(GND_net), .O(n30236));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15829_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54724 (.I0(n11999), .I1(n434), .I2(current[7]), 
            .I3(duty[23]), .O(n70939));
    defparam n11999_bdd_4_lut_54724.LUT_INIT = 16'he4aa;
    SB_LUT4 n70939_bdd_4_lut (.I0(n70939), .I1(duty[7]), .I2(n263), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n70939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i54261_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n63490), 
            .O(n2049));
    defparam i54261_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(n4_adj_5960), .I1(n5_adj_5959), .I2(n518), 
            .I3(n6_adj_5958), .O(n5_adj_6069));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'heeea;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1315_3_lut (.I0(n1928), 
            .I1(n1995), .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11999_bdd_4_lut_54719 (.I0(n11999), .I1(n435), .I2(current[6]), 
            .I3(duty[23]), .O(n70933));
    defparam n11999_bdd_4_lut_54719.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1821 (.I0(n2126), .I1(n2125), .I2(GND_net), .I3(GND_net), 
            .O(n63244));
    defparam i1_2_lut_adj_1821.LUT_INIT = 16'heeee;
    SB_LUT4 n70933_bdd_4_lut (.I0(n70933), .I1(duty[6]), .I2(n264), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n70933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30565_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n44869));
    defparam i30565_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n2122), .I1(n2128), .I2(n63244), .I3(n2127), 
            .O(n63248));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 n11999_bdd_4_lut_54714 (.I0(n11999), .I1(n436), .I2(current[5]), 
            .I3(duty[23]), .O(n70927));
    defparam n11999_bdd_4_lut_54714.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n2120), .I1(n2121), .I2(n2123), .I3(n2124), 
            .O(n63258));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 n70927_bdd_4_lut (.I0(n70927), .I1(duty[5]), .I2(n265), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n70927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(n2129), .I1(n63248), .I2(n44869), .I3(n2130), 
            .O(n63250));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'heccc;
    SB_LUT4 i43766_3_lut (.I0(n7_adj_5957), .I1(n7908), .I2(n59878), .I3(GND_net), 
            .O(n59887));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n2116), .I1(n2117), .I2(n2119), .I3(n63258), 
            .O(n63264));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 n11999_bdd_4_lut_54709 (.I0(n11999), .I1(n437), .I2(current[4]), 
            .I3(duty[23]), .O(n70921));
    defparam n11999_bdd_4_lut_54709.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_282_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i54288_4_lut (.I0(n2118), .I1(n63264), .I2(n63250), .I3(n2115), 
            .O(n2148));
    defparam i54288_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 n70921_bdd_4_lut (.I0(n70921), .I1(duty[4]), .I2(n266), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n70921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1382_3_lut (.I0(n2027), 
            .I1(n2094), .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1826 (.I0(n2224), .I1(n2223), .I2(n2227), .I3(n2225), 
            .O(n63526));
    defparam i1_4_lut_adj_1826.LUT_INIT = 16'hfffe;
    SB_LUT4 i43767_3_lut (.I0(encoder0_position_scaled_23__N_319[26]), .I1(n59887), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2226), .I1(n2221), .I2(n2222), .I3(n2228), 
            .O(n63528));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 n11999_bdd_4_lut_54704 (.I0(n11999), .I1(n438), .I2(current[3]), 
            .I3(duty[23]), .O(n70915));
    defparam n11999_bdd_4_lut_54704.LUT_INIT = 16'he4aa;
    SB_LUT4 i30499_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n44803));
    defparam i30499_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 n70915_bdd_4_lut (.I0(n70915), .I1(duty[3]), .I2(n267), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n70915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_277_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_115[20]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15980_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n59994), 
            .I3(GND_net), .O(n30387));   // verilog/coms.v(130[12] 305[6])
    defparam i15980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15830_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n78), .I3(GND_net), .O(n30237));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15830_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2126_3_lut (.I0(n3123), 
            .I1(n3190), .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n2219), .I1(n2220), .I2(n63528), .I3(n63526), 
            .O(n63534));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n2229), .I1(n44803), .I2(n2230), .I3(n2231), 
            .O(n60788));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1830 (.I0(n2217), .I1(n60788), .I2(n2218), .I3(n63534), 
            .O(n63540));
    defparam i1_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    SB_LUT4 i54031_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n63540), 
            .O(n2247));
    defparam i54031_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1449_3_lut (.I0(n2126), 
            .I1(n2193), .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15974_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n59994), 
            .I3(GND_net), .O(n30381));   // verilog/coms.v(130[12] 305[6])
    defparam i15974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1831 (.I0(n2324), .I1(n2327), .I2(GND_net), .I3(GND_net), 
            .O(n63080));
    defparam i1_2_lut_adj_1831.LUT_INIT = 16'heeee;
    SB_LUT4 i15971_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n59994), 
            .I3(GND_net), .O(n30378));   // verilog/coms.v(130[12] 305[6])
    defparam i15971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n2326), .I1(n63080), .I2(n2325), .I3(n2328), 
            .O(n63086));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i30495_3_lut (.I0(n948), .I1(n2332), .I2(n2333), .I3(GND_net), 
            .O(n44799));
    defparam i30495_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n2321), .I1(n2322), .I2(n63086), .I3(n2323), 
            .O(n63092));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i15968_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n59994), 
            .I3(GND_net), .O(n30375));   // verilog/coms.v(130[12] 305[6])
    defparam i15968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_29_lut (.I0(GND_net), 
            .I1(n3107), .I2(VCC_net), .I3(n52331), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_4 (.CI(n52251), 
            .I0(n2932), .I1(GND_net), .CO(n52252));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_12 (.CI(n52161), 
            .I0(n2524), .I1(VCC_net), .CO(n52162));
    SB_LUT4 i1_4_lut_adj_1834 (.I0(n2329), .I1(n44799), .I2(n2330), .I3(n2331), 
            .O(n60768));
    defparam i1_4_lut_adj_1834.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_4 (.CI(n52031), 
            .I0(n2032), .I1(GND_net), .CO(n52032));
    SB_LUT4 i15964_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n59994), 
            .I3(GND_net), .O(n30371));   // verilog/coms.v(130[12] 305[6])
    defparam i15964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_282_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_115[21]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15961_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n59994), 
            .I3(GND_net), .O(n30368));   // verilog/coms.v(130[12] 305[6])
    defparam i15961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15831_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[1]), .I2(n6_adj_5883), 
            .I3(n25971), .O(n30238));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15831_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2125_3_lut (.I0(n3122), 
            .I1(n3189), .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_282_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_115[22]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15958_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n59994), 
            .I3(GND_net), .O(n30365));   // verilog/coms.v(130[12] 305[6])
    defparam i15958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15954_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n28801), 
            .I3(GND_net), .O(n30361));   // verilog/coms.v(130[12] 305[6])
    defparam i15954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15832_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[2]), .I2(n6_adj_5883), 
            .I3(n25977), .O(n30239));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15832_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15945_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n28801), 
            .I3(GND_net), .O(n30352));   // verilog/coms.v(130[12] 305[6])
    defparam i15945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15941_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n28801), 
            .I3(GND_net), .O(n30348));   // verilog/coms.v(130[12] 305[6])
    defparam i15941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15833_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[3]), .I2(n6_adj_5883), 
            .I3(n25966), .O(n30240));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15833_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15935_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n28801), 
            .I3(GND_net), .O(n30342));   // verilog/coms.v(130[12] 305[6])
    defparam i15935_3_lut.LUT_INIT = 16'hacac;
    SB_DFF read_222 (.Q(state_7__N_4045[0]), .C(clk16MHz), .D(n62248));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i15931_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n28801), 
            .I3(GND_net), .O(n30338));   // verilog/coms.v(130[12] 305[6])
    defparam i15931_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n58604));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i15834_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[4]), .I2(n6_adj_5915), 
            .I3(n25959), .O(n30241));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15834_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_3_lut (.I0(GND_net), 
            .I1(n2033), .I2(VCC_net), .I3(n52030), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_3_lut (.I0(GND_net), 
            .I1(n2933), .I2(VCC_net), .I3(n52250), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_3 (.CI(n52250), 
            .I0(n2933), .I1(VCC_net), .CO(n52251));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1972_2_lut (.I0(GND_net), 
            .I1(n954), .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_20_lut (.I0(GND_net), .I1(n5413), .I2(n5438), .I3(n51637), 
            .O(n423)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23786_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n23164), .I3(GND_net), .O(n30664));
    defparam i23786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15835_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[5]), .I2(n6_adj_5915), 
            .I3(n25971), .O(n30242));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15835_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16262_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n59086), .I3(GND_net), .O(n30669));   // verilog/coms.v(130[12] 305[6])
    defparam i16262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15836_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[6]), .I2(n6_adj_5915), 
            .I3(n25977), .O(n30243));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15836_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_262_8 (.CI(n51342), .I0(duty[9]), .I1(n70691), .CO(n51343));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i973_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_264_11 (.CI(n51322), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n51323));
    SB_CARRY add_1125_20 (.CI(n51637), .I0(n5413), .I1(n5438), .CO(n51638));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1040_3_lut (.I0(n1525), 
            .I1(n1592), .I2(n1554_adj_5994), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16265_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n23230), .I3(GND_net), .O(n30672));   // verilog/coms.v(130[12] 305[6])
    defparam i16265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1835 (.I0(\data_in_frame[18] [7]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[7]), .O(n58256));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1835.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16267_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n59086), .I3(GND_net), .O(n30674));   // verilog/coms.v(130[12] 305[6])
    defparam i16267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16270_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n23164), .I3(GND_net), .O(n30677));   // verilog/coms.v(130[12] 305[6])
    defparam i16270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1836 (.I0(\data_in_frame[18] [6]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[6]), .O(n58260));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1836.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15460_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n28778), .I3(GND_net), .O(n29867));   // verilog/coms.v(130[12] 305[6])
    defparam i15460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15837_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[7]), .I2(n6_adj_5915), 
            .I3(n25966), .O(n30244));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15837_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12_4_lut_adj_1837 (.I0(\data_in_frame[18] [4]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[4]), .O(n58264));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1837.LUT_INIT = 16'h3a0a;
    SB_LUT4 add_264_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n51315), .O(encoder1_position_scaled_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2124_3_lut (.I0(n3121), 
            .I1(n3188), .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1107_3_lut (.I0(n1624), 
            .I1(n1691), .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_262_7_lut (.I0(current[5]), .I1(duty[8]), .I2(n70691), 
            .I3(n51341), .O(n265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i15838_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[8]), .I2(n6_adj_5914), 
            .I3(n25959), .O(n30245));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15838_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1174_3_lut (.I0(n1723), 
            .I1(n1790), .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15454_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n28778), .I3(GND_net), .O(n29861));   // verilog/coms.v(130[12] 305[6])
    defparam i15454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_264_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n51321), .O(encoder1_position_scaled_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1838 (.I0(\data_in_frame[18] [2]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[2]), .O(n58268));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1838.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15839_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[9]), .I2(n6_adj_5914), 
            .I3(n25971), .O(n30246));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15839_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_29 (.CI(n52331), 
            .I0(n3107), .I1(VCC_net), .CO(n52332));
    SB_LUT4 i12_4_lut_adj_1839 (.I0(\data_in_frame[18] [1]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[1]), .O(n58272));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1839.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15840_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[10]), .I2(n6_adj_5914), 
            .I3(n25977), .O(n30247));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15840_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_3 (.CI(n52030), 
            .I0(n2033), .I1(VCC_net), .CO(n52031));
    SB_LUT4 i15841_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[11]), .I2(n6_adj_5914), 
            .I3(n25966), .O(n30248));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15841_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12_4_lut_adj_1840 (.I0(\data_in_frame[18] [0]), .I1(n28719), 
            .I2(n28778), .I3(rx_data[0]), .O(n58274));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1840.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15842_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[12]), .I2(n43986), 
            .I3(n25959), .O(n30249));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15842_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12_4_lut_adj_1841 (.I0(\data_in_frame[17] [7]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[7]), .O(n58278));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1841.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1842 (.I0(\data_in_frame[17] [6]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[6]), .O(n58282));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1842.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15843_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[15]), .I2(n43986), 
            .I3(n25966), .O(n30250));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15843_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12_4_lut_adj_1843 (.I0(\data_in_frame[17] [5]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[5]), .O(n58286));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1843.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1844 (.I0(\data_in_frame[17] [4]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[4]), .O(n58290));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1844.LUT_INIT = 16'h3a0a;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_adj_1845 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n59011));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_1845.LUT_INIT = 16'h2222;
    SB_DFFESR dti_counter_2046__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n28182), 
            .D(n45), .R(n29536));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28100), 
            .D(n1561), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28100), 
            .D(n1560), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28100), 
            .D(n1559), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28100), 
            .D(n1558), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28100), 
            .D(n1557), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28100), 
            .D(n1556), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28100), 
            .D(n1555), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28100), 
            .D(n1554), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28100), 
            .D(n1553), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n28100), 
            .D(n1552), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n28100), 
            .D(n1551), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n28100), 
            .D(n1550), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n28100), 
            .D(n1549), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n28100), 
            .D(n1548), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n28100), 
            .D(n1547), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n28100), 
            .D(n1546), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n28100), 
            .D(n1545), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n28100), 
            .D(n1544), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n28100), 
            .D(n1543), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n28100), 
            .D(n1542), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n28100), 
            .D(n1541), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n28100), 
            .D(n1540), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n28100), 
            .D(n1539), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n28100), 
            .D(n1538), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n28100), 
            .D(n1537), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n28100), 
            .D(n1536), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i1_4_lut_adj_1846 (.I0(n2319), .I1(n2320), .I2(n60768), .I3(n63092), 
            .O(n63098));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1847 (.I0(\data_in_frame[17] [3]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[3]), .O(n58294));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1847.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n63098), 
            .O(n63104));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54057_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n63104), 
            .O(n2346));
    defparam i54057_4_lut.LUT_INIT = 16'h0001;
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n28100), 
            .D(n1535), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1516_3_lut (.I0(n2225), 
            .I1(n2292), .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i23_3_lut (.I0(encoder0_position_scaled_23__N_319[22]), 
            .I1(n11_adj_5953), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n936));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1241_3_lut (.I0(n1822), 
            .I1(n1889), .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1583_3_lut (.I0(n2324), 
            .I1(n2391), .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1650_3_lut (.I0(n2423), 
            .I1(n2490), .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n28100), 
            .D(n1534), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n28100), 
            .D(n1533), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i16283_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n59086), .I3(GND_net), .O(n30690));   // verilog/coms.v(130[12] 305[6])
    defparam i16283_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_262_7 (.CI(n51341), .I0(duty[8]), .I1(n70691), .CO(n51342));
    SB_LUT4 add_1125_19_lut (.I0(GND_net), .I1(n5414), .I2(n5439), .I3(n51636), 
            .O(n424)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1717_3_lut (.I0(n2522), 
            .I1(n2589), .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16286_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n23230), .I3(GND_net), .O(n30693));   // verilog/coms.v(130[12] 305[6])
    defparam i16286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1369_2_lut (.I0(GND_net), 
            .I1(n945), .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_6_lut (.I0(current[4]), .I1(duty[7]), .I2(n70691), 
            .I3(n51340), .O(n266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1369_2 (.CI(VCC_net), 
            .I0(n945), .I1(GND_net), .CO(n52030));
    SB_CARRY add_262_6 (.CI(n51340), .I0(duty[7]), .I1(n70691), .CO(n51341));
    SB_LUT4 i15845_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n62764), 
            .I3(n27_adj_5989), .O(n30252));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15845_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(control_mode[6]), .I1(control_mode[2]), 
            .I2(control_mode[4]), .I3(control_mode[5]), .O(n63892));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1850 (.I0(n63892), .I1(control_mode[7]), .I2(control_mode[3]), 
            .I3(GND_net), .O(n35592));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_3_lut_adj_1850.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1851 (.I0(control_mode[1]), .I1(n35592), .I2(control_mode[0]), 
            .I3(GND_net), .O(n61039));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_3_lut_adj_1851.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_282_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_28_lut (.I0(GND_net), 
            .I1(n3108), .I2(VCC_net), .I3(n52330), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1308_3_lut (.I0(n1921), 
            .I1(n1988), .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_277_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_115[23]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i24_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_28 (.CI(n52330), 
            .I0(n3108), .I1(VCC_net), .CO(n52331));
    SB_LUT4 add_262_5_lut (.I0(current[3]), .I1(duty[6]), .I2(n70691), 
            .I3(n51339), .O(n267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1375_3_lut (.I0(n2020), 
            .I1(n2087), .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1972_2 (.CI(VCC_net), 
            .I0(n954), .I1(GND_net), .CO(n52250));
    SB_CARRY add_262_5 (.CI(n51339), .I0(duty[6]), .I1(n70691), .CO(n51340));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1784_3_lut (.I0(n2621), 
            .I1(n2688), .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1851_3_lut (.I0(n2720), 
            .I1(n2787), .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1852_3_lut (.I0(n2721), 
            .I1(n2788), .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1919_3_lut (.I0(n2820), 
            .I1(n2887), .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1918_3_lut (.I0(n2819), 
            .I1(n2886), .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30493_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n44797));
    defparam i30493_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n2426), .I1(n2425), .I2(n2428), .I3(n2427), 
            .O(n63554));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 i15846_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n62780), 
            .I3(n27_adj_5989), .O(n30253));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15846_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n2423), .I1(n2420), .I2(n2424), .I3(n2421), 
            .O(n63556));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1854 (.I0(n2429), .I1(n44797), .I2(n2430), .I3(n2431), 
            .O(n60803));
    defparam i1_4_lut_adj_1854.LUT_INIT = 16'ha080;
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n28100), 
            .D(n1532), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i1_4_lut_adj_1855 (.I0(n60803), .I1(n2417), .I2(n63556), .I3(n63554), 
            .O(n63562));
    defparam i1_4_lut_adj_1855.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1856 (.I0(n2418), .I1(n2419), .I2(n2422), .I3(GND_net), 
            .O(n63606));
    defparam i1_3_lut_adj_1856.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n63606), .I1(n2415), .I2(n63562), .I3(n2416), 
            .O(n63566));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 i54172_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n63566), 
            .O(n2445));
    defparam i54172_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i10_3_lut (.I0(encoder0_position_scaled_23__N_319[9]), 
            .I1(n24_adj_5940), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n2525), .I1(n2526), .I2(n2524), .I3(n2528), 
            .O(n63116));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n2521), .I1(n63116), .I2(n2523), .I3(n2527), 
            .O(n63120));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'hfffe;
    SB_LUT4 i30491_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n44795));
    defparam i30491_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n28100), 
            .D(n1531), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n2529), .I1(n44795), .I2(n2530), .I3(n2531), 
            .O(n60777));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n2516), .I1(n2518), .I2(n60777), .I3(n2522), 
            .O(n63318));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n2517), .I1(n2519), .I2(n2520), .I3(n63120), 
            .O(n63126));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(n2514), .I1(n2513), .I2(n2515), .I3(n63318), 
            .O(n62091));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'hfffe;
    SB_LUT4 i54200_4_lut (.I0(n2512), .I1(n2511), .I2(n62091), .I3(n63126), 
            .O(n2544));
    defparam i54200_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i30527_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n44831));
    defparam i30527_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(n2624), .I1(n2621), .I2(n2626), .I3(n2620), 
            .O(n63598));
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1865 (.I0(\data_in_frame[17] [1]), .I1(n28725), 
            .I2(n28780), .I3(rx_data[1]), .O(n58296));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1865.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15847_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n62748), 
            .I3(n27_adj_5989), .O(n30254));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15847_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_1866 (.I0(n2627), .I1(n2623), .I2(GND_net), .I3(GND_net), 
            .O(n63498));
    defparam i1_2_lut_adj_1866.LUT_INIT = 16'heeee;
    SB_LUT4 i30555_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n44859));
    defparam i30555_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(n2617), .I1(n63498), .I2(n2619), .I3(n2625), 
            .O(n63504));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n2629), .I1(n63504), .I2(n44859), .I3(n2630), 
            .O(n63506));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'heccc;
    SB_LUT4 i16295_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n23230), .I3(GND_net), .O(n30702));   // verilog/coms.v(130[12] 305[6])
    defparam i16295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1869 (.I0(n2614), .I1(n2615), .I2(n63506), .I3(n2616), 
            .O(n63512));
    defparam i1_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1870 (.I0(n63598), .I1(n2622), .I2(n2628), .I3(GND_net), 
            .O(n63600));
    defparam i1_3_lut_adj_1870.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_14_lut (.I0(n70570), 
            .I1(n1422), .I2(VCC_net), .I3(n51826), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16296_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n23230), .I3(GND_net), .O(n30703));   // verilog/coms.v(130[12] 305[6])
    defparam i16296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_11_lut (.I0(GND_net), 
            .I1(n2525), .I2(VCC_net), .I3(n52160), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1871 (.I0(n2612), .I1(n2610), .I2(n2613), .I3(n63512), 
            .O(n62060));
    defparam i1_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 i54229_4_lut (.I0(n2618), .I1(n62060), .I2(n2611), .I3(n63600), 
            .O(n2643));
    defparam i54229_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i30647_4_lut (.I0(n829), .I1(n828), .I2(n44831), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i30647_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1728_3_lut (.I0(n2533), 
            .I1(n2600), .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1872 (.I0(n2726), .I1(n2724), .I2(GND_net), .I3(GND_net), 
            .O(n63298));
    defparam i1_2_lut_adj_1872.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1873 (.I0(n2725), .I1(n63298), .I2(n2722), .I3(n2728), 
            .O(n63302));
    defparam i1_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_LUT4 i43758_3_lut (.I0(n3_adj_5961), .I1(n7904), .I2(n59878), .I3(GND_net), 
            .O(n59879));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43759_3_lut (.I0(encoder0_position_scaled_23__N_319[30]), .I1(n59879), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam i43759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30553_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n44857));
    defparam i30553_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15848_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n62828), 
            .I3(n27_adj_5989), .O(n30255));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15848_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1442_3_lut (.I0(n2119), 
            .I1(n2186), .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1874 (.I0(n42166), .I1(n8_adj_5843), .I2(GND_net), 
            .I3(GND_net), .O(n28780));
    defparam i1_2_lut_adj_1874.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1875 (.I0(n2717), .I1(n2718), .I2(n2720), .I3(n63302), 
            .O(n63308));
    defparam i1_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_LUT4 i15849_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n62812), 
            .I3(n27_adj_5989), .O(n30256));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15849_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1876 (.I0(n2716), .I1(n2729), .I2(n44857), .I3(n2730), 
            .O(n63462));
    defparam i1_4_lut_adj_1876.LUT_INIT = 16'heaaa;
    SB_LUT4 i16298_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n23230), .I3(GND_net), .O(n30705));   // verilog/coms.v(130[12] 305[6])
    defparam i16298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16299_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n23164), .I3(GND_net), .O(n30706));   // verilog/coms.v(130[12] 305[6])
    defparam i16299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16300_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n23230), .I3(GND_net), .O(n30707));   // verilog/coms.v(130[12] 305[6])
    defparam i16300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [3]), 
            .O(n58959));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i16303_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n23230), .I3(GND_net), .O(n30710));   // verilog/coms.v(130[12] 305[6])
    defparam i16303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [4]), 
            .O(n58958));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [5]), 
            .O(n58957));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [6]), 
            .O(n58825));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [7]), 
            .O(n58956));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [0]), 
            .O(n58955));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2123_3_lut (.I0(n3120), 
            .I1(n3187), .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_27_lut (.I0(GND_net), 
            .I1(n3109), .I2(VCC_net), .I3(n52329), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n57536));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_11 (.CI(n52160), 
            .I0(n2525), .I1(VCC_net), .CO(n52161));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i28_3_lut (.I0(encoder0_position_scaled_23__N_319[27]), 
            .I1(n6_adj_5958), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_28_lut (.I0(GND_net), 
            .I1(n2808), .I2(VCC_net), .I3(n52249), .O(n2875)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_13_lut (.I0(GND_net), 
            .I1(n1423), .I2(VCC_net), .I3(n51825), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15850_3_lut (.I0(\data_in_frame[2] [6]), .I1(rx_data[6]), .I2(n59079), 
            .I3(GND_net), .O(n30257));   // verilog/coms.v(130[12] 305[6])
    defparam i15850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [1]), 
            .O(n58954));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_13 (.CI(n51825), 
            .I0(n1423), .I1(VCC_net), .CO(n51826));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [2]), 
            .O(n58953));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i29_3_lut (.I0(encoder0_position_scaled_23__N_319[28]), 
            .I1(n5_adj_5959), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [3]), 
            .O(n58952));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_27_lut (.I0(GND_net), 
            .I1(n2809), .I2(VCC_net), .I3(n52248), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_27 (.CI(n52248), 
            .I0(n2809), .I1(VCC_net), .CO(n52249));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1509_3_lut (.I0(n2218), 
            .I1(n2285), .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_26_lut (.I0(GND_net), 
            .I1(n2810), .I2(VCC_net), .I3(n52247), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_27 (.CI(n52329), 
            .I0(n3109), .I1(VCC_net), .CO(n52330));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1576_3_lut (.I0(n2317), 
            .I1(n2384), .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n58640));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_26_lut (.I0(GND_net), 
            .I1(n3110), .I2(VCC_net), .I3(n52328), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [4]), 
            .O(n58951));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [5]), 
            .O(n58950));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [6]), 
            .O(n58949));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[9] [7]), 
            .O(n58948));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [0]), 
            .O(n58947));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [5]), 
            .O(n58972));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_10_lut (.I0(GND_net), 
            .I1(n2526), .I2(VCC_net), .I3(n52159), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_12_lut (.I0(GND_net), 
            .I1(n1424), .I2(VCC_net), .I3(n51824), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n43842), .O(n57618));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [1]), 
            .O(n58946));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [6]), 
            .O(n58971));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n2719), .I1(n2723), .I2(n2721), .I3(n2727), 
            .O(n63232));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [2]), 
            .O(n58945));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_12 (.CI(n51824), 
            .I0(n1424), .I1(VCC_net), .CO(n51825));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [3]), 
            .O(n58944));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_LUT4 i15628_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [6]), .I1(rx_data[6]), 
            .I2(reset), .I3(n51), .O(n30035));   // verilog/coms.v(130[12] 305[6])
    defparam i15628_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [4]), 
            .O(n58943));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 i15624_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n51), .O(n30031));   // verilog/coms.v(130[12] 305[6])
    defparam i15624_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15621_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(reset), .I3(n51), .O(n30028));   // verilog/coms.v(130[12] 305[6])
    defparam i15621_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15609_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [3]), .I1(rx_data[3]), 
            .I2(reset), .I3(n51), .O(n30016));   // verilog/coms.v(130[12] 305[6])
    defparam i15609_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_26 (.CI(n52328), 
            .I0(n3110), .I1(VCC_net), .CO(n52329));
    SB_LUT4 i15573_3_lut_4_lut_4_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(reset), .I3(n51), .O(n29980));   // verilog/coms.v(130[12] 305[6])
    defparam i15573_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [5]), 
            .O(n58942));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [6]), 
            .O(n58941));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[10] [7]), 
            .O(n58940));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i16335_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n23164), .I3(GND_net), .O(n30742));   // verilog/coms.v(130[12] 305[6])
    defparam i16335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [0]), 
            .O(n58939));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [1]), 
            .O(n58938));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i16337_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n23230), .I3(GND_net), .O(n30744));   // verilog/coms.v(130[12] 305[6])
    defparam i16337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(n15_adj_5909), .I1(n23298), .I2(dti), 
            .I3(GND_net), .O(n28033));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [2]), 
            .O(n58937));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [3]), 
            .O(n58936));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [4]), 
            .O(n58935));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i30463_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n44767));
    defparam i30463_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [5]), 
            .O(n58934));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 i16342_3_lut (.I0(current[11]), .I1(data_adj_6147[11]), .I2(n28109), 
            .I3(GND_net), .O(n30749));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16342_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_10 (.CI(n52159), 
            .I0(n2526), .I1(VCC_net), .CO(n52160));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_26 (.CI(n52247), 
            .I0(n2810), .I1(VCC_net), .CO(n52248));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_25_lut (.I0(GND_net), 
            .I1(n2811), .I2(VCC_net), .I3(n52246), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16343_3_lut (.I0(current[10]), .I1(data_adj_6147[10]), .I2(n28109), 
            .I3(GND_net), .O(n30750));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29440_3_lut (.I0(current[9]), .I1(data_adj_6147[9]), .I2(n28109), 
            .I3(GND_net), .O(n30751));
    defparam i29440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [6]), 
            .O(n58933));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[11] [7]), 
            .O(n58932));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i16345_3_lut (.I0(current[8]), .I1(data_adj_6147[8]), .I2(n28109), 
            .I3(GND_net), .O(n30752));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16346_3_lut (.I0(current[7]), .I1(data_adj_6147[7]), .I2(n28109), 
            .I3(GND_net), .O(n30753));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [0]), 
            .O(n58931));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [1]), 
            .O(n58930));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [2]), 
            .O(n58929));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i16347_3_lut (.I0(current[6]), .I1(data_adj_6147[6]), .I2(n28109), 
            .I3(GND_net), .O(n30754));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16348_3_lut (.I0(current[5]), .I1(data_adj_6147[5]), .I2(n28109), 
            .I3(GND_net), .O(n30755));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16349_3_lut (.I0(current[4]), .I1(data_adj_6147[4]), .I2(n28109), 
            .I3(GND_net), .O(n30756));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16350_3_lut (.I0(current[3]), .I1(data_adj_6147[3]), .I2(n28109), 
            .I3(GND_net), .O(n30757));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [3]), 
            .O(n58928));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 i29322_3_lut (.I0(current[2]), .I1(data_adj_6147[2]), .I2(n28109), 
            .I3(GND_net), .O(n30758));
    defparam i29322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16352_3_lut (.I0(current[1]), .I1(data_adj_6147[1]), .I2(n28109), 
            .I3(GND_net), .O(n30759));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16353_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n23230), .I3(GND_net), .O(n30760));   // verilog/coms.v(130[12] 305[6])
    defparam i16353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16354_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n23230), .I3(GND_net), .O(n30761));   // verilog/coms.v(130[12] 305[6])
    defparam i16354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [4]), 
            .O(n58927));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 i16356_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n23230), .I3(GND_net), .O(n30763));   // verilog/coms.v(130[12] 305[6])
    defparam i16356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [5]), 
            .O(n58926));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 i16358_3_lut (.I0(baudrate[31]), .I1(data_adj_6138[7]), .I2(n62253), 
            .I3(GND_net), .O(n30765));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16358_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16359_3_lut (.I0(baudrate[30]), .I1(data_adj_6138[6]), .I2(n62253), 
            .I3(GND_net), .O(n30766));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16359_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16360_3_lut (.I0(baudrate[29]), .I1(data_adj_6138[5]), .I2(n62253), 
            .I3(GND_net), .O(n30767));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16360_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i30_3_lut (.I0(encoder0_position_scaled_23__N_319[29]), 
            .I1(n4_adj_5960), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16361_3_lut (.I0(baudrate[28]), .I1(data_adj_6138[4]), .I2(n62253), 
            .I3(GND_net), .O(n30768));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1184_3_lut (.I0(n1733), 
            .I1(n1800), .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1251_3_lut (.I0(n1832), 
            .I1(n1899), .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16362_3_lut (.I0(baudrate[27]), .I1(data_adj_6138[3]), .I2(n62253), 
            .I3(GND_net), .O(n30769));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1318_3_lut (.I0(n1931), 
            .I1(n1998), .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1385_3_lut (.I0(n2030), 
            .I1(n2097), .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1643_3_lut (.I0(n2416), 
            .I1(n2483), .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1710_3_lut (.I0(n2515), 
            .I1(n2582), .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [6]), 
            .O(n58925));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 i16363_3_lut (.I0(baudrate[26]), .I1(data_adj_6138[2]), .I2(n62253), 
            .I3(GND_net), .O(n30770));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15853_3_lut (.I0(\data_in_frame[2] [7]), .I1(rx_data[7]), .I2(n59079), 
            .I3(GND_net), .O(n30260));   // verilog/coms.v(130[12] 305[6])
    defparam i15853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16364_3_lut (.I0(baudrate[25]), .I1(data_adj_6138[1]), .I2(n62253), 
            .I3(GND_net), .O(n30771));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16364_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1777_3_lut (.I0(n2614), 
            .I1(n2681), .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[12] [7]), 
            .O(n58924));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i16365_3_lut (.I0(baudrate[24]), .I1(data_adj_6138[0]), .I2(n62253), 
            .I3(GND_net), .O(n30772));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16366_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n23230), .I3(GND_net), .O(n30773));   // verilog/coms.v(130[12] 305[6])
    defparam i16366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16728_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3358));   // verilog/coms.v(130[12] 305[6])
    defparam i16728_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2122_3_lut (.I0(n3119), 
            .I1(n3186), .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [0]), 
            .O(n58826));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1844_3_lut (.I0(n2713), 
            .I1(n2780), .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_25_lut (.I0(GND_net), 
            .I1(n3111), .I2(VCC_net), .I3(n52327), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i31_3_lut (.I0(encoder0_position_scaled_23__N_319[30]), 
            .I1(n3_adj_5961), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6605_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_468));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6605_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2121_3_lut (.I0(n3118), 
            .I1(n3185), .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1917 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [1]), 
            .O(n58923));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1917.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2120_3_lut (.I0(n3117), 
            .I1(n3184), .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6607_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_485));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6607_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1845_3_lut (.I0(n2714), 
            .I1(n2781), .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [2]), 
            .O(n58922));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [3]), 
            .O(n58921));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 i6609_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_490));
    defparam i6609_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [4]), 
            .O(n58920));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2119_3_lut (.I0(n3116), 
            .I1(n3183), .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2118_3_lut (.I0(n3115), 
            .I1(n3182), .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2117_3_lut (.I0(n3114), 
            .I1(n3181), .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2116_3_lut (.I0(n3113), 
            .I1(n3180), .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_25 (.CI(n52246), 
            .I0(n2811), .I1(VCC_net), .CO(n52247));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2115_3_lut (.I0(n3112), 
            .I1(n3179), .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [5]), 
            .O(n58919));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h2300;
    SB_LUT4 i6611_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_499));
    defparam i6611_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [6]), 
            .O(n58918));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[13] [7]), 
            .O(n58917));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [0]), 
            .O(n58916));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [1]), 
            .O(n58915));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [2]), 
            .O(n58914));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [3]), 
            .O(n58913));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [4]), 
            .O(n58912));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h2300;
    SB_LUT4 i53793_2_lut (.I0(state_7__N_4253[3]), .I1(n11_adj_5912), .I2(GND_net), 
            .I3(GND_net), .O(n62));
    defparam i53793_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [5]), 
            .O(n58911));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [6]), 
            .O(n58910));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1931 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[14] [7]), 
            .O(n58909));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1931.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [0]), 
            .O(n58908));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_LUT4 add_6183_32_lut (.I0(GND_net), .I1(encoder0_position[31]), .I2(VCC_net), 
            .I3(n53140), .O(encoder0_position_scaled_23__N_319[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6183_31_lut (.I0(GND_net), .I1(encoder0_position[30]), .I2(VCC_net), 
            .I3(n53139), .O(encoder0_position_scaled_23__N_319[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_31 (.CI(n53139), .I0(encoder0_position[30]), .I1(VCC_net), 
            .CO(n53140));
    SB_LUT4 add_6183_30_lut (.I0(GND_net), .I1(encoder0_position[29]), .I2(VCC_net), 
            .I3(n53138), .O(encoder0_position_scaled_23__N_319[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_30 (.CI(n53138), .I0(encoder0_position[29]), .I1(VCC_net), 
            .CO(n53139));
    SB_LUT4 add_6183_29_lut (.I0(GND_net), .I1(encoder0_position[28]), .I2(VCC_net), 
            .I3(n53137), .O(encoder0_position_scaled_23__N_319[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_29 (.CI(n53137), .I0(encoder0_position[28]), .I1(VCC_net), 
            .CO(n53138));
    SB_LUT4 add_6183_28_lut (.I0(GND_net), .I1(encoder0_position[27]), .I2(VCC_net), 
            .I3(n53136), .O(encoder0_position_scaled_23__N_319[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_28 (.CI(n53136), .I0(encoder0_position[27]), .I1(VCC_net), 
            .CO(n53137));
    SB_LUT4 add_6183_27_lut (.I0(GND_net), .I1(encoder0_position[26]), .I2(VCC_net), 
            .I3(n53135), .O(encoder0_position_scaled_23__N_319[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_27 (.CI(n53135), .I0(encoder0_position[26]), .I1(VCC_net), 
            .CO(n53136));
    SB_LUT4 add_6183_26_lut (.I0(GND_net), .I1(encoder0_position[25]), .I2(VCC_net), 
            .I3(n53134), .O(encoder0_position_scaled_23__N_319[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_26 (.CI(n53134), .I0(encoder0_position[25]), .I1(VCC_net), 
            .CO(n53135));
    SB_LUT4 add_6183_25_lut (.I0(GND_net), .I1(encoder0_position[24]), .I2(VCC_net), 
            .I3(n53133), .O(encoder0_position_scaled_23__N_319[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_25 (.CI(n53133), .I0(encoder0_position[24]), .I1(VCC_net), 
            .CO(n53134));
    SB_LUT4 add_6183_24_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(VCC_net), 
            .I3(n53132), .O(encoder0_position_scaled_23__N_319[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_24 (.CI(n53132), .I0(encoder0_position[23]), .I1(VCC_net), 
            .CO(n53133));
    SB_LUT4 add_6183_23_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(VCC_net), 
            .I3(n53131), .O(encoder0_position_scaled_23__N_319[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_23 (.CI(n53131), .I0(encoder0_position[22]), .I1(VCC_net), 
            .CO(n53132));
    SB_LUT4 add_6183_22_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(VCC_net), 
            .I3(n53130), .O(encoder0_position_scaled_23__N_319[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_22 (.CI(n53130), .I0(encoder0_position[21]), .I1(VCC_net), 
            .CO(n53131));
    SB_LUT4 add_6183_21_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(VCC_net), 
            .I3(n53129), .O(encoder0_position_scaled_23__N_319[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_21 (.CI(n53129), .I0(encoder0_position[20]), .I1(VCC_net), 
            .CO(n53130));
    SB_LUT4 add_6183_20_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(VCC_net), 
            .I3(n53128), .O(encoder0_position_scaled_23__N_319[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_20 (.CI(n53128), .I0(encoder0_position[19]), .I1(VCC_net), 
            .CO(n53129));
    SB_LUT4 add_6183_19_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(VCC_net), 
            .I3(n53127), .O(encoder0_position_scaled_23__N_319[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_19 (.CI(n53127), .I0(encoder0_position[18]), .I1(VCC_net), 
            .CO(n53128));
    SB_LUT4 add_6183_18_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(VCC_net), 
            .I3(n53126), .O(encoder0_position_scaled_23__N_319[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_18 (.CI(n53126), .I0(encoder0_position[17]), .I1(VCC_net), 
            .CO(n53127));
    SB_LUT4 add_6183_17_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(VCC_net), 
            .I3(n53125), .O(encoder0_position_scaled_23__N_319[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_17 (.CI(n53125), .I0(encoder0_position[16]), .I1(VCC_net), 
            .CO(n53126));
    SB_LUT4 add_6183_16_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(VCC_net), 
            .I3(n53124), .O(encoder0_position_scaled_23__N_319[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_16 (.CI(n53124), .I0(encoder0_position[15]), .I1(VCC_net), 
            .CO(n53125));
    SB_LUT4 add_6183_15_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(VCC_net), 
            .I3(n53123), .O(encoder0_position_scaled_23__N_319[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_15 (.CI(n53123), .I0(encoder0_position[14]), .I1(VCC_net), 
            .CO(n53124));
    SB_LUT4 add_6183_14_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(VCC_net), 
            .I3(n53122), .O(encoder0_position_scaled_23__N_319[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_14 (.CI(n53122), .I0(encoder0_position[13]), .I1(VCC_net), 
            .CO(n53123));
    SB_LUT4 add_6183_13_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(VCC_net), 
            .I3(n53121), .O(encoder0_position_scaled_23__N_319[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_13 (.CI(n53121), .I0(encoder0_position[12]), .I1(VCC_net), 
            .CO(n53122));
    SB_LUT4 add_6183_12_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(VCC_net), 
            .I3(n53120), .O(encoder0_position_scaled_23__N_319[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_12 (.CI(n53120), .I0(encoder0_position[11]), .I1(VCC_net), 
            .CO(n53121));
    SB_LUT4 add_6183_11_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(VCC_net), 
            .I3(n53119), .O(encoder0_position_scaled_23__N_319[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_11 (.CI(n53119), .I0(encoder0_position[10]), .I1(VCC_net), 
            .CO(n53120));
    SB_LUT4 add_6183_10_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(VCC_net), 
            .I3(n53118), .O(encoder0_position_scaled_23__N_319[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_10 (.CI(n53118), .I0(encoder0_position[9]), .I1(VCC_net), 
            .CO(n53119));
    SB_LUT4 add_6183_9_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(VCC_net), 
            .I3(n53117), .O(encoder0_position_scaled_23__N_319[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_9 (.CI(n53117), .I0(encoder0_position[8]), .I1(VCC_net), 
            .CO(n53118));
    SB_LUT4 add_6183_8_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(VCC_net), 
            .I3(n53116), .O(encoder0_position_scaled_23__N_319[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_8 (.CI(n53116), .I0(encoder0_position[7]), .I1(VCC_net), 
            .CO(n53117));
    SB_LUT4 add_6183_7_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(VCC_net), 
            .I3(n53115), .O(encoder0_position_scaled_23__N_319[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_7 (.CI(n53115), .I0(encoder0_position[6]), .I1(VCC_net), 
            .CO(n53116));
    SB_LUT4 add_6183_6_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(VCC_net), 
            .I3(n53114), .O(encoder0_position_scaled_23__N_319[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_6 (.CI(n53114), .I0(encoder0_position[5]), .I1(VCC_net), 
            .CO(n53115));
    SB_LUT4 add_6183_5_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(VCC_net), 
            .I3(n53113), .O(encoder0_position_scaled_23__N_319[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_5 (.CI(n53113), .I0(encoder0_position[4]), .I1(VCC_net), 
            .CO(n53114));
    SB_LUT4 add_6183_4_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(VCC_net), 
            .I3(n53112), .O(encoder0_position_scaled_23__N_319[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_4 (.CI(n53112), .I0(encoder0_position[3]), .I1(VCC_net), 
            .CO(n53113));
    SB_LUT4 add_6183_3_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(VCC_net), 
            .I3(n53111), .O(encoder0_position_scaled_23__N_319[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_3 (.CI(n53111), .I0(encoder0_position[2]), .I1(VCC_net), 
            .CO(n53112));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [1]), 
            .O(n58907));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 add_6183_2_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(VCC_net), 
            .I3(n53110), .O(encoder0_position_scaled_23__N_319[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_2 (.CI(n53110), .I0(encoder0_position[1]), .I1(VCC_net), 
            .CO(n53111));
    SB_CARRY add_6183_1 (.CI(GND_net), .I0(encoder0_position[0]), .I1(encoder0_position[0]), 
            .CO(n53110));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [2]), 
            .O(n58906));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [3]), 
            .O(n58905));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [4]), 
            .O(n58904));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [5]), 
            .O(n58903));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1912_3_lut (.I0(n2813), 
            .I1(n2880), .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i18_3_lut (.I0(encoder0_position_scaled_23__N_319[17]), 
            .I1(n16_adj_5948), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1911_3_lut (.I0(n2812), 
            .I1(n2879), .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30203_2_lut_2_lut (.I0(duty[23]), .I1(n296), .I2(GND_net), 
            .I3(GND_net), .O(n5433));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30203_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [6]), 
            .O(n58902));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 i16383_3_lut (.I0(baudrate[7]), .I1(data_adj_6138[7]), .I2(n61238), 
            .I3(GND_net), .O(n30790));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16384_3_lut (.I0(baudrate[6]), .I1(data_adj_6138[6]), .I2(n61238), 
            .I3(GND_net), .O(n30791));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[15] [7]), 
            .O(n58901));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [0]), 
            .O(n58900));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i16385_3_lut (.I0(baudrate[5]), .I1(data_adj_6138[5]), .I2(n61238), 
            .I3(GND_net), .O(n30792));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1941 (.I0(n2713), .I1(n63462), .I2(n63308), .I3(n2715), 
            .O(n63312));
    defparam i1_4_lut_adj_1941.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1942 (.I0(n2710), .I1(n2712), .I2(n2714), .I3(n63232), 
            .O(n63238));
    defparam i1_4_lut_adj_1942.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [1]), 
            .O(n58899));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1910_3_lut (.I0(n2811), 
            .I1(n2878), .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16386_3_lut (.I0(baudrate[4]), .I1(data_adj_6138[4]), .I2(n61238), 
            .I3(GND_net), .O(n30793));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6115_2_lut (.I0(n2_adj_5962), .I1(encoder0_position_scaled_23__N_319[31]), 
            .I2(GND_net), .I3(GND_net), .O(n621));
    defparam i6115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [2]), 
            .O(n58829));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i500_4_lut (.I0(n621), .I1(n7903), 
            .I2(n63466), .I3(n5_adj_6069), .O(n828));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i500_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5900));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5901));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5897));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5898));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i24_3_lut (.I0(encoder0_position_scaled_23__N_319[23]), 
            .I1(n10_adj_5954), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n935));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16387_3_lut (.I0(baudrate[3]), .I1(data_adj_6138[3]), .I2(n61238), 
            .I3(GND_net), .O(n30794));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16388_3_lut (.I0(baudrate[2]), .I1(data_adj_6138[2]), .I2(n61238), 
            .I3(GND_net), .O(n30795));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i5_2_lut (.I0(current[2]), .I1(duty[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5906));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i9_3_lut (.I0(encoder0_position_scaled_23__N_319[8]), 
            .I1(n25_adj_5939), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5904));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5903));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51580_4_lut (.I0(n9_adj_5903), .I1(n7_adj_5904), .I2(n5_adj_5906), 
            .I3(current[0]), .O(n67754));
    defparam i51580_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1796_3_lut (.I0(n2633), 
            .I1(n2700), .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i709_3_lut (.I0(n935), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_11_lut (.I0(GND_net), 
            .I1(n1425), .I2(VCC_net), .I3(n51823), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_11 (.CI(n51823), 
            .I0(n1425), .I1(VCC_net), .CO(n51824));
    SB_LUT4 i16389_3_lut (.I0(baudrate[1]), .I1(data_adj_6138[1]), .I2(n61238), 
            .I3(GND_net), .O(n30796));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [3]), 
            .O(n58832));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i14_3_lut (.I0(n6_adj_5905), .I1(duty[8]), .I2(n17_adj_5897), 
            .I3(GND_net), .O(n14_adj_5899));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_25 (.CI(n52327), 
            .I0(n3111), .I1(VCC_net), .CO(n52328));
    SB_LUT4 i20574_3_lut (.I0(duty[1]), .I1(current[1]), .I2(duty[0]), 
            .I3(GND_net), .O(n34970));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i20574_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i53171_3_lut (.I0(n34970), .I1(duty[4]), .I2(n9_adj_5903), 
            .I3(GND_net), .O(n69346));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53172_3_lut (.I0(n69346), .I1(duty[5]), .I2(n11_adj_5901), 
            .I3(GND_net), .O(n69347));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51572_4_lut (.I0(n15_adj_5898), .I1(n13_adj_5900), .I2(n11_adj_5901), 
            .I3(n67754), .O(n67746));
    defparam i51572_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53462_4_lut (.I0(n14_adj_5899), .I1(n4_adj_5907), .I2(n17_adj_5897), 
            .I3(n67742), .O(n69637));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53462_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51956_3_lut (.I0(n69347), .I1(duty[6]), .I2(n13_adj_5900), 
            .I3(GND_net), .O(n68130));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53672_4_lut (.I0(n68130), .I1(n69637), .I2(n17_adj_5897), 
            .I3(n67746), .O(n69847));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53672_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_9_lut (.I0(GND_net), 
            .I1(n2527), .I2(VCC_net), .I3(n52158), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11999_bdd_4_lut_54699 (.I0(n11999), .I1(n439), .I2(current[2]), 
            .I3(duty[23]), .O(n70897));
    defparam n11999_bdd_4_lut_54699.LUT_INIT = 16'he4aa;
    SB_LUT4 n70897_bdd_4_lut (.I0(n70897), .I1(duty[2]), .I2(n268), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n70897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1946 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n63278));
    defparam i1_2_lut_adj_1946.LUT_INIT = 16'h8888;
    SB_LUT4 n11999_bdd_4_lut_54684 (.I0(n11999), .I1(n440), .I2(current[1]), 
            .I3(duty[23]), .O(n70891));
    defparam n11999_bdd_4_lut_54684.LUT_INIT = 16'he4aa;
    SB_LUT4 n70891_bdd_4_lut (.I0(n70891), .I1(duty[1]), .I2(n269), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n70891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1947 (.I0(n927), .I1(n63278), .I2(n928), .I3(n44767), 
            .O(n960));
    defparam i1_4_lut_adj_1947.LUT_INIT = 16'hfefa;
    SB_LUT4 n11999_bdd_4_lut_54679 (.I0(n11999), .I1(n441), .I2(current[0]), 
            .I3(duty[23]), .O(n70885));
    defparam n11999_bdd_4_lut_54679.LUT_INIT = 16'he4aa;
    SB_LUT4 n70885_bdd_4_lut (.I0(n70885), .I1(duty[0]), .I2(n270), .I3(duty[23]), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n70885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30461_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n44765));
    defparam i30461_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1948 (.I0(n1029), .I1(n44765), .I2(n1030), .I3(n1031), 
            .O(n60705));
    defparam i1_4_lut_adj_1948.LUT_INIT = 16'ha080;
    SB_LUT4 i16390_3_lut (.I0(baudrate[0]), .I1(data_adj_6138[0]), .I2(n61238), 
            .I3(GND_net), .O(n30797));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16390_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54470_4_lut (.I0(n1026), .I1(n60705), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i54470_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54661 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n70861));
    defparam byte_transmit_counter_0__bdd_4_lut_54661.LUT_INIT = 16'he4aa;
    SB_LUT4 n70861_bdd_4_lut (.I0(n70861), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n70864));
    defparam n70861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [4]), 
            .O(n58833));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 i16391_3_lut (.I0(ID[7]), .I1(data_adj_6138[7]), .I2(n59065), 
            .I3(GND_net), .O(n30798));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [5]), 
            .O(n58834));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [6]), 
            .O(n58835));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2111_3_lut (.I0(n3108), 
            .I1(n3175), .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53673_3_lut (.I0(n69847), .I1(duty[9]), .I2(current[9]), 
            .I3(GND_net), .O(n69848));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53673_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54087_4_lut (.I0(n63238), .I1(n2709), .I2(n63312), .I3(n2711), 
            .O(n2742));
    defparam i54087_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53580_3_lut (.I0(n69848), .I1(duty[10]), .I2(current[10]), 
            .I3(GND_net), .O(n69755));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53580_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16392_3_lut (.I0(ID[6]), .I1(data_adj_6138[6]), .I2(n59065), 
            .I3(GND_net), .O(n30799));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n69755), .I1(duty[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5896));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_24_lut (.I0(GND_net), 
            .I1(n3112), .I2(VCC_net), .I3(n52326), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16393_3_lut (.I0(ID[5]), .I1(data_adj_6138[5]), .I2(n59065), 
            .I3(GND_net), .O(n30800));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i977_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_9 (.CI(n52158), 
            .I0(n2527), .I1(VCC_net), .CO(n52159));
    SB_LUT4 i16394_3_lut (.I0(ID[4]), .I1(data_adj_6138[4]), .I2(n59065), 
            .I3(GND_net), .O(n30801));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16394_3_lut.LUT_INIT = 16'hacac;
    SB_DFF reset_223 (.Q(reset), .C(clk16MHz), .D(n57618));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[16] [7]), 
            .O(n58836));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i16395_3_lut (.I0(ID[3]), .I1(data_adj_6138[3]), .I2(n59065), 
            .I3(GND_net), .O(n30802));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut (.I0(duty[14]), .I1(n24_adj_5896), .I2(duty[12]), 
            .I3(duty[13]), .O(n61279));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [0]), 
            .O(n58841));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_1954 (.I0(duty[14]), .I1(n24_adj_5896), .I2(duty[12]), 
            .I3(duty[13]), .O(n61284));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1954.LUT_INIT = 16'h8000;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_24 (.CI(n52326), 
            .I0(n3112), .I1(VCC_net), .CO(n52327));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1044_3_lut (.I0(n1529), 
            .I1(n1596), .I2(n1554_adj_5994), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1955 (.I0(duty[15]), .I1(current[15]), .I2(n61284), 
            .I3(n61279), .O(n32));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1955.LUT_INIT = 16'hb3a2;
    SB_CARRY add_1125_19 (.CI(n51636), .I0(n5414), .I1(n5439), .CO(n51637));
    SB_LUT4 i16396_3_lut (.I0(ID[2]), .I1(data_adj_6138[2]), .I2(n59065), 
            .I3(GND_net), .O(n30803));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16397_3_lut (.I0(ID[1]), .I1(data_adj_6138[1]), .I2(n59065), 
            .I3(GND_net), .O(n30804));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1956 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n61347));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1956.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1957 (.I0(duty[18]), .I1(n32), .I2(duty[16]), 
            .I3(duty[17]), .O(n61350));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1957.LUT_INIT = 16'h8000;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1111_3_lut (.I0(n1628), 
            .I1(n1695), .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1958 (.I0(duty[19]), .I1(current[15]), .I2(n61350), 
            .I3(n61347), .O(n40));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_adj_1958.LUT_INIT = 16'hb3a2;
    SB_LUT4 add_262_4_lut (.I0(current[2]), .I1(duty[5]), .I2(n70691), 
            .I3(n51338), .O(n268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_10_lut (.I0(GND_net), 
            .I1(n1426), .I2(VCC_net), .I3(n51822), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_10 (.CI(n51822), 
            .I0(n1426), .I1(VCC_net), .CO(n51823));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_24_lut (.I0(GND_net), 
            .I1(n2812), .I2(VCC_net), .I3(n52245), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_23_lut (.I0(GND_net), 
            .I1(n3113), .I2(VCC_net), .I3(n52325), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1959 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n61440));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1959.LUT_INIT = 16'hfffe;
    SB_LUT4 add_1125_18_lut (.I0(GND_net), .I1(n5415), .I2(n5440), .I3(n51635), 
            .O(n425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1960 (.I0(duty[22]), .I1(n40), .I2(duty[20]), 
            .I3(duty[21]), .O(n61445));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i3_4_lut_adj_1960.LUT_INIT = 16'h8000;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_9_lut (.I0(GND_net), 
            .I1(n1427), .I2(VCC_net), .I3(n51821), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16398_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3844 [23]), 
            .I2(control_update), .I3(GND_net), .O(n30805));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_8_lut (.I0(GND_net), 
            .I1(n2528), .I2(VCC_net), .I3(n52157), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_9 (.CI(n51821), 
            .I0(n1427), .I1(VCC_net), .CO(n51822));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [1]), 
            .O(n58843));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [2]), 
            .O(n58847));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i16399_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3844 [22]), 
            .I2(control_update), .I3(GND_net), .O(n30806));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [3]), 
            .O(n58848));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1178_3_lut (.I0(n1727), 
            .I1(n1794), .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16400_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3844 [21]), 
            .I2(control_update), .I3(GND_net), .O(n30807));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16401_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3844 [20]), 
            .I2(control_update), .I3(GND_net), .O(n30808));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5846));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_24 (.CI(n52245), 
            .I0(n2812), .I1(VCC_net), .CO(n52246));
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28100), 
            .D(n1562), .R(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_8_lut (.I0(GND_net), 
            .I1(n1428), .I2(VCC_net), .I3(n51820), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_18 (.CI(n51635), .I0(n5415), .I1(n5440), .CO(n51636));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_8 (.CI(n51820), 
            .I0(n1428), .I1(VCC_net), .CO(n51821));
    SB_LUT4 add_1125_17_lut (.I0(GND_net), .I1(n5416), .I2(n5441), .I3(n51634), 
            .O(n426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_23 (.CI(n52325), 
            .I0(n3113), .I1(VCC_net), .CO(n52326));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_7_lut (.I0(GND_net), 
            .I1(n1429), .I2(GND_net), .I3(n51819), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_7 (.CI(n51819), 
            .I0(n1429), .I1(GND_net), .CO(n51820));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_6_lut (.I0(GND_net), 
            .I1(n1430), .I2(GND_net), .I3(n51818), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_6 (.CI(n51818), 
            .I0(n1430), .I1(GND_net), .CO(n51819));
    SB_LUT4 LessThan_17_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5844));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_91[23]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_91[22]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 LessThan_17_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_91[21]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_91[20]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_91[19]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_91[18]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_91[17]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_91[16]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_91[15]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_91[14]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_91[13]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_91[12]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_91[11]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_91[10]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_91[9]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_91[8]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_91[7]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_91[6]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_91[5]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_91[4]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_91[3]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_91[2]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_91[1]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 i16402_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(\PID_CONTROLLER.integral_23__N_3844 [19]), 
            .I2(control_update), .I3(GND_net), .O(n30809));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16402_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR GHC_215 (.Q(GHC), .C(clk16MHz), .E(n28059), .D(GHC_N_504), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_213 (.Q(GHB), .C(clk16MHz), .E(n28059), .D(GHB_N_490), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_211 (.Q(GHA), .C(clk16MHz), .E(n28059), .D(GHA_N_468), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_6090), .D(commutation_state_7__N_256[0]), .S(commutation_state_7__N_264));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_212 (.Q(INLA_c_0), .C(clk16MHz), .E(n28059), .D(GLA_N_485), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[23]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[22]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 i51615_4_lut (.I0(n11), .I1(n9_adj_5844), .I2(n7_adj_5846), 
            .I3(n5), .O(n67789));
    defparam i51615_4_lut.LUT_INIT = 16'haaab;
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[21]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_LUT4 i22656_3_lut (.I0(n136), .I1(n188), .I2(n181), .I3(GND_net), 
            .O(n37022));
    defparam i22656_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[20]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[19]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[18]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[17]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[16]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[15]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[14]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[13]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[12]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[11]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_67[10]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[9]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[8]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[7]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[6]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[5]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[4]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[3]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[2]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_67[1]));   // verilog/TinyFPGA_B.v(323[10] 336[6])
    SB_DFFESR GLB_214 (.Q(INLB_c_0), .C(clk16MHz), .E(n28059), .D(GLB_N_499), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_216 (.Q(INLC_c_0), .C(clk16MHz), .E(n28059), .D(GLC_N_513), 
            .R(n29221));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i22657_3_lut (.I0(n37022), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(n37023));
    defparam i22657_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_8 (.CI(n52157), 
            .I0(n2528), .I1(VCC_net), .CO(n52158));
    SB_CARRY add_262_4 (.CI(n51338), .I0(duty[5]), .I1(n70691), .CO(n51339));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_5_lut (.I0(GND_net), 
            .I1(n1431), .I2(VCC_net), .I3(n51817), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_17 (.CI(n51634), .I0(n5416), .I1(n5441), .CO(n51635));
    SB_LUT4 add_262_3_lut (.I0(current[1]), .I1(duty[4]), .I2(n70691), 
            .I3(n51337), .O(n269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_1125_16_lut (.I0(GND_net), .I1(n5417), .I2(n5442), .I3(n51633), 
            .O(n427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_5 (.CI(n51817), 
            .I0(n1431), .I1(VCC_net), .CO(n51818));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_4_lut (.I0(GND_net), 
            .I1(n1432), .I2(GND_net), .I3(n51816), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_4 (.CI(n51816), 
            .I0(n1432), .I1(GND_net), .CO(n51817));
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5845), .I1(current_limit[9]), 
            .I2(n19), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_3_lut (.I0(GND_net), 
            .I1(n1433), .I2(VCC_net), .I3(n51815), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_10 (.CI(n51321), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n51322));
    SB_LUT4 i22658_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n37023), 
            .I2(control_update), .I3(GND_net), .O(n30810));   // verilog/motorControl.v(20[7:21])
    defparam i22658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_22_lut (.I0(GND_net), 
            .I1(n3114), .I2(VCC_net), .I3(n52324), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_3 (.CI(n51815), 
            .I0(n1433), .I1(VCC_net), .CO(n51816));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_967_2_lut (.I0(GND_net), 
            .I1(n939), .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_967_2 (.CI(VCC_net), 
            .I0(n939), .I1(GND_net), .CO(n51815));
    SB_CARRY add_1125_16 (.CI(n51633), .I0(n5417), .I1(n5442), .CO(n51634));
    SB_CARRY add_262_3 (.CI(n51337), .I0(duty[4]), .I1(n70691), .CO(n51338));
    SB_LUT4 add_1125_15_lut (.I0(GND_net), .I1(n5418), .I2(n5443), .I3(n51632), 
            .O(n428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_22 (.CI(n52324), 
            .I0(n3114), .I1(VCC_net), .CO(n52325));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_7_lut (.I0(GND_net), 
            .I1(n2529), .I2(GND_net), .I3(n52156), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_262_2_lut (.I0(GND_net), .I1(duty[3]), .I2(n211), .I3(GND_net), 
            .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_262_2 (.CI(GND_net), .I0(duty[3]), .I1(n211), .CO(n51337));
    SB_LUT4 add_264_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n51336), .O(encoder1_position_scaled_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_15 (.CI(n51632), .I0(n5418), .I1(n5443), .CO(n51633));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_7 (.CI(n52156), 
            .I0(n2529), .I1(GND_net), .CO(n52157));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_23_lut (.I0(GND_net), 
            .I1(n2813), .I2(VCC_net), .I3(n52244), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_6_lut (.I0(GND_net), 
            .I1(n2530), .I2(GND_net), .I3(n52155), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_6 (.CI(n52155), 
            .I0(n2530), .I1(GND_net), .CO(n52156));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_23 (.CI(n52244), 
            .I0(n2813), .I1(VCC_net), .CO(n52245));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_21_lut (.I0(GND_net), 
            .I1(n3115), .I2(VCC_net), .I3(n52323), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_14_lut (.I0(GND_net), .I1(n5419), .I2(n5444), .I3(n51631), 
            .O(n429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_21 (.CI(n52323), 
            .I0(n3115), .I1(VCC_net), .CO(n52324));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_20_lut (.I0(GND_net), 
            .I1(n3116), .I2(VCC_net), .I3(n52322), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_22_lut (.I0(GND_net), 
            .I1(n2814), .I2(VCC_net), .I3(n52243), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_5_lut (.I0(GND_net), 
            .I1(n2531), .I2(VCC_net), .I3(n52154), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16404_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(\PID_CONTROLLER.integral_23__N_3844 [17]), 
            .I2(control_update), .I3(GND_net), .O(n30811));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16404_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_22 (.CI(n52243), 
            .I0(n2814), .I1(VCC_net), .CO(n52244));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_20 (.CI(n52322), 
            .I0(n3116), .I1(VCC_net), .CO(n52323));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_19_lut (.I0(GND_net), 
            .I1(n3117), .I2(VCC_net), .I3(n52321), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_5 (.CI(n52154), 
            .I0(n2531), .I1(VCC_net), .CO(n52155));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_4_lut (.I0(GND_net), 
            .I1(n2532), .I2(GND_net), .I3(n52153), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_21_lut (.I0(GND_net), 
            .I1(n2815), .I2(VCC_net), .I3(n52242), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_21 (.CI(n52242), 
            .I0(n2815), .I1(VCC_net), .CO(n52243));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_19 (.CI(n52321), 
            .I0(n3117), .I1(VCC_net), .CO(n52322));
    SB_LUT4 i16405_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3844 [16]), 
            .I2(control_update), .I3(GND_net), .O(n30812));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16405_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_4 (.CI(n52153), 
            .I0(n2532), .I1(GND_net), .CO(n52154));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_3_lut (.I0(GND_net), 
            .I1(n2533), .I2(VCC_net), .I3(n52152), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_20_lut (.I0(GND_net), 
            .I1(n2816), .I2(VCC_net), .I3(n52241), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_20 (.CI(n52241), 
            .I0(n2816), .I1(VCC_net), .CO(n52242));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_18_lut (.I0(GND_net), 
            .I1(n3118), .I2(VCC_net), .I3(n52320), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_18 (.CI(n52320), 
            .I0(n3118), .I1(VCC_net), .CO(n52321));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i25_3_lut (.I0(encoder0_position_scaled_23__N_319[24]), 
            .I1(n9_adj_5955), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n934));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_3 (.CI(n52152), 
            .I0(n2533), .I1(VCC_net), .CO(n52153));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1704_2_lut (.I0(GND_net), 
            .I1(n950), .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_14 (.CI(n51631), .I0(n5419), .I1(n5444), .CO(n51632));
    SB_LUT4 LessThan_17_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1704_2 (.CI(VCC_net), 
            .I0(n950), .I1(GND_net), .CO(n52152));
    SB_LUT4 i53175_3_lut (.I0(n4), .I1(current_limit[5]), .I2(n11), .I3(GND_net), 
            .O(n69350));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53176_3_lut (.I0(n69350), .I1(current_limit[6]), .I2(n13), 
            .I3(GND_net), .O(n69351));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_24_lut (.I0(n70321), 
            .I1(n2412), .I2(VCC_net), .I3(n52151), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_23_lut (.I0(GND_net), 
            .I1(n2413), .I2(VCC_net), .I3(n52150), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_19_lut (.I0(GND_net), 
            .I1(n2817), .I2(VCC_net), .I3(n52240), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_17_lut (.I0(GND_net), 
            .I1(n3119), .I2(VCC_net), .I3(n52319), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_13_lut (.I0(GND_net), .I1(n5420), .I2(n5445), .I3(n51630), 
            .O(n430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_19 (.CI(n52240), 
            .I0(n2817), .I1(VCC_net), .CO(n52241));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_17 (.CI(n52319), 
            .I0(n3119), .I1(VCC_net), .CO(n52320));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_23 (.CI(n52150), 
            .I0(n2413), .I1(VCC_net), .CO(n52151));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_22_lut (.I0(GND_net), 
            .I1(n2414), .I2(VCC_net), .I3(n52149), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_22 (.CI(n52149), 
            .I0(n2414), .I1(VCC_net), .CO(n52150));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_16_lut (.I0(GND_net), 
            .I1(n3120), .I2(VCC_net), .I3(n52318), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_13 (.CI(n51630), .I0(n5420), .I1(n5445), .CO(n51631));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_21_lut (.I0(GND_net), 
            .I1(n2415), .I2(VCC_net), .I3(n52148), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51596_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n67789), 
            .O(n67770));
    defparam i51596_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_1125_12_lut (.I0(GND_net), .I1(n5421), .I2(n5446), .I3(n51629), 
            .O(n431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_12 (.CI(n51629), .I0(n5421), .I1(n5446), .CO(n51630));
    SB_LUT4 i16406_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3844 [15]), 
            .I2(control_update), .I3(GND_net), .O(n30813));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_18_lut (.I0(GND_net), 
            .I1(n2818), .I2(VCC_net), .I3(n52239), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_11_lut (.I0(GND_net), .I1(n5422), .I2(n5447), .I3(n51628), 
            .O(n432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_18 (.CI(n52239), 
            .I0(n2818), .I1(VCC_net), .CO(n52240));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_21 (.CI(n52148), 
            .I0(n2415), .I1(VCC_net), .CO(n52149));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_16 (.CI(n52318), 
            .I0(n3120), .I1(VCC_net), .CO(n52319));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_15_lut (.I0(GND_net), 
            .I1(n3121), .I2(VCC_net), .I3(n52317), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_11 (.CI(n51628), .I0(n5422), .I1(n5447), .CO(n51629));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_17_lut (.I0(GND_net), 
            .I1(n2819), .I2(VCC_net), .I3(n52238), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16407_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3844 [14]), 
            .I2(control_update), .I3(GND_net), .O(n30814));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_255), 
            .I3(n51412), .O(n356)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_20_lut (.I0(GND_net), 
            .I1(n2416), .I2(VCC_net), .I3(n52147), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_15 (.CI(n52317), 
            .I0(n3121), .I1(VCC_net), .CO(n52318));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_17 (.CI(n52238), 
            .I0(n2819), .I1(VCC_net), .CO(n52239));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_20 (.CI(n52147), 
            .I0(n2416), .I1(VCC_net), .CO(n52148));
    SB_LUT4 add_1125_10_lut (.I0(GND_net), .I1(n5423), .I2(n5448), .I3(n51627), 
            .O(n433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_19_lut (.I0(GND_net), 
            .I1(n2417), .I2(VCC_net), .I3(n52146), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_10 (.CI(n51627), .I0(n5423), .I1(n5448), .CO(n51628));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_14_lut (.I0(GND_net), 
            .I1(n3122), .I2(VCC_net), .I3(n52316), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_9_lut (.I0(GND_net), .I1(n5424), .I2(n5449), .I3(n51626), 
            .O(n434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_19 (.CI(n52146), 
            .I0(n2417), .I1(VCC_net), .CO(n52147));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_18_lut (.I0(GND_net), 
            .I1(n2418), .I2(VCC_net), .I3(n52145), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(n5246), .I1(GND_net), .I2(pwm_setpoint_23__N_255), 
            .I3(n51411), .O(n5411)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_14 (.CI(n52316), 
            .I0(n3122), .I1(VCC_net), .CO(n52317));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_16_lut (.I0(GND_net), 
            .I1(n2820), .I2(VCC_net), .I3(n52237), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_16 (.CI(n52237), 
            .I0(n2820), .I1(VCC_net), .CO(n52238));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_18 (.CI(n52145), 
            .I0(n2418), .I1(VCC_net), .CO(n52146));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_17_lut (.I0(GND_net), 
            .I1(n2419), .I2(VCC_net), .I3(n52144), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_13_lut (.I0(GND_net), 
            .I1(n3123), .I2(VCC_net), .I3(n52315), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_15_lut (.I0(GND_net), 
            .I1(n2821), .I2(VCC_net), .I3(n52236), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_19_lut (.I0(n70464), 
            .I1(n1917), .I2(VCC_net), .I3(n52008), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_13 (.CI(n52315), 
            .I0(n3123), .I1(VCC_net), .CO(n52316));
    SB_CARRY unary_minus_21_add_3_25 (.CI(n51411), .I0(GND_net), .I1(pwm_setpoint_23__N_255), 
            .CO(n51412));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_18_lut (.I0(GND_net), 
            .I1(n1918), .I2(VCC_net), .I3(n52007), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_17 (.CI(n52144), 
            .I0(n2419), .I1(VCC_net), .CO(n52145));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_18 (.CI(n52007), 
            .I0(n1918), .I1(VCC_net), .CO(n52008));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_16_lut (.I0(GND_net), 
            .I1(n2420), .I2(VCC_net), .I3(n52143), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_17_lut (.I0(GND_net), 
            .I1(n1919), .I2(VCC_net), .I3(n52006), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_17 (.CI(n52006), 
            .I0(n1919), .I1(VCC_net), .CO(n52007));
    SB_CARRY add_1125_9 (.CI(n51626), .I0(n5424), .I1(n5449), .CO(n51627));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_16_lut (.I0(GND_net), 
            .I1(n1920), .I2(VCC_net), .I3(n52005), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_12_lut (.I0(GND_net), 
            .I1(n3124), .I2(VCC_net), .I3(n52314), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_15 (.CI(n52236), 
            .I0(n2821), .I1(VCC_net), .CO(n52237));
    SB_LUT4 add_1125_8_lut (.I0(GND_net), .I1(n5425), .I2(n5450), .I3(n51625), 
            .O(n435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_16 (.CI(n52143), 
            .I0(n2420), .I1(VCC_net), .CO(n52144));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_15_lut (.I0(GND_net), 
            .I1(n2421), .I2(VCC_net), .I3(n52142), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2114_3_lut (.I0(n3111), 
            .I1(n3178), .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_16 (.CI(n52005), 
            .I0(n1920), .I1(VCC_net), .CO(n52006));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_15 (.CI(n52142), 
            .I0(n2421), .I1(VCC_net), .CO(n52143));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_14_lut (.I0(GND_net), 
            .I1(n2822), .I2(VCC_net), .I3(n52235), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16408_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3844 [13]), 
            .I2(control_update), .I3(GND_net), .O(n30815));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(n5246), .I1(GND_net), .I2(n3), 
            .I3(n51410), .O(n5412)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1125_8 (.CI(n51625), .I0(n5425), .I1(n5450), .CO(n51626));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_14 (.CI(n52235), 
            .I0(n2822), .I1(VCC_net), .CO(n52236));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_14_lut (.I0(GND_net), 
            .I1(n2422), .I2(VCC_net), .I3(n52141), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_7_lut (.I0(GND_net), .I1(n5426), .I2(n5451), .I3(n51624), 
            .O(n436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_14 (.CI(n52141), 
            .I0(n2422), .I1(VCC_net), .CO(n52142));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_13_lut (.I0(GND_net), 
            .I1(n2823), .I2(VCC_net), .I3(n52234), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_15_lut (.I0(GND_net), 
            .I1(n1921), .I2(VCC_net), .I3(n52004), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_15 (.CI(n52004), 
            .I0(n1921), .I1(VCC_net), .CO(n52005));
    SB_CARRY add_1125_7 (.CI(n51624), .I0(n5426), .I1(n5451), .CO(n51625));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_12 (.CI(n52314), 
            .I0(n3124), .I1(VCC_net), .CO(n52315));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_13_lut (.I0(GND_net), 
            .I1(n1323), .I2(VCC_net), .I3(n51792), .O(n1390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_6_lut (.I0(GND_net), .I1(n5427), .I2(n5452), .I3(n51623), 
            .O(n437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_12_lut (.I0(GND_net), 
            .I1(n1324), .I2(VCC_net), .I3(n51791), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_12 (.CI(n51791), 
            .I0(n1324), .I1(VCC_net), .CO(n51792));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [4]), 
            .O(n58849));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_14_lut (.I0(GND_net), 
            .I1(n1922), .I2(VCC_net), .I3(n52003), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_11_lut (.I0(GND_net), 
            .I1(n1325), .I2(VCC_net), .I3(n51790), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_11 (.CI(n51790), 
            .I0(n1325), .I1(VCC_net), .CO(n51791));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_10_lut (.I0(GND_net), 
            .I1(n1326), .I2(VCC_net), .I3(n51789), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_24 (.CI(n51410), .I0(GND_net), .I1(n3), 
            .CO(n51411));
    SB_CARRY add_1125_6 (.CI(n51623), .I0(n5427), .I1(n5452), .CO(n51624));
    SB_LUT4 i53464_4_lut (.I0(n16), .I1(n6), .I2(n19), .I3(n67768), 
            .O(n69639));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53464_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i22283_3_lut (.I0(n219), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844 [12]));
    defparam i22283_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_13 (.CI(n52234), 
            .I0(n2823), .I1(VCC_net), .CO(n52235));
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(n5246), .I1(GND_net), .I2(n4_adj_5849), 
            .I3(n51409), .O(n5413)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n51409), .I0(GND_net), .I1(n4_adj_5849), 
            .CO(n51410));
    SB_LUT4 i22284_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3844 [12]), 
            .I2(control_update), .I3(GND_net), .O(n30816));   // verilog/motorControl.v(20[7:21])
    defparam i22284_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_14 (.CI(n52003), 
            .I0(n1922), .I1(VCC_net), .CO(n52004));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_10 (.CI(n51789), 
            .I0(n1326), .I1(VCC_net), .CO(n51790));
    SB_LUT4 add_1125_5_lut (.I0(GND_net), .I1(n5428), .I2(n5453), .I3(n51622), 
            .O(n438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_11_lut (.I0(GND_net), 
            .I1(n3125), .I2(VCC_net), .I3(n52313), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_4 (.CI(n51315), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n51316));
    SB_LUT4 i51950_3_lut (.I0(n69351), .I1(current_limit[7]), .I2(n15), 
            .I3(GND_net), .O(n68124));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i51950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_9_lut (.I0(GND_net), 
            .I1(n1327), .I2(VCC_net), .I3(n51788), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(n5246), .I1(GND_net), .I2(n5_adj_5850), 
            .I3(n51408), .O(n5414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_12_lut (.I0(GND_net), 
            .I1(n2824), .I2(VCC_net), .I3(n52233), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_5 (.CI(n51622), .I0(n5428), .I1(n5453), .CO(n51623));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_13_lut (.I0(GND_net), 
            .I1(n2423), .I2(VCC_net), .I3(n52140), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_12 (.CI(n52233), 
            .I0(n2824), .I1(VCC_net), .CO(n52234));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_11 (.CI(n52313), 
            .I0(n3125), .I1(VCC_net), .CO(n52314));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_13 (.CI(n52140), 
            .I0(n2423), .I1(VCC_net), .CO(n52141));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_13_lut (.I0(GND_net), 
            .I1(n1923), .I2(VCC_net), .I3(n52002), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_9 (.CI(n51788), 
            .I0(n1327), .I1(VCC_net), .CO(n51789));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_8_lut (.I0(GND_net), 
            .I1(n1328), .I2(VCC_net), .I3(n51787), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_13 (.CI(n52002), 
            .I0(n1923), .I1(VCC_net), .CO(n52003));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_8 (.CI(n51787), 
            .I0(n1328), .I1(VCC_net), .CO(n51788));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_10_lut (.I0(GND_net), 
            .I1(n3126), .I2(VCC_net), .I3(n52312), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_7_lut (.I0(GND_net), 
            .I1(n1329), .I2(GND_net), .I3(n51786), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_12_lut (.I0(GND_net), 
            .I1(n1924), .I2(VCC_net), .I3(n52001), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1125_4_lut (.I0(GND_net), .I1(n5429), .I2(n5454), .I3(n51621), 
            .O(n439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_7 (.CI(n51786), 
            .I0(n1329), .I1(GND_net), .CO(n51787));
    SB_CARRY add_1125_4 (.CI(n51621), .I0(n5429), .I1(n5454), .CO(n51622));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_6_lut (.I0(GND_net), 
            .I1(n1330), .I2(GND_net), .I3(n51785), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_10 (.CI(n52312), 
            .I0(n3126), .I1(VCC_net), .CO(n52313));
    SB_LUT4 i53652_4_lut (.I0(n68124), .I1(n69639), .I2(n19), .I3(n67770), 
            .O(n69827));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53652_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_6 (.CI(n51785), 
            .I0(n1330), .I1(GND_net), .CO(n51786));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_12_lut (.I0(GND_net), 
            .I1(n2424), .I2(VCC_net), .I3(n52139), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_12 (.CI(n52001), 
            .I0(n1924), .I1(VCC_net), .CO(n52002));
    SB_LUT4 add_1125_3_lut (.I0(GND_net), .I1(n5430), .I2(n9_adj_6055), 
            .I3(n51620), .O(n440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1125_3 (.CI(n51620), .I0(n5430), .I1(n9_adj_6055), .CO(n51621));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_5_lut (.I0(GND_net), 
            .I1(n1331), .I2(VCC_net), .I3(n51784), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_5 (.CI(n51784), 
            .I0(n1331), .I1(VCC_net), .CO(n51785));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_12 (.CI(n52139), 
            .I0(n2424), .I1(VCC_net), .CO(n52140));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_11_lut (.I0(GND_net), 
            .I1(n2825), .I2(VCC_net), .I3(n52232), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_11_lut (.I0(GND_net), 
            .I1(n1925), .I2(VCC_net), .I3(n52000), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_11 (.CI(n52000), 
            .I0(n1925), .I1(VCC_net), .CO(n52001));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_11_lut (.I0(GND_net), 
            .I1(n2425), .I2(VCC_net), .I3(n52138), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_9_lut (.I0(GND_net), 
            .I1(n3127), .I2(VCC_net), .I3(n52311), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53653_3_lut (.I0(n69827), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n69828));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53653_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53592_3_lut (.I0(n69828), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53592_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_4_lut (.I0(GND_net), 
            .I1(n1332), .I2(GND_net), .I3(n51783), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n51408), .I0(GND_net), .I1(n5_adj_5850), 
            .CO(n51409));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_10_lut (.I0(GND_net), 
            .I1(n1926), .I2(VCC_net), .I3(n51999), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_4 (.CI(n51783), 
            .I0(n1332), .I1(GND_net), .CO(n51784));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_3_lut (.I0(GND_net), 
            .I1(n1333), .I2(VCC_net), .I3(n51782), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_9 (.CI(n52311), 
            .I0(n3127), .I1(VCC_net), .CO(n52312));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_11 (.CI(n52232), 
            .I0(n2825), .I1(VCC_net), .CO(n52233));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_3 (.CI(n51782), 
            .I0(n1333), .I1(VCC_net), .CO(n51783));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_900_2_lut (.I0(GND_net), 
            .I1(n938), .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_8_lut (.I0(GND_net), 
            .I1(n3128), .I2(VCC_net), .I3(n52310), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_10 (.CI(n51999), 
            .I0(n1926), .I1(VCC_net), .CO(n52000));
    SB_LUT4 i16410_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3844 [11]), 
            .I2(control_update), .I3(GND_net), .O(n30817));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16410_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_11 (.CI(n52138), 
            .I0(n2425), .I1(VCC_net), .CO(n52139));
    SB_LUT4 add_1125_2_lut (.I0(GND_net), .I1(n5431), .I2(n5456), .I3(GND_net), 
            .O(n441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1125_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_900_2 (.CI(VCC_net), 
            .I0(n938), .I1(GND_net), .CO(n51782));
    SB_LUT4 i1_4_lut_adj_1965 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n61264));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1965.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_8 (.CI(n52310), 
            .I0(n3128), .I1(VCC_net), .CO(n52311));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [5]), 
            .O(n58850));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(n5246), .I1(GND_net), .I2(n6_adj_5851), 
            .I3(n51407), .O(n5415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1125_2 (.CI(GND_net), .I0(n5431), .I1(n5456), .CO(n51620));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_7_lut (.I0(GND_net), 
            .I1(n3129), .I2(GND_net), .I3(n52309), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_9_lut (.I0(GND_net), 
            .I1(n1927), .I2(VCC_net), .I3(n51998), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_10_lut (.I0(GND_net), 
            .I1(n2426), .I2(VCC_net), .I3(n52137), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_21 (.CI(n51407), .I0(GND_net), .I1(n6_adj_5851), 
            .CO(n51408));
    SB_LUT4 unary_minus_19_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51619), .O(n330)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(n5246), .I1(GND_net), .I2(n7_adj_5852), 
            .I3(n51406), .O(n5416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_20 (.CI(n51406), .I0(GND_net), .I1(n7_adj_5852), 
            .CO(n51407));
    SB_LUT4 add_264_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n51335), .O(encoder1_position_scaled_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_10_lut (.I0(GND_net), 
            .I1(n2826), .I2(VCC_net), .I3(n52231), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_10 (.CI(n52137), 
            .I0(n2426), .I1(VCC_net), .CO(n52138));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_9 (.CI(n51998), 
            .I0(n1927), .I1(VCC_net), .CO(n51999));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_9_lut (.I0(GND_net), 
            .I1(n2427), .I2(VCC_net), .I3(n52136), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_24 (.CI(n51335), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n51336));
    SB_LUT4 unary_minus_19_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n51618), .O(n334)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_8_lut (.I0(GND_net), 
            .I1(n1928), .I2(VCC_net), .I3(n51997), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_8 (.CI(n51997), 
            .I0(n1928), .I1(VCC_net), .CO(n51998));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_7 (.CI(n52309), 
            .I0(n3129), .I1(GND_net), .CO(n52310));
    SB_LUT4 i1_4_lut_adj_1967 (.I0(current_limit[13]), .I1(n24), .I2(current_limit[14]), 
            .I3(current_limit[12]), .O(n61267));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1967.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1968 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n61267), .I3(n61264), .O(n296));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1968.LUT_INIT = 16'hb3a2;
    SB_LUT4 add_264_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n51320), .O(encoder1_position_scaled_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_7_lut (.I0(GND_net), 
            .I1(n1929), .I2(GND_net), .I3(n51996), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(n5246), .I1(GND_net), .I2(n8_adj_5853), 
            .I3(n51405), .O(n5417)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_19_add_3_14 (.CI(n51618), .I0(GND_net), .I1(n2), 
            .CO(n51619));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_9 (.CI(n52136), 
            .I0(n2427), .I1(VCC_net), .CO(n52137));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_7 (.CI(n51996), 
            .I0(n1929), .I1(GND_net), .CO(n51997));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_6_lut (.I0(GND_net), 
            .I1(n1930), .I2(GND_net), .I3(n51995), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_6_lut (.I0(GND_net), 
            .I1(n3130), .I2(GND_net), .I3(n52308), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n51334), .O(encoder1_position_scaled_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_6 (.CI(n52308), 
            .I0(n3130), .I1(GND_net), .CO(n52309));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_8_lut (.I0(GND_net), 
            .I1(n2428), .I2(VCC_net), .I3(n52135), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_6 (.CI(n51995), 
            .I0(n1930), .I1(GND_net), .CO(n51996));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_10 (.CI(n52231), 
            .I0(n2826), .I1(VCC_net), .CO(n52232));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_5_lut (.I0(GND_net), 
            .I1(n3131), .I2(VCC_net), .I3(n52307), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_5_lut (.I0(GND_net), 
            .I1(n1931), .I2(VCC_net), .I3(n51994), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_8 (.CI(n52135), 
            .I0(n2428), .I1(VCC_net), .CO(n52136));
    SB_CARRY unary_minus_21_add_3_19 (.CI(n51405), .I0(GND_net), .I1(n8_adj_5853), 
            .CO(n51406));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_9_lut (.I0(GND_net), 
            .I1(n2827), .I2(VCC_net), .I3(n52230), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_5 (.CI(n52307), 
            .I0(n3131), .I1(VCC_net), .CO(n52308));
    SB_LUT4 i16411_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3844 [10]), 
            .I2(control_update), .I3(GND_net), .O(n30818));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_7_lut (.I0(GND_net), 
            .I1(n2429), .I2(GND_net), .I3(n52134), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2578_25_lut (.I0(n70642), .I1(n2_adj_6019), .I2(n1059), 
            .I3(n52387), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_25_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_5 (.CI(n51994), 
            .I0(n1931), .I1(VCC_net), .CO(n51995));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_4_lut (.I0(GND_net), 
            .I1(n1932), .I2(GND_net), .I3(n51993), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_9 (.CI(n52230), 
            .I0(n2827), .I1(VCC_net), .CO(n52231));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1245_3_lut (.I0(n1826), 
            .I1(n1893), .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_19_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5863), 
            .I3(n51617), .O(n335)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(n5246), .I1(GND_net), .I2(n9_adj_5854), 
            .I3(n51404), .O(n5418)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_8_lut (.I0(GND_net), 
            .I1(n2828), .I2(VCC_net), .I3(n52229), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_13 (.CI(n51617), .I0(GND_net), .I1(n14_adj_5863), 
            .CO(n51618));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_4_lut (.I0(GND_net), 
            .I1(n3132), .I2(GND_net), .I3(n52306), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_4 (.CI(n52306), 
            .I0(n3132), .I1(GND_net), .CO(n52307));
    SB_LUT4 add_2578_24_lut (.I0(n70582), .I1(n2_adj_6019), .I2(n1158), 
            .I3(n52386), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_19_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5864), 
            .I3(n51616), .O(n336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_24 (.CI(n52386), .I0(n2_adj_6019), .I1(n1158), .CO(n52387));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_7 (.CI(n52134), 
            .I0(n2429), .I1(GND_net), .CO(n52135));
    SB_LUT4 add_2578_23_lut (.I0(n70599), .I1(n2_adj_6019), .I2(n1257), 
            .I3(n52385), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_262_17_lut (.I0(current[15]), .I1(duty[18]), .I2(n70691), 
            .I3(n51351), .O(n255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_262_17_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_6_lut (.I0(GND_net), 
            .I1(n2430), .I2(GND_net), .I3(n52133), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_8 (.CI(n52229), 
            .I0(n2828), .I1(VCC_net), .CO(n52230));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_4 (.CI(n51993), 
            .I0(n1932), .I1(GND_net), .CO(n51994));
    SB_CARRY unary_minus_19_add_3_12 (.CI(n51616), .I0(GND_net), .I1(n15_adj_5864), 
            .CO(n51617));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_6 (.CI(n52133), 
            .I0(n2430), .I1(GND_net), .CO(n52134));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_3_lut (.I0(GND_net), 
            .I1(n3133), .I2(VCC_net), .I3(n52305), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_23 (.CI(n52385), .I0(n2_adj_6019), .I1(n1257), .CO(n52386));
    SB_LUT4 add_2578_22_lut (.I0(n70629), .I1(n2_adj_6019), .I2(n1356), 
            .I3(n52384), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i30535_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n44839));
    defparam i30535_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16412_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3844 [9]), 
            .I2(control_update), .I3(GND_net), .O(n30819));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_19_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5865), 
            .I3(n51615), .O(n337)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_3_lut (.I0(GND_net), 
            .I1(n1933), .I2(VCC_net), .I3(n51992), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_3 (.CI(n51992), 
            .I0(n1933), .I1(VCC_net), .CO(n51993));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1302_2_lut (.I0(GND_net), 
            .I1(n944), .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_22 (.CI(n52384), .I0(n2_adj_6019), .I1(n1356), .CO(n52385));
    SB_CARRY add_264_23 (.CI(n51334), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n51335));
    SB_CARRY unary_minus_19_add_3_11 (.CI(n51615), .I0(GND_net), .I1(n16_adj_5865), 
            .CO(n51616));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1302_2 (.CI(VCC_net), 
            .I0(n944), .I1(GND_net), .CO(n51992));
    SB_LUT4 add_2578_21_lut (.I0(n70570), .I1(n2_adj_6019), .I2(n1455), 
            .I3(n52383), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_21_add_3_18 (.CI(n51404), .I0(GND_net), .I1(n9_adj_5854), 
            .CO(n51405));
    SB_LUT4 unary_minus_19_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5866), 
            .I3(n51614), .O(n338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_7_lut (.I0(GND_net), 
            .I1(n2829), .I2(GND_net), .I3(n52228), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(n5246), .I1(GND_net), .I2(n10_adj_5855), 
            .I3(n51403), .O(n5419)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [6]), 
            .O(n58844));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_19_add_3_10 (.CI(n51614), .I0(GND_net), .I1(n17_adj_5866), 
            .CO(n51615));
    SB_LUT4 LessThan_20_i13_2_lut (.I0(duty[6]), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5888));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2578_21 (.CI(n52383), .I0(n2_adj_6019), .I1(n1455), .CO(n52384));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_7 (.CI(n52228), 
            .I0(n2829), .I1(GND_net), .CO(n52229));
    SB_LUT4 i16413_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3844 [8]), 
            .I2(control_update), .I3(GND_net), .O(n30820));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i15_2_lut (.I0(duty[7]), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5887));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2578_20_lut (.I0(n70548), .I1(n2_adj_6019), .I2(n1554_adj_5994), 
            .I3(n52382), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_19_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5867), 
            .I3(n51613), .O(n339)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_3 (.CI(n52305), 
            .I0(n3133), .I1(VCC_net), .CO(n52306));
    SB_CARRY add_2578_20 (.CI(n52382), .I0(n2_adj_6019), .I1(n1554_adj_5994), 
            .CO(n52383));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_5_lut (.I0(GND_net), 
            .I1(n2431), .I2(VCC_net), .I3(n52132), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1970 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n63034));
    defparam i1_3_lut_adj_1970.LUT_INIT = 16'hfefe;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(duty[9]), .I1(n337), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5884));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_5 (.CI(n52132), 
            .I0(n2431), .I1(VCC_net), .CO(n52133));
    SB_LUT4 i16414_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3844 [7]), 
            .I2(control_update), .I3(GND_net), .O(n30821));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_6_lut (.I0(GND_net), 
            .I1(n2830), .I2(GND_net), .I3(n52227), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2106_2_lut (.I0(GND_net), 
            .I1(n956), .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(duty[8]), .I1(n338), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5885));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16415_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3844 [6]), 
            .I2(control_update), .I3(GND_net), .O(n30822));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i7_2_lut (.I0(duty[3]), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5892));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1971 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n63292));
    defparam i1_2_lut_adj_1971.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(duty[4]), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5890));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i11_2_lut (.I0(duty[5]), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5889));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i5_2_lut (.I0(duty[2]), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5894));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_4_lut (.I0(GND_net), 
            .I1(n2432), .I2(GND_net), .I3(n52131), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51659_4_lut (.I0(n11_adj_5889), .I1(n9_adj_5890), .I2(n7_adj_5892), 
            .I3(n5_adj_5894), .O(n67833));
    defparam i51659_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n342), .I1(n338), .I2(n17_adj_5885), 
            .I3(GND_net), .O(n8_adj_5891));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2106_2 (.CI(VCC_net), 
            .I0(n956), .I1(GND_net), .CO(n52305));
    SB_LUT4 add_2578_19_lut (.I0(n70527), .I1(n2_adj_6019), .I2(n1653), 
            .I3(n52381), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_21_add_3_17 (.CI(n51403), .I0(GND_net), .I1(n10_adj_5855), 
            .CO(n51404));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_4 (.CI(n52131), 
            .I0(n2432), .I1(GND_net), .CO(n52132));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_6 (.CI(n52227), 
            .I0(n2830), .I1(GND_net), .CO(n52228));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_30_lut (.I0(n70055), 
            .I1(n3006), .I2(VCC_net), .I3(n52304), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 LessThan_20_i6_3_lut (.I0(n344), .I1(n343), .I2(n7_adj_5892), 
            .I3(GND_net), .O(n6_adj_5893));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i16_3_lut (.I0(n8_adj_5891), .I1(n337), .I2(n19_adj_5884), 
            .I3(GND_net), .O(n16_adj_5886));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47889_3_lut (.I0(duty[21]), .I1(duty[14]), .I2(n330), .I3(GND_net), 
            .O(n64052));
    defparam i47889_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i47893_3_lut (.I0(duty[16]), .I1(duty[19]), .I2(n330), .I3(GND_net), 
            .O(n64056));
    defparam i47893_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i48028_4_lut (.I0(duty[22]), .I1(n64052), .I2(duty[15]), .I3(n330), 
            .O(n64193));
    defparam i48028_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 LessThan_20_i4_3_lut (.I0(n66923), .I1(n345), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5895));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53177_3_lut (.I0(n4_adj_5895), .I1(n341), .I2(n11_adj_5889), 
            .I3(GND_net), .O(n69352));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53178_3_lut (.I0(n69352), .I1(n340), .I2(n13_adj_5888), .I3(GND_net), 
            .O(n69353));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51647_4_lut (.I0(n17_adj_5885), .I1(n15_adj_5887), .I2(n13_adj_5888), 
            .I3(n67833), .O(n67821));
    defparam i51647_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53484_4_lut (.I0(n16_adj_5886), .I1(n6_adj_5893), .I2(n19_adj_5884), 
            .I3(n67819), .O(n69659));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53484_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51948_3_lut (.I0(n69353), .I1(n339), .I2(n15_adj_5887), .I3(GND_net), 
            .O(n68122));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53664_4_lut (.I0(n68122), .I1(n69659), .I2(n19_adj_5884), 
            .I3(n67821), .O(n69839));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53664_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53665_3_lut (.I0(n69839), .I1(n336), .I2(duty[10]), .I3(GND_net), 
            .O(n69840));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53665_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53588_3_lut (.I0(n69840), .I1(n335), .I2(duty[11]), .I3(GND_net), 
            .O(n69763));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53588_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i16416_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3844 [5]), 
            .I2(control_update), .I3(GND_net), .O(n30823));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i26_3_lut (.I0(n69763), .I1(n334), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_20_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7_4_lut (.I0(duty[20]), .I1(n26), .I2(n330), .I3(duty[23]), 
            .O(n20_adj_6079));
    defparam i7_4_lut.LUT_INIT = 16'h2100;
    SB_CARRY add_2578_19 (.CI(n52381), .I0(n2_adj_6019), .I1(n1653), .CO(n52382));
    SB_LUT4 i11_4_lut_adj_1972 (.I0(n330), .I1(n64193), .I2(n64056), .I3(duty[13]), 
            .O(n24_adj_6078));
    defparam i11_4_lut_adj_1972.LUT_INIT = 16'h0200;
    SB_LUT4 i51110_4_lut (.I0(duty[18]), .I1(n20_adj_6079), .I2(duty[17]), 
            .I3(n330), .O(n67072));
    defparam i51110_4_lut.LUT_INIT = 16'h8004;
    SB_LUT4 i2_2_lut_4_lut_4_lut (.I0(state_adj_6170[2]), .I1(state_adj_6170[3]), 
            .I2(state_adj_6170[0]), .I3(state_adj_6170[1]), .O(n6_adj_6010));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i2_2_lut_4_lut_4_lut.LUT_INIT = 16'hfdbd;
    SB_LUT4 i14_4_lut_adj_1973 (.I0(n67072), .I1(pwm_setpoint_23__N_255), 
            .I2(n296), .I3(n24_adj_6078), .O(n11999));
    defparam i14_4_lut_adj_1973.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_29_lut (.I0(GND_net), 
            .I1(n3007), .I2(VCC_net), .I3(n52303), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_5_lut (.I0(GND_net), 
            .I1(n2831), .I2(VCC_net), .I3(n52226), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_1106_i15_2_lut (.I0(r_Clock_Count_adj_6162[7]), .I1(o_Rx_DV_N_3617[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_6007));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1106_i9_2_lut (.I0(r_Clock_Count_adj_6162[4]), .I1(o_Rx_DV_N_3617[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_6004));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16417_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3844 [4]), 
            .I2(control_update), .I3(GND_net), .O(n30824));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1106_i13_2_lut (.I0(r_Clock_Count_adj_6162[6]), .I1(o_Rx_DV_N_3617[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_6006));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1106_i11_2_lut (.I0(r_Clock_Count_adj_6162[5]), .I1(o_Rx_DV_N_3617[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_6005));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[17] [7]), 
            .O(n58851));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_12_lut (.I0(n70599), 
            .I1(n1224), .I2(VCC_net), .I3(n51767), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_29 (.CI(n52303), 
            .I0(n3007), .I1(VCC_net), .CO(n52304));
    SB_CARRY unary_minus_19_add_3_9 (.CI(n51613), .I0(GND_net), .I1(n18_adj_5867), 
            .CO(n51614));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_11_lut (.I0(GND_net), 
            .I1(n1225), .I2(VCC_net), .I3(n51766), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_28_lut (.I0(GND_net), 
            .I1(n3008), .I2(VCC_net), .I3(n52302), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5868), 
            .I3(n51612), .O(n340)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_5 (.CI(n52226), 
            .I0(n2831), .I1(VCC_net), .CO(n52227));
    SB_LUT4 add_2578_18_lut (.I0(n70489), .I1(n2_adj_6019), .I2(n1752), 
            .I3(n52380), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_11 (.CI(n51766), 
            .I0(n1225), .I1(VCC_net), .CO(n51767));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_10_lut (.I0(GND_net), 
            .I1(n1226), .I2(VCC_net), .I3(n51765), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_10 (.CI(n51765), 
            .I0(n1226), .I1(VCC_net), .CO(n51766));
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(n5246), .I1(GND_net), .I2(n11_adj_5856), 
            .I3(n51402), .O(n5420)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_19_add_3_8 (.CI(n51612), .I0(GND_net), .I1(n19_adj_5868), 
            .CO(n51613));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_3_lut (.I0(GND_net), 
            .I1(n2433), .I2(VCC_net), .I3(n52130), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_16 (.CI(n51402), .I0(GND_net), .I1(n11_adj_5856), 
            .CO(n51403));
    SB_LUT4 unary_minus_19_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5869), 
            .I3(n51611), .O(n341)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_9_lut (.I0(GND_net), 
            .I1(n1227), .I2(VCC_net), .I3(n51764), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_9 (.CI(n51764), 
            .I0(n1227), .I1(VCC_net), .CO(n51765));
    SB_CARRY unary_minus_19_add_3_7 (.CI(n51611), .I0(GND_net), .I1(n20_adj_5869), 
            .CO(n51612));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_8_lut (.I0(GND_net), 
            .I1(n1228), .I2(VCC_net), .I3(n51763), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_9 (.CI(n51320), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n51321));
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(n5246), .I1(GND_net), .I2(n12), 
            .I3(n51401), .O(n5421)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_19_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5870), 
            .I3(n51610), .O(n342)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_3 (.CI(n52130), 
            .I0(n2433), .I1(VCC_net), .CO(n52131));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_8 (.CI(n51763), 
            .I0(n1228), .I1(VCC_net), .CO(n51764));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_7_lut (.I0(GND_net), 
            .I1(n1229), .I2(GND_net), .I3(n51762), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_19_add_3_6 (.CI(n51610), .I0(GND_net), .I1(n21_adj_5870), 
            .CO(n51611));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_7 (.CI(n51762), 
            .I0(n1229), .I1(GND_net), .CO(n51763));
    SB_LUT4 unary_minus_19_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5871), 
            .I3(n51609), .O(n343)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1637_2_lut (.I0(GND_net), 
            .I1(n949), .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_6_lut (.I0(GND_net), 
            .I1(n1230), .I2(GND_net), .I3(n51761), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_4_lut (.I0(GND_net), 
            .I1(n2832), .I2(GND_net), .I3(n52225), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_6 (.CI(n51761), 
            .I0(n1230), .I1(GND_net), .CO(n51762));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1637_2 (.CI(VCC_net), 
            .I0(n949), .I1(GND_net), .CO(n52130));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_5_lut (.I0(GND_net), 
            .I1(n1231), .I2(VCC_net), .I3(n51760), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_5 (.CI(n51760), 
            .I0(n1231), .I1(VCC_net), .CO(n51761));
    SB_CARRY unary_minus_19_add_3_5 (.CI(n51609), .I0(GND_net), .I1(n22_adj_5871), 
            .CO(n51610));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_4_lut (.I0(GND_net), 
            .I1(n1232), .I2(GND_net), .I3(n51759), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5872), 
            .I3(n51608), .O(n344)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n51333), .O(encoder1_position_scaled_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_4 (.CI(n51759), 
            .I0(n1232), .I1(GND_net), .CO(n51760));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_3_lut (.I0(GND_net), 
            .I1(n1233), .I2(VCC_net), .I3(n51758), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_3 (.CI(n51758), 
            .I0(n1233), .I1(VCC_net), .CO(n51759));
    SB_CARRY unary_minus_19_add_3_4 (.CI(n51608), .I0(GND_net), .I1(n23_adj_5872), 
            .CO(n51609));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_833_2_lut (.I0(GND_net), 
            .I1(n937), .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_19_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5873), 
            .I3(n51607), .O(n345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_18 (.CI(n52380), .I0(n2_adj_6019), .I1(n1752), .CO(n52381));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_28 (.CI(n52302), 
            .I0(n3008), .I1(VCC_net), .CO(n52303));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_833_2 (.CI(VCC_net), 
            .I0(n937), .I1(GND_net), .CO(n51758));
    SB_CARRY unary_minus_21_add_3_15 (.CI(n51401), .I0(GND_net), .I1(n12), 
            .CO(n51402));
    SB_CARRY unary_minus_19_add_3_3 (.CI(n51607), .I0(GND_net), .I1(n24_adj_5873), 
            .CO(n51608));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_4 (.CI(n52225), 
            .I0(n2832), .I1(GND_net), .CO(n52226));
    SB_LUT4 unary_minus_19_add_3_2_lut (.I0(n34987), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(n66923)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_19_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_23_lut (.I0(n70229), 
            .I1(n2313), .I2(VCC_net), .I3(n52129), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_19_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n51607));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_22_lut (.I0(GND_net), 
            .I1(n2314), .I2(VCC_net), .I3(n52128), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_22 (.CI(n51333), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n51334));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_22 (.CI(n52128), 
            .I0(n2314), .I1(VCC_net), .CO(n52129));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(n5246), .I1(GND_net), .I2(n13_adj_5857), 
            .I3(n51400), .O(n5422)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2578_17_lut (.I0(n70294), .I1(n2_adj_6019), .I2(n1851), 
            .I3(n52379), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_21_lut (.I0(GND_net), 
            .I1(n2315), .I2(VCC_net), .I3(n52127), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_17 (.CI(n52379), .I0(n2_adj_6019), .I1(n1851), .CO(n52380));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_21 (.CI(n52127), 
            .I0(n2315), .I1(VCC_net), .CO(n52128));
    SB_LUT4 add_264_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n51332), .O(encoder1_position_scaled_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_3_lut (.I0(GND_net), 
            .I1(n2833), .I2(VCC_net), .I3(n52224), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n51319), .O(encoder1_position_scaled_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_27_lut (.I0(GND_net), 
            .I1(n3009), .I2(VCC_net), .I3(n52301), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_27 (.CI(n52301), 
            .I0(n3009), .I1(VCC_net), .CO(n52302));
    SB_CARRY unary_minus_21_add_3_14 (.CI(n51400), .I0(GND_net), .I1(n13_adj_5857), 
            .CO(n51401));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_20_lut (.I0(GND_net), 
            .I1(n2316), .I2(VCC_net), .I3(n52126), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_3 (.CI(n52224), 
            .I0(n2833), .I1(VCC_net), .CO(n52225));
    SB_LUT4 add_264_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n51314), .O(encoder1_position_scaled_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1905_2_lut (.I0(GND_net), 
            .I1(n953), .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_20 (.CI(n52126), 
            .I0(n2316), .I1(VCC_net), .CO(n52127));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_26_lut (.I0(GND_net), 
            .I1(n3010), .I2(VCC_net), .I3(n52300), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1905_2 (.CI(VCC_net), 
            .I0(n953), .I1(GND_net), .CO(n52224));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_27_lut (.I0(n70259), 
            .I1(n2709), .I2(VCC_net), .I3(n52223), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_19_lut (.I0(GND_net), 
            .I1(n2317), .I2(VCC_net), .I3(n52125), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(n5246), .I1(GND_net), .I2(n14), 
            .I3(n51399), .O(n5423)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_21_add_3_13 (.CI(n51399), .I0(GND_net), .I1(n14), 
            .CO(n51400));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_26 (.CI(n52300), 
            .I0(n3010), .I1(VCC_net), .CO(n52301));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_19 (.CI(n52125), 
            .I0(n2317), .I1(VCC_net), .CO(n52126));
    SB_CARRY add_264_3 (.CI(n51314), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n51315));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_18_lut (.I0(GND_net), 
            .I1(n2318), .I2(VCC_net), .I3(n52124), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(n5246), .I1(GND_net), .I2(n15_adj_5858), 
            .I3(n51398), .O(n5424)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_18 (.CI(n52124), 
            .I0(n2318), .I1(VCC_net), .CO(n52125));
    SB_CARRY unary_minus_21_add_3_12 (.CI(n51398), .I0(GND_net), .I1(n15_adj_5858), 
            .CO(n51399));
    SB_CARRY add_264_8 (.CI(n51319), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n51320));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_25_lut (.I0(GND_net), 
            .I1(n3011), .I2(VCC_net), .I3(n52299), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_26_lut (.I0(GND_net), 
            .I1(n2710), .I2(VCC_net), .I3(n52222), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(n5246), .I1(GND_net), .I2(n16_adj_5859), 
            .I3(n51397), .O(n5425)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_264_21 (.CI(n51332), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n51333));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_26 (.CI(n52222), 
            .I0(n2710), .I1(VCC_net), .CO(n52223));
    SB_LUT4 add_264_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n51331), .O(encoder1_position_scaled_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_25 (.CI(n52299), 
            .I0(n3011), .I1(VCC_net), .CO(n52300));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_17_lut (.I0(GND_net), 
            .I1(n2319), .I2(VCC_net), .I3(n52123), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_25_lut (.I0(GND_net), 
            .I1(n2711), .I2(VCC_net), .I3(n52221), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_17 (.CI(n52123), 
            .I0(n2319), .I1(VCC_net), .CO(n52124));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_25 (.CI(n52221), 
            .I0(n2711), .I1(VCC_net), .CO(n52222));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_16_lut (.I0(GND_net), 
            .I1(n2320), .I2(VCC_net), .I3(n52122), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_11_lut (.I0(n70582), 
            .I1(n1125), .I2(VCC_net), .I3(n51738), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2578_16_lut (.I0(n70464), .I1(n2_adj_6019), .I2(n1950), 
            .I3(n52378), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_16 (.CI(n52122), 
            .I0(n2320), .I1(VCC_net), .CO(n52123));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_10_lut (.I0(GND_net), 
            .I1(n1126), .I2(VCC_net), .I3(n51737), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_10 (.CI(n51737), 
            .I0(n1126), .I1(VCC_net), .CO(n51738));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_9_lut (.I0(GND_net), 
            .I1(n1127), .I2(VCC_net), .I3(n51736), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_9 (.CI(n51736), 
            .I0(n1127), .I1(VCC_net), .CO(n51737));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_18_lut (.I0(n70294), 
            .I1(n1818), .I2(VCC_net), .I3(n51971), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_8_lut (.I0(GND_net), 
            .I1(n1128), .I2(VCC_net), .I3(n51735), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_8 (.CI(n51735), 
            .I0(n1128), .I1(VCC_net), .CO(n51736));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_7_lut (.I0(GND_net), 
            .I1(n1129), .I2(GND_net), .I3(n51734), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n51397), .I0(GND_net), .I1(n16_adj_5859), 
            .CO(n51398));
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(n5246), .I1(GND_net), .I2(n17_adj_5860), 
            .I3(n51396), .O(n5426)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_7 (.CI(n51734), 
            .I0(n1129), .I1(GND_net), .CO(n51735));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_24_lut (.I0(GND_net), 
            .I1(n2712), .I2(VCC_net), .I3(n52220), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_24 (.CI(n52220), 
            .I0(n2712), .I1(VCC_net), .CO(n52221));
    SB_CARRY unary_minus_21_add_3_10 (.CI(n51396), .I0(GND_net), .I1(n17_adj_5860), 
            .CO(n51397));
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(n5246), .I1(GND_net), .I2(n18), 
            .I3(n51395), .O(n5427)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_264_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_351), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_17_lut (.I0(GND_net), 
            .I1(n1819), .I2(VCC_net), .I3(n51970), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_6_lut (.I0(GND_net), 
            .I1(n1130), .I2(GND_net), .I3(n51733), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_15_lut (.I0(GND_net), 
            .I1(n2321), .I2(VCC_net), .I3(n52121), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n51318), .O(encoder1_position_scaled_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_20 (.CI(n51331), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n51332));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_6 (.CI(n51733), 
            .I0(n1130), .I1(GND_net), .CO(n51734));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_15 (.CI(n52121), 
            .I0(n2321), .I1(VCC_net), .CO(n52122));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_17 (.CI(n51970), 
            .I0(n1819), .I1(VCC_net), .CO(n51971));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_16_lut (.I0(GND_net), 
            .I1(n1820), .I2(VCC_net), .I3(n51969), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_5_lut (.I0(GND_net), 
            .I1(n1131), .I2(VCC_net), .I3(n51732), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_5 (.CI(n51732), 
            .I0(n1131), .I1(VCC_net), .CO(n51733));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_4_lut (.I0(GND_net), 
            .I1(n1132), .I2(GND_net), .I3(n51731), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_4 (.CI(n51731), 
            .I0(n1132), .I1(GND_net), .CO(n51732));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_24_lut (.I0(GND_net), 
            .I1(n3012), .I2(VCC_net), .I3(n52298), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_24 (.CI(n52298), 
            .I0(n3012), .I1(VCC_net), .CO(n52299));
    SB_CARRY add_264_7 (.CI(n51318), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n51319));
    SB_LUT4 add_264_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n51330), .O(encoder1_position_scaled_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n51395), .I0(GND_net), .I1(n18), 
            .CO(n51396));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_16 (.CI(n51969), 
            .I0(n1820), .I1(VCC_net), .CO(n51970));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [0]), 
            .O(n58852));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 add_264_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n51317), .O(encoder1_position_scaled_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(n5246), .I1(GND_net), .I2(n19_adj_5861), 
            .I3(n51394), .O(n5428)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_264_19 (.CI(n51330), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n51331));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_15_lut (.I0(GND_net), 
            .I1(n1821), .I2(VCC_net), .I3(n51968), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_3_lut (.I0(GND_net), 
            .I1(n1133), .I2(VCC_net), .I3(n51730), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_3 (.CI(n51730), 
            .I0(n1133), .I1(VCC_net), .CO(n51731));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_766_2_lut (.I0(GND_net), 
            .I1(n936), .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_14_lut (.I0(GND_net), 
            .I1(n2322), .I2(VCC_net), .I3(n52120), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_766_2 (.CI(VCC_net), 
            .I0(n936), .I1(GND_net), .CO(n51730));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_14 (.CI(n52120), 
            .I0(n2322), .I1(VCC_net), .CO(n52121));
    SB_CARRY add_2578_16 (.CI(n52378), .I0(n2_adj_6019), .I1(n1950), .CO(n52379));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_23_lut (.I0(GND_net), 
            .I1(n2713), .I2(VCC_net), .I3(n52219), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_15 (.CI(n51968), 
            .I0(n1821), .I1(VCC_net), .CO(n51969));
    SB_LUT4 add_2578_15_lut (.I0(n70433), .I1(n2_adj_6019), .I2(n2049), 
            .I3(n52377), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_14_lut (.I0(GND_net), 
            .I1(n1822), .I2(VCC_net), .I3(n51967), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_13_lut (.I0(GND_net), 
            .I1(n2323), .I2(VCC_net), .I3(n52119), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_23_lut (.I0(GND_net), 
            .I1(n3013), .I2(VCC_net), .I3(n52297), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_23 (.CI(n52219), 
            .I0(n2713), .I1(VCC_net), .CO(n52220));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_13 (.CI(n52119), 
            .I0(n2323), .I1(VCC_net), .CO(n52120));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_14 (.CI(n51967), 
            .I0(n1822), .I1(VCC_net), .CO(n51968));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_13_lut (.I0(GND_net), 
            .I1(n1823), .I2(VCC_net), .I3(n51966), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_22_lut (.I0(GND_net), 
            .I1(n2714), .I2(VCC_net), .I3(n52218), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_13 (.CI(n51966), 
            .I0(n1823), .I1(VCC_net), .CO(n51967));
    SB_CARRY unary_minus_21_add_3_8 (.CI(n51394), .I0(GND_net), .I1(n19_adj_5861), 
            .CO(n51395));
    SB_LUT4 add_264_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n51329), .O(encoder1_position_scaled_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_12_lut (.I0(GND_net), 
            .I1(n1824), .I2(VCC_net), .I3(n51965), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_351), 
            .CO(n51314));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_22 (.CI(n52218), 
            .I0(n2714), .I1(VCC_net), .CO(n52219));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_12_lut (.I0(GND_net), 
            .I1(n2324), .I2(VCC_net), .I3(n52118), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(n5246), .I1(GND_net), .I2(n20), 
            .I3(n51393), .O(n5429)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2578_15 (.CI(n52377), .I0(n2_adj_6019), .I1(n2049), .CO(n52378));
    SB_CARRY add_264_6 (.CI(n51317), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n51318));
    SB_CARRY add_264_18 (.CI(n51329), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n51330));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_12 (.CI(n52118), 
            .I0(n2324), .I1(VCC_net), .CO(n52119));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_23 (.CI(n52297), 
            .I0(n3013), .I1(VCC_net), .CO(n52298));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_12 (.CI(n51965), 
            .I0(n1824), .I1(VCC_net), .CO(n51966));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_21_lut (.I0(GND_net), 
            .I1(n2715), .I2(VCC_net), .I3(n52217), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_11_lut (.I0(GND_net), 
            .I1(n2325), .I2(VCC_net), .I3(n52117), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_22_lut (.I0(GND_net), 
            .I1(n3014), .I2(VCC_net), .I3(n52296), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_11_lut (.I0(GND_net), 
            .I1(n1825), .I2(VCC_net), .I3(n51964), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_11 (.CI(n51964), 
            .I0(n1825), .I1(VCC_net), .CO(n51965));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_10_lut (.I0(GND_net), 
            .I1(n1826), .I2(VCC_net), .I3(n51963), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_10 (.CI(n51963), 
            .I0(n1826), .I1(VCC_net), .CO(n51964));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_11 (.CI(n52117), 
            .I0(n2325), .I1(VCC_net), .CO(n52118));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_9_lut (.I0(GND_net), 
            .I1(n1827), .I2(VCC_net), .I3(n51962), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_9 (.CI(n51962), 
            .I0(n1827), .I1(VCC_net), .CO(n51963));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_8_lut (.I0(GND_net), 
            .I1(n1828), .I2(VCC_net), .I3(n51961), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_21 (.CI(n52217), 
            .I0(n2715), .I1(VCC_net), .CO(n52218));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n51393), .I0(GND_net), .I1(n20), 
            .CO(n51394));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_10_lut (.I0(GND_net), 
            .I1(n2326), .I2(VCC_net), .I3(n52116), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n51328), .O(encoder1_position_scaled_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_20_lut (.I0(GND_net), 
            .I1(n2716), .I2(VCC_net), .I3(n52216), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_10 (.CI(n52116), 
            .I0(n2326), .I1(VCC_net), .CO(n52117));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_8 (.CI(n51961), 
            .I0(n1828), .I1(VCC_net), .CO(n51962));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_20 (.CI(n52216), 
            .I0(n2716), .I1(VCC_net), .CO(n52217));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_7_lut (.I0(GND_net), 
            .I1(n1829), .I2(GND_net), .I3(n51960), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_9_lut (.I0(GND_net), 
            .I1(n2327), .I2(VCC_net), .I3(n52115), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(n5246), .I1(GND_net), .I2(n21), 
            .I3(n51392), .O(n5430)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_7 (.CI(n51960), 
            .I0(n1829), .I1(GND_net), .CO(n51961));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_6_lut (.I0(GND_net), 
            .I1(n1830), .I2(GND_net), .I3(n51959), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_19_lut (.I0(GND_net), 
            .I1(n2717), .I2(VCC_net), .I3(n52215), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_6 (.CI(n51959), 
            .I0(n1830), .I1(GND_net), .CO(n51960));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_22 (.CI(n52296), 
            .I0(n3014), .I1(VCC_net), .CO(n52297));
    SB_CARRY unary_minus_21_add_3_6 (.CI(n51392), .I0(GND_net), .I1(n21), 
            .CO(n51393));
    SB_CARRY add_264_17 (.CI(n51328), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n51329));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(n296), .I1(GND_net), .I2(n22), 
            .I3(n51391), .O(n5431)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n51391), .I0(GND_net), .I1(n22), 
            .CO(n51392));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_9 (.CI(n52115), 
            .I0(n2327), .I1(VCC_net), .CO(n52116));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_5_lut (.I0(GND_net), 
            .I1(n1831), .I2(VCC_net), .I3(n51958), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_21_lut (.I0(GND_net), 
            .I1(n3015), .I2(VCC_net), .I3(n52295), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n51327), .O(encoder1_position_scaled_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_16 (.CI(n51327), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n51328));
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(n379), .I1(GND_net), .I2(n23), 
            .I3(n51390), .O(n4_adj_5902)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_5 (.CI(n51958), 
            .I0(n1831), .I1(VCC_net), .CO(n51959));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_19 (.CI(n52215), 
            .I0(n2717), .I1(VCC_net), .CO(n52216));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_8_lut (.I0(GND_net), 
            .I1(n2328), .I2(VCC_net), .I3(n52114), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_4_lut (.I0(GND_net), 
            .I1(n1832), .I2(GND_net), .I3(n51957), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2578_14_lut (.I0(n70460), .I1(n2_adj_6019), .I2(n2148), 
            .I3(n52376), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_1106_i4_4_lut (.I0(r_Clock_Count_adj_6162[0]), .I1(o_Rx_DV_N_3617[1]), 
            .I2(r_Clock_Count_adj_6162[1]), .I3(o_Rx_DV_N_3617[0]), .O(n4_adj_6001));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i16418_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3844 [3]), 
            .I2(control_update), .I3(GND_net), .O(n30825));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16418_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_4 (.CI(n51957), 
            .I0(n1832), .I1(GND_net), .CO(n51958));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n51390), .I0(GND_net), .I1(n23), 
            .CO(n51391));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5862), 
            .I3(n51389), .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_3_lut (.I0(GND_net), 
            .I1(n1833), .I2(VCC_net), .I3(n51956), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_3 (.CI(n51956), 
            .I0(n1833), .I1(VCC_net), .CO(n51957));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_10_lut (.I0(GND_net), 
            .I1(n1026), .I2(VCC_net), .I3(n51717), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_8 (.CI(n52114), 
            .I0(n2328), .I1(VCC_net), .CO(n52115));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1235_2_lut (.I0(GND_net), 
            .I1(n943), .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_7_lut (.I0(GND_net), 
            .I1(n2329), .I2(GND_net), .I3(n52113), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_9_lut (.I0(GND_net), 
            .I1(n1027), .I2(VCC_net), .I3(n51716), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1235_2 (.CI(VCC_net), 
            .I0(n943), .I1(GND_net), .CO(n51956));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_9 (.CI(n51716), 
            .I0(n1027), .I1(VCC_net), .CO(n51717));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_8_lut (.I0(GND_net), 
            .I1(n1028), .I2(VCC_net), .I3(n51715), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_8 (.CI(n51715), 
            .I0(n1028), .I1(VCC_net), .CO(n51716));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_18_lut (.I0(GND_net), 
            .I1(n2718), .I2(VCC_net), .I3(n52214), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n51389), .I0(GND_net), .I1(n24_adj_5862), 
            .CO(n51390));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n4_adj_5902), .I1(GND_net), 
            .I2(n34987), .I3(VCC_net), .O(n66911)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n34987), 
            .CO(n51389));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_7_lut (.I0(GND_net), 
            .I1(n1029), .I2(GND_net), .I3(n51714), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_7 (.CI(n52113), 
            .I0(n2329), .I1(GND_net), .CO(n52114));
    SB_LUT4 add_264_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n51326), .O(encoder1_position_scaled_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_6_lut (.I0(GND_net), 
            .I1(n2330), .I2(GND_net), .I3(n52112), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_7 (.CI(n51714), 
            .I0(n1029), .I1(GND_net), .CO(n51715));
    SB_LUT4 add_174_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n51388), .O(n1531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_264_15 (.CI(n51326), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n51327));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_6_lut (.I0(GND_net), 
            .I1(n1030), .I2(GND_net), .I3(n51713), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_21 (.CI(n52295), 
            .I0(n3015), .I1(VCC_net), .CO(n52296));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_6 (.CI(n52112), 
            .I0(n2330), .I1(GND_net), .CO(n52113));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_6 (.CI(n51713), 
            .I0(n1030), .I1(GND_net), .CO(n51714));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_18 (.CI(n52214), 
            .I0(n2718), .I1(VCC_net), .CO(n52215));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_5_lut (.I0(GND_net), 
            .I1(n2331), .I2(VCC_net), .I3(n52111), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_5_lut (.I0(GND_net), 
            .I1(n1031), .I2(VCC_net), .I3(n51712), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_14 (.CI(n52376), .I0(n2_adj_6019), .I1(n2148), .CO(n52377));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_5 (.CI(n51712), 
            .I0(n1031), .I1(VCC_net), .CO(n51713));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_4_lut (.I0(GND_net), 
            .I1(n1032), .I2(GND_net), .I3(n51711), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_5 (.CI(n52111), 
            .I0(n2331), .I1(VCC_net), .CO(n52112));
    SB_LUT4 add_174_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n51387), .O(n1532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_4 (.CI(n51711), 
            .I0(n1032), .I1(GND_net), .CO(n51712));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_20_lut (.I0(GND_net), 
            .I1(n3016), .I2(VCC_net), .I3(n52294), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_17_lut (.I0(GND_net), 
            .I1(n2719), .I2(VCC_net), .I3(n52213), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_3_lut (.I0(GND_net), 
            .I1(n1033), .I2(VCC_net), .I3(n51710), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_4_lut (.I0(GND_net), 
            .I1(n2332), .I2(GND_net), .I3(n52110), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_174_32 (.CI(n51387), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n51388));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_3 (.CI(n51710), 
            .I0(n1033), .I1(VCC_net), .CO(n51711));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_699_2_lut (.I0(GND_net), 
            .I1(n935), .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_264_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n51325), .O(encoder1_position_scaled_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_264_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_4 (.CI(n52110), 
            .I0(n2332), .I1(GND_net), .CO(n52111));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_3_lut (.I0(GND_net), 
            .I1(n2333), .I2(VCC_net), .I3(n52109), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_699_2 (.CI(VCC_net), 
            .I0(n935), .I1(GND_net), .CO(n51710));
    SB_LUT4 add_2578_13_lut (.I0(n70182), .I1(n2_adj_6019), .I2(n2247), 
            .I3(n52375), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_174_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n51386), .O(n1533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53060_3_lut (.I0(n4_adj_6001), .I1(o_Rx_DV_N_3617[5]), .I2(n11_adj_6005), 
            .I3(GND_net), .O(n69235));   // verilog/uart_tx.v(117[17:57])
    defparam i53060_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_17 (.CI(n52213), 
            .I0(n2719), .I1(VCC_net), .CO(n52214));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_3 (.CI(n52109), 
            .I0(n2333), .I1(VCC_net), .CO(n52110));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1570_2_lut (.I0(GND_net), 
            .I1(n948), .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_20 (.CI(n52294), 
            .I0(n3016), .I1(VCC_net), .CO(n52295));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_19_lut (.I0(GND_net), 
            .I1(n3017), .I2(VCC_net), .I3(n52293), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_13 (.CI(n52375), .I0(n2_adj_6019), .I1(n2247), .CO(n52376));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_16_lut (.I0(GND_net), 
            .I1(n2720), .I2(VCC_net), .I3(n52212), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1570_2 (.CI(VCC_net), 
            .I0(n948), .I1(GND_net), .CO(n52109));
    SB_LUT4 add_2578_12_lut (.I0(n70229), .I1(n2_adj_6019), .I2(n2346), 
            .I3(n52374), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_22_lut (.I0(n70182), 
            .I1(n2214), .I2(VCC_net), .I3(n52108), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_16 (.CI(n52212), 
            .I0(n2720), .I1(VCC_net), .CO(n52213));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_21_lut (.I0(GND_net), 
            .I1(n2215), .I2(VCC_net), .I3(n52107), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_21 (.CI(n52107), 
            .I0(n2215), .I1(VCC_net), .CO(n52108));
    SB_CARRY add_2578_12 (.CI(n52374), .I0(n2_adj_6019), .I1(n2346), .CO(n52375));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_15_lut (.I0(GND_net), 
            .I1(n2721), .I2(VCC_net), .I3(n52211), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_19 (.CI(n52293), 
            .I0(n3017), .I1(VCC_net), .CO(n52294));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_15 (.CI(n52211), 
            .I0(n2721), .I1(VCC_net), .CO(n52212));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_20_lut (.I0(GND_net), 
            .I1(n2216), .I2(VCC_net), .I3(n52106), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_20 (.CI(n52106), 
            .I0(n2216), .I1(VCC_net), .CO(n52107));
    SB_CARRY add_174_31 (.CI(n51386), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n51387));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_14_lut (.I0(GND_net), 
            .I1(n2722), .I2(VCC_net), .I3(n52210), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_19_lut (.I0(GND_net), 
            .I1(n2217), .I2(VCC_net), .I3(n52105), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_19 (.CI(n52105), 
            .I0(n2217), .I1(VCC_net), .CO(n52106));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_18_lut (.I0(GND_net), 
            .I1(n3018), .I2(VCC_net), .I3(n52292), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_14 (.CI(n52210), 
            .I0(n2722), .I1(VCC_net), .CO(n52211));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_18_lut (.I0(GND_net), 
            .I1(n2218), .I2(VCC_net), .I3(n52104), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_18 (.CI(n52104), 
            .I0(n2218), .I1(VCC_net), .CO(n52105));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_18 (.CI(n52292), 
            .I0(n3018), .I1(VCC_net), .CO(n52293));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_13_lut (.I0(GND_net), 
            .I1(n2723), .I2(VCC_net), .I3(n52209), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_17_lut (.I0(GND_net), 
            .I1(n2219), .I2(VCC_net), .I3(n52103), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_17 (.CI(n52103), 
            .I0(n2219), .I1(VCC_net), .CO(n52104));
    SB_LUT4 add_174_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n51385), .O(n1534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_174_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2578_11_lut (.I0(n70321), .I1(n2_adj_6019), .I2(n2445), 
            .I3(n52373), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_17_lut (.I0(GND_net), 
            .I1(n3019), .I2(VCC_net), .I3(n52291), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_13 (.CI(n52209), 
            .I0(n2723), .I1(VCC_net), .CO(n52210));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_16_lut (.I0(GND_net), 
            .I1(n2220), .I2(VCC_net), .I3(n52102), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_11 (.CI(n52373), .I0(n2_adj_6019), .I1(n2445), .CO(n52374));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_16 (.CI(n52102), 
            .I0(n2220), .I1(VCC_net), .CO(n52103));
    SB_LUT4 add_2578_10_lut (.I0(n70372), .I1(n2_adj_6019), .I2(n2544), 
            .I3(n52372), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_12_lut (.I0(GND_net), 
            .I1(n2724), .I2(VCC_net), .I3(n52208), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_10 (.CI(n52372), .I0(n2_adj_6019), .I1(n2544), .CO(n52373));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_15_lut (.I0(GND_net), 
            .I1(n2221), .I2(VCC_net), .I3(n52101), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_17 (.CI(n52291), 
            .I0(n3019), .I1(VCC_net), .CO(n52292));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_15 (.CI(n52101), 
            .I0(n2221), .I1(VCC_net), .CO(n52102));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_16_lut (.I0(GND_net), 
            .I1(n3020), .I2(VCC_net), .I3(n52290), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_14_lut (.I0(GND_net), 
            .I1(n2222), .I2(VCC_net), .I3(n52100), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_16 (.CI(n52290), 
            .I0(n3020), .I1(VCC_net), .CO(n52291));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_12 (.CI(n52208), 
            .I0(n2724), .I1(VCC_net), .CO(n52209));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_14 (.CI(n52100), 
            .I0(n2222), .I1(VCC_net), .CO(n52101));
    SB_LUT4 add_2578_9_lut (.I0(n70401), .I1(n2_adj_6019), .I2(n2643), 
            .I3(n52371), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_11_lut (.I0(GND_net), 
            .I1(n2725), .I2(VCC_net), .I3(n52207), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_13_lut (.I0(GND_net), 
            .I1(n2223), .I2(VCC_net), .I3(n52099), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_17_lut (.I0(n70489), 
            .I1(n1719), .I2(VCC_net), .I3(n51927), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_13 (.CI(n52099), 
            .I0(n2223), .I1(VCC_net), .CO(n52100));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_16_lut (.I0(GND_net), 
            .I1(n1720), .I2(VCC_net), .I3(n51926), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_11 (.CI(n52207), 
            .I0(n2725), .I1(VCC_net), .CO(n52208));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_12_lut (.I0(GND_net), 
            .I1(n2224), .I2(VCC_net), .I3(n52098), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_16 (.CI(n51926), 
            .I0(n1720), .I1(VCC_net), .CO(n51927));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_15_lut (.I0(GND_net), 
            .I1(n1721), .I2(VCC_net), .I3(n51925), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_10_lut (.I0(GND_net), 
            .I1(n2726), .I2(VCC_net), .I3(n52206), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_12 (.CI(n52098), 
            .I0(n2224), .I1(VCC_net), .CO(n52099));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_15 (.CI(n51925), 
            .I0(n1721), .I1(VCC_net), .CO(n51926));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_14_lut (.I0(GND_net), 
            .I1(n1722), .I2(VCC_net), .I3(n51924), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_14 (.CI(n51924), 
            .I0(n1722), .I1(VCC_net), .CO(n51925));
    SB_CARRY add_264_14 (.CI(n51325), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n51326));
    SB_CARRY add_2578_9 (.CI(n52371), .I0(n2_adj_6019), .I1(n2643), .CO(n52372));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_15_lut (.I0(GND_net), 
            .I1(n3021), .I2(VCC_net), .I3(n52289), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_11_lut (.I0(GND_net), 
            .I1(n2225), .I2(VCC_net), .I3(n52097), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_10 (.CI(n52206), 
            .I0(n2726), .I1(VCC_net), .CO(n52207));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_11 (.CI(n52097), 
            .I0(n2225), .I1(VCC_net), .CO(n52098));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_13_lut (.I0(GND_net), 
            .I1(n1723), .I2(VCC_net), .I3(n51923), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_10_lut (.I0(GND_net), 
            .I1(n2226), .I2(VCC_net), .I3(n52096), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_13 (.CI(n51923), 
            .I0(n1723), .I1(VCC_net), .CO(n51924));
    SB_LUT4 add_2578_8_lut (.I0(n70259), .I1(n2_adj_6019), .I2(n2742), 
            .I3(n52370), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_12_lut (.I0(GND_net), 
            .I1(n1724), .I2(VCC_net), .I3(n51922), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_12 (.CI(n51922), 
            .I0(n1724), .I1(VCC_net), .CO(n51923));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_10 (.CI(n52096), 
            .I0(n2226), .I1(VCC_net), .CO(n52097));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_11_lut (.I0(GND_net), 
            .I1(n1725), .I2(VCC_net), .I3(n51921), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_9_lut (.I0(GND_net), 
            .I1(n2227), .I2(VCC_net), .I3(n52095), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_11 (.CI(n51921), 
            .I0(n1725), .I1(VCC_net), .CO(n51922));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_10_lut (.I0(GND_net), 
            .I1(n1726), .I2(VCC_net), .I3(n51920), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_10 (.CI(n51920), 
            .I0(n1726), .I1(VCC_net), .CO(n51921));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_9_lut (.I0(GND_net), 
            .I1(n1727), .I2(VCC_net), .I3(n51919), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_9 (.CI(n52095), 
            .I0(n2227), .I1(VCC_net), .CO(n52096));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_9_lut (.I0(GND_net), 
            .I1(n2727), .I2(VCC_net), .I3(n52205), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_9 (.CI(n51919), 
            .I0(n1727), .I1(VCC_net), .CO(n51920));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_9 (.CI(n52205), 
            .I0(n2727), .I1(VCC_net), .CO(n52206));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_8_lut (.I0(GND_net), 
            .I1(n2228), .I2(VCC_net), .I3(n52094), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_8 (.CI(n52370), .I0(n2_adj_6019), .I1(n2742), .CO(n52371));
    SB_LUT4 add_2578_7_lut (.I0(n70290), .I1(n2_adj_6019), .I2(n2841), 
            .I3(n52369), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_8_lut (.I0(GND_net), 
            .I1(n1728), .I2(VCC_net), .I3(n51918), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_7 (.CI(n52369), .I0(n2_adj_6019), .I1(n2841), .CO(n52370));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_8 (.CI(n52094), 
            .I0(n2228), .I1(VCC_net), .CO(n52095));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_6019), .I3(n52866), .O(n2_adj_5962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2578_6_lut (.I0(n70178), .I1(n2_adj_6019), .I2(n2940), 
            .I3(n52368), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i16419_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3844 [2]), 
            .I2(control_update), .I3(GND_net), .O(n30826));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53061_3_lut (.I0(n69235), .I1(o_Rx_DV_N_3617[6]), .I2(n13_adj_6006), 
            .I3(GND_net), .O(n69236));   // verilog/uart_tx.v(117[17:57])
    defparam i53061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_8_lut (.I0(GND_net), 
            .I1(n2728), .I2(VCC_net), .I3(n52204), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52380_4_lut (.I0(n13_adj_6006), .I1(n11_adj_6005), .I2(n9_adj_6004), 
            .I3(n67674), .O(n68554));
    defparam i52380_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_6020), .I3(n52865), .O(n3_adj_5961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_1106_i8_3_lut (.I0(n6_adj_6002), .I1(o_Rx_DV_N_3617[4]), 
            .I2(n9_adj_6004), .I3(GND_net), .O(n8_adj_6003));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_32 (.CI(n52865), 
            .I0(GND_net), .I1(n3_adj_6020), .CO(n52866));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_6021), .I3(n52864), .O(n4_adj_5960)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_31 (.CI(n52864), 
            .I0(GND_net), .I1(n4_adj_6021), .CO(n52865));
    SB_CARRY add_2578_6 (.CI(n52368), .I0(n2_adj_6019), .I1(n2940), .CO(n52369));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_6022), .I3(n52863), .O(n5_adj_5959)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_7_lut (.I0(GND_net), 
            .I1(n2229), .I2(GND_net), .I3(n52093), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_7 (.CI(n52093), 
            .I0(n2229), .I1(GND_net), .CO(n52094));
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_30 (.CI(n52863), 
            .I0(GND_net), .I1(n5_adj_6022), .CO(n52864));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_8 (.CI(n52204), 
            .I0(n2728), .I1(VCC_net), .CO(n52205));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_15 (.CI(n52289), 
            .I0(n3021), .I1(VCC_net), .CO(n52290));
    SB_LUT4 i52048_3_lut (.I0(n69236), .I1(o_Rx_DV_N_3617[7]), .I2(n15_adj_6007), 
            .I3(GND_net), .O(n68222));   // verilog/uart_tx.v(117[17:57])
    defparam i52048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53006_4_lut (.I0(n68222), .I1(n8_adj_6003), .I2(n15_adj_6007), 
            .I3(n68554), .O(n69181));   // verilog/uart_tx.v(117[17:57])
    defparam i53006_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53007_3_lut (.I0(n69181), .I1(o_Rx_DV_N_3617[8]), .I2(r_Clock_Count_adj_6162[8]), 
            .I3(GND_net), .O(n5257));   // verilog/uart_tx.v(117[17:57])
    defparam i53007_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_6023), .I3(n52862), .O(n6_adj_5958)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_29 (.CI(n52862), 
            .I0(GND_net), .I1(n6_adj_6023), .CO(n52863));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_6024), .I3(n52861), .O(n7_adj_5957)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_28 (.CI(n52861), 
            .I0(GND_net), .I1(n7_adj_6024), .CO(n52862));
    SB_LUT4 i16420_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3844 [1]), 
            .I2(control_update), .I3(GND_net), .O(n30827));   // verilog/motorControl.v(41[14] 61[8])
    defparam i16420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16421_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n23164), .I3(GND_net), .O(n30828));   // verilog/coms.v(130[12] 305[6])
    defparam i16421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [1]), 
            .O(n58846));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [2]), 
            .O(n58853));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1103_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3617[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_6014));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1103_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [3]), 
            .O(n58854));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [4]), 
            .O(n58855));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1103_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3617[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3617[0]), .O(n4_adj_6011));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1103_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1103_i8_3_lut (.I0(n6_adj_6012), .I1(o_Rx_DV_N_3617[4]), 
            .I2(n9_adj_6014), .I3(GND_net), .O(n8_adj_6013));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1103_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53440_4_lut (.I0(n8_adj_6013), .I1(n4_adj_6011), .I2(n9_adj_6014), 
            .I3(n67659), .O(n69615));   // verilog/uart_rx.v(119[17:57])
    defparam i53440_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53441_3_lut (.I0(n69615), .I1(o_Rx_DV_N_3617[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n69616));   // verilog/uart_rx.v(119[17:57])
    defparam i53441_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [5]), 
            .O(n58856));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i53348_3_lut (.I0(n69616), .I1(o_Rx_DV_N_3617[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n69523));   // verilog/uart_rx.v(119[17:57])
    defparam i53348_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_6025), .I3(n52860), .O(n8_adj_5956)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52076_3_lut (.I0(n69523), .I1(o_Rx_DV_N_3617[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5254));   // verilog/uart_rx.v(119[17:57])
    defparam i52076_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_27 (.CI(n52860), 
            .I0(GND_net), .I1(n8_adj_6025), .CO(n52861));
    SB_LUT4 i15683_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n30090));   // verilog/coms.v(130[12] 305[6])
    defparam i15683_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_6026), .I3(n52859), .O(n9_adj_5955)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_26 (.CI(n52859), 
            .I0(GND_net), .I1(n9_adj_6026), .CO(n52860));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_6027), .I3(n52858), .O(n10_adj_5954)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_25 (.CI(n52858), 
            .I0(GND_net), .I1(n10_adj_6027), .CO(n52859));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_6_lut (.I0(GND_net), 
            .I1(n2230), .I2(GND_net), .I3(n52092), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_6028), .I3(n52857), .O(n11_adj_5953)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_24 (.CI(n52857), 
            .I0(GND_net), .I1(n11_adj_6028), .CO(n52858));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_6029), .I3(n52856), .O(n12_adj_5952)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [6]), 
            .O(n58857));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[18] [7]), 
            .O(n58858));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_23 (.CI(n52856), 
            .I0(GND_net), .I1(n12_adj_6029), .CO(n52857));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_6030), .I3(n52855), .O(n13_adj_5951)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_22 (.CI(n52855), 
            .I0(GND_net), .I1(n13_adj_6030), .CO(n52856));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_6031), .I3(n52854), .O(n14_adj_5950)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2578_5_lut (.I0(n70055), .I1(n2_adj_6019), .I2(n3039), 
            .I3(n52367), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_7_lut (.I0(GND_net), 
            .I1(n2729), .I2(GND_net), .I3(n52203), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_21 (.CI(n52854), 
            .I0(GND_net), .I1(n14_adj_6031), .CO(n52855));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_6032), .I3(n52853), .O(n15_adj_5949)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_14_lut (.I0(GND_net), 
            .I1(n3022), .I2(VCC_net), .I3(n52288), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_20 (.CI(n52853), 
            .I0(GND_net), .I1(n15_adj_6032), .CO(n52854));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_6033), .I3(n52852), .O(n16_adj_5948)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_19 (.CI(n52852), 
            .I0(GND_net), .I1(n16_adj_6033), .CO(n52853));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_6034), .I3(n52851), .O(n17_adj_5947)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_18 (.CI(n52851), 
            .I0(GND_net), .I1(n17_adj_6034), .CO(n52852));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_6035), .I3(n52850), .O(n18_adj_5946)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_17 (.CI(n52850), 
            .I0(GND_net), .I1(n18_adj_6035), .CO(n52851));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_6036), .I3(n52849), .O(n19_adj_5945)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_16 (.CI(n52849), 
            .I0(GND_net), .I1(n19_adj_6036), .CO(n52850));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_6037), .I3(n52848), .O(n20_adj_5944)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_15 (.CI(n52848), 
            .I0(GND_net), .I1(n20_adj_6037), .CO(n52849));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_6 (.CI(n52092), 
            .I0(n2230), .I1(GND_net), .CO(n52093));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_6038), .I3(n52847), .O(n21_adj_5943)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_14 (.CI(n52847), 
            .I0(GND_net), .I1(n21_adj_6038), .CO(n52848));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [0]), 
            .O(n58859));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_5_lut (.I0(GND_net), 
            .I1(n2231), .I2(VCC_net), .I3(n52091), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_6039), .I3(n52846), .O(n22_adj_5942)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [1]), 
            .O(n58827));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [2]), 
            .O(n58860));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [3]), 
            .O(n58861));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_13 (.CI(n52846), 
            .I0(GND_net), .I1(n22_adj_6039), .CO(n52847));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_6040), .I3(n52845), .O(n23_adj_5941)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_9_lut (.I0(n960), 
            .I1(n927), .I2(VCC_net), .I3(n51693), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [4]), 
            .O(n58862));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_12 (.CI(n52845), 
            .I0(GND_net), .I1(n23_adj_6040), .CO(n52846));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1312_3_lut (.I0(n1925), 
            .I1(n1992), .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2110_3_lut (.I0(n3107), 
            .I1(n3174), .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2043_3_lut (.I0(n3008), 
            .I1(n3075), .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2046_3_lut (.I0(n3011), 
            .I1(n3078), .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [5]), 
            .O(n58863));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2045_3_lut (.I0(n3010), 
            .I1(n3077), .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2044_3_lut (.I0(n3009), 
            .I1(n3076), .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2049_3_lut (.I0(n3014), 
            .I1(n3081), .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51464_3_lut (.I0(state_7__N_4237[0]), .I1(n11_adj_5913), .I2(enable_slow_N_4340), 
            .I3(GND_net), .O(n67126));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i51464_3_lut.LUT_INIT = 16'h4c4c;
    SB_CARRY add_2578_5 (.CI(n52367), .I0(n2_adj_6019), .I1(n3039), .CO(n52368));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_14 (.CI(n52288), 
            .I0(n3022), .I1(VCC_net), .CO(n52289));
    SB_LUT4 i16_4_lut_adj_1989 (.I0(state_adj_6170[0]), .I1(n67126), .I2(n6878), 
            .I3(n6_adj_6010), .O(n8_adj_6087));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_1989.LUT_INIT = 16'h3afa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2048_3_lut (.I0(n3013), 
            .I1(n3080), .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2047_3_lut (.I0(n3012), 
            .I1(n3079), .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2051_3_lut (.I0(n3016), 
            .I1(n3083), .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2050_3_lut (.I0(n3015), 
            .I1(n3082), .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1990 (.I0(hall3), .I1(commutation_state[1]), .I2(hall2), 
            .I3(hall1), .O(n58640));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_1990.LUT_INIT = 16'hd054;
    SB_LUT4 add_2578_4_lut (.I0(n70089), .I1(n2_adj_6019), .I2(n3138), 
            .I3(n52366), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_13_lut (.I0(GND_net), 
            .I1(n3023), .I2(VCC_net), .I3(n52287), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_8 (.CI(n51918), 
            .I0(n1728), .I1(VCC_net), .CO(n51919));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2054_3_lut (.I0(n3019), 
            .I1(n3086), .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2053_3_lut (.I0(n3018), 
            .I1(n3085), .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_13 (.CI(n52287), 
            .I0(n3023), .I1(VCC_net), .CO(n52288));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2052_3_lut (.I0(n3017), 
            .I1(n3084), .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2067_3_lut (.I0(n3032), 
            .I1(n3099), .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2066_3_lut (.I0(n3031), 
            .I1(n3098), .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_6041), .I3(n52844), .O(n24_adj_5940)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2578_4 (.CI(n52366), .I0(n2_adj_6019), .I1(n3138), .CO(n52367));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2065_3_lut (.I0(n3030), 
            .I1(n3097), .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2062_3_lut (.I0(n3027), 
            .I1(n3094), .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16434_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[0]), 
            .I2(n10_adj_6065), .I3(n49984), .O(n30841));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16434_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2055_3_lut (.I0(n3020), 
            .I1(n3087), .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2061_3_lut (.I0(n3026), 
            .I1(n3093), .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2063_3_lut (.I0(n3028), 
            .I1(n3095), .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2059_3_lut (.I0(n3024), 
            .I1(n3091), .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2060_3_lut (.I0(n3025), 
            .I1(n3092), .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1795_3_lut (.I0(n2632), 
            .I1(n2699), .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_11 (.CI(n52844), 
            .I0(GND_net), .I1(n24_adj_6041), .CO(n52845));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_6042), .I3(n52843), .O(n25_adj_5939)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i43883_3_lut (.I0(reset), .I1(n8_adj_5908), .I2(n59093), .I3(GND_net), 
            .O(n60009));
    defparam i43883_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2058_3_lut (.I0(n3023), 
            .I1(n3090), .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2056_3_lut (.I0(n3021), 
            .I1(n3088), .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16435_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n60009), 
            .I3(GND_net), .O(n30842));   // verilog/coms.v(130[12] 305[6])
    defparam i16435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2057_3_lut (.I0(n3022), 
            .I1(n3089), .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2064_3_lut (.I0(n3029), 
            .I1(n3096), .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i13_3_lut (.I0(encoder0_position_scaled_23__N_319[12]), 
            .I1(n21_adj_5943), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16440_3_lut (.I0(n60079), .I1(r_Bit_Index_adj_6163[0]), .I2(n28320), 
            .I3(GND_net), .O(n30847));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i16440_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i16443_3_lut (.I0(n60053), .I1(r_Bit_Index[0]), .I2(n28324), 
            .I3(GND_net), .O(n30850));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16443_3_lut.LUT_INIT = 16'h1414;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_10 (.CI(n52843), 
            .I0(GND_net), .I1(n25_adj_6042), .CO(n52844));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_6043), .I3(n52842), .O(n26_adj_5938)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_12_lut (.I0(GND_net), 
            .I1(n3024), .I2(VCC_net), .I3(n52286), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1168_7_lut (.I0(GND_net), 
            .I1(n1729), .I2(GND_net), .I3(n51917), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_5 (.CI(n52091), 
            .I0(n2231), .I1(VCC_net), .CO(n52092));
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_9 (.CI(n52842), 
            .I0(GND_net), .I1(n26_adj_6043), .CO(n52843));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_12 (.CI(n52286), 
            .I0(n3024), .I1(VCC_net), .CO(n52287));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_6044), .I3(n52841), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_7 (.CI(n52203), 
            .I0(n2729), .I1(GND_net), .CO(n52204));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1503_4_lut (.I0(GND_net), 
            .I1(n2232), .I2(GND_net), .I3(n52090), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_8 (.CI(n52841), 
            .I0(GND_net), .I1(n27_adj_6044), .CO(n52842));
    SB_LUT4 add_2578_3_lut (.I0(n70125), .I1(n2_adj_6019), .I2(n3237), 
            .I3(n52365), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_6045), .I3(n52840), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_11_lut (.I0(GND_net), 
            .I1(n3025), .I2(VCC_net), .I3(n52285), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1168_7 (.CI(n51917), 
            .I0(n1729), .I1(GND_net), .CO(n51918));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_11 (.CI(n52285), 
            .I0(n3025), .I1(VCC_net), .CO(n52286));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_10_lut (.I0(GND_net), 
            .I1(n3026), .I2(VCC_net), .I3(n52284), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1524_3_lut (.I0(n2233), 
            .I1(n2300), .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1591_3_lut (.I0(n2332), 
            .I1(n2399), .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_7 (.CI(n52840), 
            .I0(GND_net), .I1(n28_adj_6045), .CO(n52841));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1379_3_lut (.I0(n2024), 
            .I1(n2091), .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1658_3_lut (.I0(n2431), 
            .I1(n2498), .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1725_3_lut (.I0(n2530), 
            .I1(n2597), .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_6046), .I3(n52839), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1792_3_lut (.I0(n2629), 
            .I1(n2696), .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1859_3_lut (.I0(n2728), 
            .I1(n2795), .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_6 (.CI(n52839), 
            .I0(GND_net), .I1(n29_adj_6046), .CO(n52840));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_6047), .I3(n52838), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53731_3_lut (.I0(\data_out_frame[15] [7]), .I1(n54003), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n69906));
    defparam i53731_3_lut.LUT_INIT = 16'h6969;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_5 (.CI(n52838), 
            .I0(GND_net), .I1(n30_adj_6047), .CO(n52839));
    SB_LUT4 i1_3_lut_adj_1991 (.I0(n2815), .I1(n2824), .I2(n2828), .I3(GND_net), 
            .O(n63730));
    defparam i1_3_lut_adj_1991.LUT_INIT = 16'hfefe;
    SB_LUT4 i30551_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n44855));
    defparam i30551_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_6048), .I3(n52837), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1992 (.I0(n2816), .I1(n2817), .I2(n2825), .I3(n2821), 
            .O(n63624));
    defparam i1_4_lut_adj_1992.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1993 (.I0(n2812), .I1(n2813), .I2(n2814), .I3(n63730), 
            .O(n63736));
    defparam i1_4_lut_adj_1993.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_4 (.CI(n52837), 
            .I0(GND_net), .I1(n31_adj_6048), .CO(n52838));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_6049), .I3(n52836), .O(n32_adj_5937)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1926_3_lut (.I0(n2827), 
            .I1(n2894), .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16447_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n62796), 
            .I3(n27_adj_5989), .O(n30854));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16447_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1976_3_lut (.I0(n2909), 
            .I1(n2976), .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16448_4_lut (.I0(CS_MISO_c), .I1(data_adj_6147[0]), .I2(n11_adj_5928), 
            .I3(state_7__N_4446), .O(n30855));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16448_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1975_3_lut (.I0(n2908), 
            .I1(n2975), .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1979_3_lut (.I0(n2912), 
            .I1(n2979), .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54420_4_lut (.I0(n63292), .I1(n1125), .I2(n63034), .I3(n44839), 
            .O(n1158));
    defparam i54420_4_lut.LUT_INIT = 16'h0103;
    SB_CARRY add_2578_3 (.CI(n52365), .I0(n2_adj_6019), .I1(n3237), .CO(n52366));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1978_3_lut (.I0(n2911), 
            .I1(n2978), .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_10 (.CI(n52284), 
            .I0(n3026), .I1(VCC_net), .CO(n52285));
    SB_LUT4 add_2578_2_lut (.I0(n70130), .I1(n2_adj_6019), .I2(n44815), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2578_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1977_3_lut (.I0(n2910), 
            .I1(n2977), .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1982_3_lut (.I0(n2915), 
            .I1(n2982), .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1981_3_lut (.I0(n2914), 
            .I1(n2981), .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1980_3_lut (.I0(n2913), 
            .I1(n2980), .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [6]), 
            .O(n58864));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_9_lut (.I0(GND_net), 
            .I1(n3027), .I2(VCC_net), .I3(n52283), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1983_3_lut (.I0(n2916), 
            .I1(n2983), .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1997_3_lut (.I0(n2930), 
            .I1(n2997), .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1985_3_lut (.I0(n2918), 
            .I1(n2985), .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30_4_lut (.I0(state_7__N_4045[0]), .I1(n5_adj_6076), .I2(state_adj_6139[1]), 
            .I3(n6_adj_6075), .O(n12_adj_6088));   // verilog/eeprom.v(35[8] 81[4])
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12_adj_6088), .I1(n67130), .I2(state_adj_6139[0]), 
            .I3(state_adj_6139[2]), .O(n58352));   // verilog/eeprom.v(35[8] 81[4])
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_3 (.CI(n52836), 
            .I0(GND_net), .I1(n32_adj_6049), .CO(n52837));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1984_3_lut (.I0(n2917), 
            .I1(n2984), .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_9 (.CI(n52283), 
            .I0(n3027), .I1(VCC_net), .CO(n52284));
    SB_CARRY add_2578_2 (.CI(VCC_net), .I0(n2_adj_6019), .I1(n44815), 
            .CO(n52365));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_8_lut (.I0(GND_net), 
            .I1(n3028), .I2(VCC_net), .I3(n52282), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[0] [2]), 
            .O(n58845));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2000_3_lut (.I0(n2933), 
            .I1(n3000), .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1999_3_lut (.I0(n2932), 
            .I1(n2999), .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i12_3_lut (.I0(encoder0_position_scaled_23__N_319[11]), 
            .I1(n22_adj_5942), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[0] [3]), 
            .O(n59003));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_33_lut (.I0(GND_net), 
            .I1(n3204), .I2(VCC_net), .I3(n52364), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1592_3_lut (.I0(n2333), 
            .I1(n2400), .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_8 (.CI(n52282), 
            .I0(n3028), .I1(VCC_net), .CO(n52283));
    SB_LUT4 i15653_3_lut_4_lut (.I0(n2275), .I1(b_prev_adj_5931), .I2(a_new_adj_6125[1]), 
            .I3(position_31__N_3956_adj_5932), .O(n30060));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15653_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2039_7_lut (.I0(GND_net), 
            .I1(n3029), .I2(GND_net), .I3(n52281), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_1838_6_lut (.I0(GND_net), 
            .I1(n2730), .I2(GND_net), .I3(n52202), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_6050), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15651_3_lut_4_lut (.I0(n2234), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3956), .O(n30058));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15651_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1659_3_lut (.I0(n2432), 
            .I1(n2499), .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1726_3_lut (.I0(n2531), 
            .I1(n2598), .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1997 (.I0(n63624), .I1(n2829), .I2(n44855), .I3(n2830), 
            .O(n63626));
    defparam i1_4_lut_adj_1997.LUT_INIT = 16'heaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_632_8_lut (.I0(GND_net), 
            .I1(n928), .I2(VCC_net), .I3(n51692), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_228_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_6050), .CO(n52836));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1503_4 (.CI(n52090), 
            .I0(n2232), .I1(GND_net), .CO(n52091));
    SB_LUT4 encoder0_position_scaled_23__I_0_228_add_2173_32_lut (.I0(GND_net), 
            .I1(n3205), .I2(VCC_net), .I3(n52363), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_228_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_1838_6 (.CI(n52202), 
            .I0(n2730), .I1(GND_net), .CO(n52203));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_2039_7 (.CI(n52281), 
            .I0(n3029), .I1(GND_net), .CO(n52282));
    SB_CARRY encoder0_position_scaled_23__I_0_228_add_632_8 (.CI(n51692), 
            .I0(n928), .I1(VCC_net), .CO(n51693));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[19] [7]), 
            .O(n58865));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1793_3_lut (.I0(n2630), 
            .I1(n2697), .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1860_3_lut (.I0(n2729), 
            .I1(n2796), .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i11_3_lut (.I0(encoder0_position_scaled_23__N_319[10]), 
            .I1(n23_adj_5941), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1660_3_lut (.I0(n2433), 
            .I1(n2500), .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1727_3_lut (.I0(n2532), 
            .I1(n2599), .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51162_4_lut (.I0(data_ready), .I1(n7082), .I2(n24_adj_6072), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n67067));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i51162_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1794_3_lut (.I0(n2631), 
            .I1(n2698), .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1861_3_lut (.I0(n2730), 
            .I1(n2797), .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1928_3_lut (.I0(n2829), 
            .I1(n2896), .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1999 (.I0(n2826), .I1(n2822), .I2(n2827), .I3(n2823), 
            .O(n63614));
    defparam i1_4_lut_adj_1999.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2000 (.I0(n2811), .I1(n63626), .I2(n2810), .I3(n63736), 
            .O(n63628));
    defparam i1_4_lut_adj_2000.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51699_2_lut (.I0(n24_adj_6072), .I1(n7082), .I2(GND_net), 
            .I3(GND_net), .O(n67070));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i51699_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n67070), .I1(n67067), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_6089), .O(n57536));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[0] [4]), 
            .O(n59002));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 i30471_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n44775));
    defparam i30471_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [0]), 
            .O(n58866));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [0]), 
            .O(n59001));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2004 (.I0(n2818), .I1(n63614), .I2(n2819), .I3(n2820), 
            .O(n63618));
    defparam i1_4_lut_adj_2004.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1927_3_lut (.I0(n2828), 
            .I1(n2895), .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1994_3_lut (.I0(n2927), 
            .I1(n2994), .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2005 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n63344));
    defparam i1_3_lut_adj_2005.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1986_3_lut (.I0(n2919), 
            .I1(n2986), .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54118_4_lut (.I0(n2808), .I1(n63618), .I2(n63628), .I3(n2809), 
            .O(n2841));
    defparam i54118_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1995_3_lut (.I0(n2928), 
            .I1(n2995), .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1862_3_lut (.I0(n2731), 
            .I1(n2798), .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i14_3_lut (.I0(encoder0_position_scaled_23__N_319[13]), 
            .I1(n20_adj_5944), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1930_3_lut (.I0(n2831), 
            .I1(n2898), .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2006 (.I0(n1229), .I1(n44775), .I2(n1230), .I3(n1231), 
            .O(n60702));
    defparam i1_4_lut_adj_2006.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1929_3_lut (.I0(n2830), 
            .I1(n2897), .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1456_3_lut (.I0(n2133), 
            .I1(n2200), .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [1]), 
            .O(n59000));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1523_3_lut (.I0(n2232), 
            .I1(n2299), .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1590_3_lut (.I0(n2331), 
            .I1(n2398), .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1657_3_lut (.I0(n2430), 
            .I1(n2497), .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [3]), 
            .O(n58999));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1724_3_lut (.I0(n2529), 
            .I1(n2596), .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1921_3_lut (.I0(n2822), 
            .I1(n2889), .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1791_3_lut (.I0(n2628), 
            .I1(n2695), .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54438_4_lut (.I0(n1225), .I1(n1224), .I2(n60702), .I3(n63344), 
            .O(n1257));
    defparam i54438_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1924_3_lut (.I0(n2825), 
            .I1(n2892), .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1858_3_lut (.I0(n2727), 
            .I1(n2794), .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [1]), 
            .O(n29319));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [2]), 
            .O(n29318));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [5]), 
            .O(n58998));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i902_3_lut (.I0(n1323), .I1(n1390), 
            .I2(n1356), .I3(GND_net), .O(n1422));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2012 (.I0(n2927), .I1(n2925), .I2(n2923), .I3(n2928), 
            .O(n63048));
    defparam i1_4_lut_adj_2012.LUT_INIT = 16'hfffe;
    SB_LUT4 i15627_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_6161[1]), 
            .I2(r_SM_Main_adj_6161[2]), .I3(n6_adj_6068), .O(n30034));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15627_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [6]), 
            .O(n58997));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1925_3_lut (.I0(n2826), 
            .I1(n2893), .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [7]), 
            .O(n58970));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i19_3_lut (.I0(encoder0_position_scaled_23__N_319[18]), 
            .I1(n15_adj_5949), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554_adj_5994), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [0]), 
            .O(n58969));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1116_3_lut (.I0(n1633), 
            .I1(n1700), .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1183_3_lut (.I0(n1732), 
            .I1(n1799), .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1250_3_lut (.I0(n1831), 
            .I1(n1898), .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1317_3_lut (.I0(n1930), 
            .I1(n1997), .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1384_3_lut (.I0(n2029), 
            .I1(n2096), .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1451_3_lut (.I0(n2128), 
            .I1(n2195), .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1518_3_lut (.I0(n2227), 
            .I1(n2294), .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1585_3_lut (.I0(n2326), 
            .I1(n2393), .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1652_3_lut (.I0(n2425), 
            .I1(n2492), .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30209_2_lut (.I0(duty[17]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5439));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30209_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1719_3_lut (.I0(n2524), 
            .I1(n2591), .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1786_3_lut (.I0(n2623), 
            .I1(n2690), .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1853_3_lut (.I0(n2722), 
            .I1(n2789), .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1920_3_lut (.I0(n2821), 
            .I1(n2888), .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15086_4_lut (.I0(n28100), .I1(n1642), .I2(n66915), .I3(n43962), 
            .O(n29464));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i15086_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1987_3_lut (.I0(n2920), 
            .I1(n2987), .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1988_3_lut (.I0(n2921), 
            .I1(n2988), .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1992_3_lut (.I0(n2925), 
            .I1(n2992), .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1991_3_lut (.I0(n2924), 
            .I1(n2991), .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i16_3_lut (.I0(encoder0_position_scaled_23__N_319[15]), 
            .I1(n18_adj_5946), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2016 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[1] [7]), 
            .O(n58996));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2016.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[3] [1]), 
            .O(n58995));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1320_3_lut (.I0(n1933), 
            .I1(n2000), .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1387_3_lut (.I0(n2032), 
            .I1(n2099), .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1454_3_lut (.I0(n2131), 
            .I1(n2198), .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1521_3_lut (.I0(n2230), 
            .I1(n2297), .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1588_3_lut (.I0(n2329), 
            .I1(n2396), .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2018 (.I0(n2922), .I1(n2920), .I2(n2926), .I3(GND_net), 
            .O(n63046));
    defparam i1_3_lut_adj_2018.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1655_3_lut (.I0(n2428), 
            .I1(n2495), .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1722_3_lut (.I0(n2527), 
            .I1(n2594), .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1789_3_lut (.I0(n2626), 
            .I1(n2693), .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1856_3_lut (.I0(n2725), 
            .I1(n2792), .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[3] [3]), 
            .O(n58994));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i17_3_lut (.I0(encoder0_position_scaled_23__N_319[16]), 
            .I1(n17_adj_5947), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2020 (.I0(n63048), .I1(n2924), .I2(n2921), .I3(GND_net), 
            .O(n63050));
    defparam i1_3_lut_adj_2020.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1252_3_lut (.I0(n1833), 
            .I1(n1900), .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1319_3_lut (.I0(n1932), 
            .I1(n1999), .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1386_3_lut (.I0(n2031), 
            .I1(n2098), .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1453_3_lut (.I0(n2130), 
            .I1(n2197), .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[3] [4]), 
            .O(n58842));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1520_3_lut (.I0(n2229), 
            .I1(n2296), .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1587_3_lut (.I0(n2328), 
            .I1(n2395), .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1654_3_lut (.I0(n2427), 
            .I1(n2494), .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1721_3_lut (.I0(n2526), 
            .I1(n2593), .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1788_3_lut (.I0(n2625), 
            .I1(n2692), .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1855_3_lut (.I0(n2724), 
            .I1(n2791), .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1922_3_lut (.I0(n2823), 
            .I1(n2890), .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1923_3_lut (.I0(n2824), 
            .I1(n2891), .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1990_3_lut (.I0(n2923), 
            .I1(n2990), .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15514_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n62846), 
            .I3(n27_adj_5989), .O(n29921));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15514_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1989_3_lut (.I0(n2922), 
            .I1(n2989), .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1996_3_lut (.I0(n2929), 
            .I1(n2996), .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1993_3_lut (.I0(n2926), 
            .I1(n2993), .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2022 (.I0(n3025), .I1(n3028), .I2(n3021), .I3(n3022), 
            .O(n63680));
    defparam i1_4_lut_adj_2022.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2023 (.I0(n3023), .I1(n3024), .I2(n3020), .I3(n3019), 
            .O(n63678));
    defparam i1_4_lut_adj_2023.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2024 (.I0(n63680), .I1(n3027), .I2(n3018), .I3(n3026), 
            .O(n63682));
    defparam i1_4_lut_adj_2024.LUT_INIT = 16'hfffe;
    SB_LUT4 i30547_4_lut (.I0(n955), .I1(n3031), .I2(n3032), .I3(n3033), 
            .O(n44851));
    defparam i30547_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2025 (.I0(n3016), .I1(n63682), .I2(n3017), .I3(n63678), 
            .O(n63688));
    defparam i1_4_lut_adj_2025.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2026 (.I0(n3029), .I1(n3030), .I2(GND_net), .I3(GND_net), 
            .O(n63794));
    defparam i1_2_lut_adj_2026.LUT_INIT = 16'h8888;
    SB_LUT4 i30483_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n44787));
    defparam i30483_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2027 (.I0(n3015), .I1(n63794), .I2(n63688), .I3(n44851), 
            .O(n63692));
    defparam i1_4_lut_adj_2027.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_2028 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n63692), 
            .O(n63698));
    defparam i1_4_lut_adj_2028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2029 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n63698), 
            .O(n63704));
    defparam i1_4_lut_adj_2029.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1045_3_lut (.I0(n1530), 
            .I1(n1597), .I2(n1554_adj_5994), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53883_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n63704), 
            .O(n3039));
    defparam i53883_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i4_3_lut (.I0(encoder0_position_scaled_23__N_319[3]), 
            .I1(n30), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n955));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2030 (.I0(n2918), .I1(n63050), .I2(n2919), .I3(n63046), 
            .O(n63056));
    defparam i1_4_lut_adj_2030.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2068_3_lut (.I0(n3033), 
            .I1(n3100), .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i3_3_lut (.I0(encoder0_position_scaled_23__N_319[2]), 
            .I1(n31), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n956));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30477_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n44781));
    defparam i30477_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2031 (.I0(n3128), .I1(n3121), .I2(n3120), .I3(n3122), 
            .O(n63192));
    defparam i1_4_lut_adj_2031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [3]), 
            .O(n29317));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2033 (.I0(n3124), .I1(n3123), .I2(n3127), .I3(n3125), 
            .O(n63194));
    defparam i1_4_lut_adj_2033.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2034 (.I0(n63194), .I1(n63192), .I2(n3119), .I3(n3126), 
            .O(n63198));
    defparam i1_4_lut_adj_2034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[3] [6]), 
            .O(n58993));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[3] [7]), 
            .O(n58992));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2037 (.I0(n3129), .I1(n44781), .I2(n3130), .I3(n3131), 
            .O(n60806));
    defparam i1_4_lut_adj_2037.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1112_3_lut (.I0(n1629), 
            .I1(n1696), .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2038 (.I0(n3116), .I1(n3117), .I2(n63198), .I3(n3118), 
            .O(n63204));
    defparam i1_4_lut_adj_2038.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2039 (.I0(n3114), .I1(n3115), .I2(n63204), .I3(n60806), 
            .O(n63210));
    defparam i1_4_lut_adj_2039.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2040 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n63210), 
            .O(n63216));
    defparam i1_4_lut_adj_2040.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2041 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n63216), 
            .O(n63222));
    defparam i1_4_lut_adj_2041.LUT_INIT = 16'hfffe;
    SB_LUT4 i53917_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n63222), 
            .O(n3138));
    defparam i53917_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2042_3_lut (.I0(n3007), 
            .I1(n3074), .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2109_3_lut (.I0(n3106), 
            .I1(n3173), .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [0]), 
            .O(n58991));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1446_3_lut (.I0(n2123), 
            .I1(n2190), .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [1]), 
            .O(n58990));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1513_3_lut (.I0(n2222), 
            .I1(n2289), .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1580_3_lut (.I0(n2321), 
            .I1(n2388), .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [2]), 
            .O(n58989));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1647_3_lut (.I0(n2420), 
            .I1(n2487), .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [3]), 
            .O(n58988));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [4]), 
            .O(n58867));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 i30208_2_lut (.I0(duty[18]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5438));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30208_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1714_3_lut (.I0(n2519), 
            .I1(n2586), .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [5]), 
            .O(n58868));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h2300;
    SB_LUT4 i5_3_lut_adj_2048 (.I0(r_SM_Main_adj_6161[0]), .I1(o_Rx_DV_N_3617[24]), 
            .I2(n27_adj_5989), .I3(GND_net), .O(n14_adj_6080));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut_adj_2048.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut_adj_2049 (.I0(n29_adj_5988), .I1(o_Rx_DV_N_3617[12]), 
            .I2(n23_adj_5990), .I3(n5257), .O(n15_adj_6077));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut_adj_2049.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut_adj_2050 (.I0(n15_adj_6077), .I1(n1), .I2(n14_adj_6080), 
            .I3(r_SM_Main_adj_6161[1]), .O(n71131));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut_adj_2050.LUT_INIT = 16'h8000;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1781_3_lut (.I0(n2618), 
            .I1(n2685), .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [4]), 
            .O(n58987));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 i15603_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n23230), .I3(GND_net), .O(n30010));   // verilog/coms.v(130[12] 305[6])
    defparam i15603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2052 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [5]), 
            .O(n58986));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2052.LUT_INIT = 16'h2300;
    SB_LUT4 i15605_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3844 [0]), 
            .I2(control_update), .I3(GND_net), .O(n30012));   // verilog/motorControl.v(41[14] 61[8])
    defparam i15605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15606_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n78), .I3(GND_net), .O(n30013));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15606_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15607_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n78), .I3(GND_net), .O(n30014));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15607_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [6]), 
            .O(n58985));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 i15608_3_lut (.I0(ID[0]), .I1(data_adj_6138[0]), .I2(n59065), 
            .I3(GND_net), .O(n30015));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2054 (.I0(n2929), .I1(n44787), .I2(n2930), .I3(n2931), 
            .O(n60797));
    defparam i1_4_lut_adj_2054.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_2055 (.I0(n3_adj_6054), .I1(data_ready), .I2(n25956), 
            .I3(state_adj_6139[2]), .O(n58524));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_2055.LUT_INIT = 16'hcec0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[4] [7]), 
            .O(n58984));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [6]), 
            .O(n58869));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    SB_LUT4 i15616_3_lut (.I0(current[0]), .I1(data_adj_6147[0]), .I2(n28109), 
            .I3(GND_net), .O(n30023));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15617_4_lut (.I0(rw), .I1(state_adj_6139[1]), .I2(state_adj_6139[2]), 
            .I3(n6196), .O(n30024));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15617_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15618_3_lut (.I0(CS_c), .I1(state_adj_6149[0]), .I2(state_adj_6149[1]), 
            .I3(GND_net), .O(n30025));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15618_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i54510_4_lut (.I0(n15_adj_5916), .I1(clk_out), .I2(state_adj_6149[0]), 
            .I3(state_adj_6149[1]), .O(n9_adj_6085));   // verilog/tli4970.v(35[10] 68[6])
    defparam i54510_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [0]), 
            .O(n58840));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h2300;
    SB_LUT4 i15634_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[1]), 
            .I2(n10_adj_6065), .I3(n25984), .O(n30041));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15634_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15635_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[2]), 
            .I2(n4_adj_5910), .I3(n49984), .O(n30042));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15635_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2059 (.I0(hall1), .I1(commutation_state[2]), .I2(hall3), 
            .I3(hall2), .O(n58604));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_4_lut_adj_2059.LUT_INIT = 16'hd054;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1179_3_lut (.I0(n1728), 
            .I1(n1795), .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15640_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[3]), 
            .I2(n4_adj_5910), .I3(n25984), .O(n30047));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15640_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2060 (.I0(n2916), .I1(n2917), .I2(n60797), .I3(n63056), 
            .O(n63062));
    defparam i1_4_lut_adj_2060.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15642_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[5]), 
            .I2(n4_adj_5911), .I3(n25984), .O(n30049));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15642_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1246_3_lut (.I0(n1827), 
            .I1(n1894), .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [1]), 
            .O(n58839));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1042_3_lut (.I0(n1527), 
            .I1(n1594), .I2(n1554_adj_5994), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15647_4_lut (.I0(state_7__N_4253[3]), .I1(data_adj_6138[7]), 
            .I2(n44006), .I3(n25984), .O(n30054));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15647_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i3_4_lut_adj_2062 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62_adj_5997), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n62248));
    defparam i3_4_lut_adj_2062.LUT_INIT = 16'h0004;
    SB_LUT4 i15650_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n23164), .I3(GND_net), .O(n30057));   // verilog/coms.v(130[12] 305[6])
    defparam i15650_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i15652_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n23164), .I3(GND_net), .O(n30059));   // verilog/coms.v(130[12] 305[6])
    defparam i15652_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(1)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n2270(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .b_prev(b_prev), .\a_new[1] (a_new[1]), 
            .n30058(n30058), .n2234(n2234), .position_31__N_3956(position_31__N_3956)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[49] 310[6])
    SB_LUT4 i15654_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n23164), .I3(GND_net), .O(n30061));   // verilog/coms.v(130[12] 305[6])
    defparam i15654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15655_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n23164), .I3(GND_net), .O(n30062));   // verilog/coms.v(130[12] 305[6])
    defparam i15655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15659_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n23164), .I3(GND_net), .O(n30066));   // verilog/coms.v(130[12] 305[6])
    defparam i15659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15660_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n23164), .I3(GND_net), .O(n30067));   // verilog/coms.v(130[12] 305[6])
    defparam i15660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15661_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n23164), .I3(GND_net), .O(n30068));   // verilog/coms.v(130[12] 305[6])
    defparam i15661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1109_3_lut (.I0(n1626), 
            .I1(n1693), .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1176_3_lut (.I0(n1725), 
            .I1(n1792), .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23792_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n23164), .I3(GND_net), .O(n30072));
    defparam i23792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15666_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n23164), .I3(GND_net), .O(n30073));   // verilog/coms.v(130[12] 305[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [2]), 
            .O(n58983));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2064 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [3]), 
            .O(n58982));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2064.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1103_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3617[3]), 
            .I2(o_Rx_DV_N_3617[2]), .I3(GND_net), .O(n6_adj_6012));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1103_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51485_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3617[3]), 
            .I2(o_Rx_DV_N_3617[2]), .I3(r_Clock_Count[2]), .O(n67659));   // verilog/uart_rx.v(119[17:57])
    defparam i51485_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [4]), 
            .O(n58981));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [7]), 
            .O(n58870));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1243_3_lut (.I0(n1824), 
            .I1(n1891), .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2067 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [0]), 
            .O(n58871));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2067.LUT_INIT = 16'h2300;
    SB_LUT4 i51500_3_lut_4_lut (.I0(r_Clock_Count_adj_6162[3]), .I1(o_Rx_DV_N_3617[3]), 
            .I2(o_Rx_DV_N_3617[2]), .I3(r_Clock_Count_adj_6162[2]), .O(n67674));   // verilog/uart_tx.v(117[17:57])
    defparam i51500_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1106_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_6162[3]), 
            .I1(o_Rx_DV_N_3617[3]), .I2(o_Rx_DV_N_3617[2]), .I3(GND_net), 
            .O(n6_adj_6002));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1106_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1310_3_lut (.I0(n1923), 
            .I1(n1990), .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [1]), 
            .O(n58968));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [1]), 
            .O(n29311));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2070 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [2]), 
            .O(n58872));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2070.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2071 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [3]), 
            .O(n58873));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2071.LUT_INIT = 16'h2300;
    SB_LUT4 i15667_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n23164), .I3(GND_net), .O(n30074));   // verilog/coms.v(130[12] 305[6])
    defparam i15667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53768_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n43842), .I3(GND_net), .O(n28100));
    defparam i53768_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i29458_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n23164), .I3(GND_net), .O(n30075));
    defparam i29458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51050_2_lut_3_lut (.I0(n62_adj_5997), .I1(delay_counter[31]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n66915));
    defparam i51050_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i29667_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n43842), .I3(GND_net), .O(n43962));
    defparam i29667_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2072 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [4]), 
            .O(n58874));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2072.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [5]), 
            .O(n58875));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_2074 (.I0(\data_out_frame[5] [1]), .I1(n59593), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n26490));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_2074.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2075 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [6]), 
            .O(n58876));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2075.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2076 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[21] [7]), 
            .O(n58877));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2076.LUT_INIT = 16'h2300;
    SB_LUT4 i5_2_lut_adj_2077 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26087));   // verilog/coms.v(100[12:26])
    defparam i5_2_lut_adj_2077.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2078 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [0]), 
            .O(n58878));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2078.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62_adj_5997), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_6089));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1642), .I3(n43842), .O(n24_adj_6072));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_adj_2079 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n63062), 
            .O(n63068));
    defparam i1_4_lut_adj_2079.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1313_3_lut (.I0(n1926), 
            .I1(n1993), .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2080 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [1]), 
            .O(n58879));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2080.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2081 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [2]), 
            .O(n58838));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2081.LUT_INIT = 16'h2300;
    SB_LUT4 i51802_2_lut_3_lut (.I0(enable_slow_N_4340), .I1(ready_prev), 
            .I2(state_adj_6139[1]), .I3(GND_net), .O(n67130));   // verilog/eeprom.v(35[8] 81[4])
    defparam i51802_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1377_3_lut (.I0(n2022), 
            .I1(n2089), .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2082 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n63068), 
            .O(n63074));
    defparam i1_4_lut_adj_2082.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1444_3_lut (.I0(n2121), 
            .I1(n2188), .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1380_3_lut (.I0(n2025), 
            .I1(n2092_adj_5995), .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2083 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [3]), 
            .O(n58880));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2083.LUT_INIT = 16'h2300;
    SB_LUT4 i54006_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n63074), 
            .O(n2940));
    defparam i54006_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1447_3_lut (.I0(n2124), 
            .I1(n2191), .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2084 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [4]), 
            .O(n58837));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2084.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1931_3_lut (.I0(n2832), 
            .I1(n2899), .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29533_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i29533_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29532_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i29532_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30207_2_lut (.I0(duty[19]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5437));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30207_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2085 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [5]), 
            .O(n58881));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2085.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1514_3_lut (.I0(n2223), 
            .I1(n2290), .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2086 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [6]), 
            .O(n58882));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2086.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2087 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [5]), 
            .O(n58980));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2087.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2088 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [6]), 
            .O(n58979));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2088.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2089 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[22] [7]), 
            .O(n58883));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2089.LUT_INIT = 16'h2300;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n28127), .O(n55126));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1511_3_lut (.I0(n2220), 
            .I1(n2287), .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1578_3_lut (.I0(n2319), 
            .I1(n2386), .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1645_3_lut (.I0(n2418), 
            .I1(n2485), .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1712_3_lut (.I0(n2517), 
            .I1(n2584), .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2090 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[5] [7]), 
            .O(n58978));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2090.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2091 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [2]), 
            .O(n58967));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2091.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2092 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [0]), 
            .O(n58977));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2092.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1581_3_lut (.I0(n2322), 
            .I1(n2389), .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1648_3_lut (.I0(n2421), 
            .I1(n2488), .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1998_3_lut (.I0(n2931), 
            .I1(n2998), .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2093 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [0]), 
            .O(n58884));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2093.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n652));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30206_2_lut (.I0(duty[20]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5436));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30206_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2094 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [3]), 
            .O(n58966));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2094.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2095 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [1]), 
            .O(n58885));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2095.LUT_INIT = 16'h2300;
    SB_LUT4 i15714_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n23230), .I3(GND_net), .O(n30121));   // verilog/coms.v(130[12] 305[6])
    defparam i15714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15716_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n23230), .I3(GND_net), .O(n30123));   // verilog/coms.v(130[12] 305[6])
    defparam i15716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30205_2_lut (.I0(duty[21]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5435));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30205_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15717_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n23230), .I3(GND_net), .O(n30124));   // verilog/coms.v(130[12] 305[6])
    defparam i15717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15718_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n23230), .I3(GND_net), .O(n30125));   // verilog/coms.v(130[12] 305[6])
    defparam i15718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15719_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n23230), .I3(GND_net), .O(n30126));   // verilog/coms.v(130[12] 305[6])
    defparam i15719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2096 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [2]), 
            .O(n58831));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2096.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2097 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [3]), 
            .O(n58830));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2097.LUT_INIT = 16'h2300;
    SB_LUT4 i51645_2_lut_4_lut (.I0(duty[8]), .I1(n338), .I2(duty[4]), 
            .I3(n342), .O(n67819));
    defparam i51645_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2098 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [4]), 
            .O(n58886));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2098.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1715_3_lut (.I0(n2520), 
            .I1(n2587), .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15720_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n23230), .I3(GND_net), .O(n30127));   // verilog/coms.v(130[12] 305[6])
    defparam i15720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15721_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n23230), .I3(GND_net), .O(n30128));   // verilog/coms.v(130[12] 305[6])
    defparam i15721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2099 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [5]), 
            .O(n58887));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2099.LUT_INIT = 16'h2300;
    SB_LUT4 i15722_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n23230), .I3(GND_net), .O(n30129));   // verilog/coms.v(130[12] 305[6])
    defparam i15722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2100 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [6]), 
            .O(n58888));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2100.LUT_INIT = 16'h2300;
    SB_LUT4 i15723_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n23230), .I3(GND_net), .O(n30130));   // verilog/coms.v(130[12] 305[6])
    defparam i15723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53733_2_lut_4_lut (.I0(\data_out_frame[15] [7]), .I1(n54003), 
            .I2(\data_out_frame[13] [7]), .I3(\data_out_frame[16] [1]), 
            .O(n69908));   // verilog/coms.v(100[12:26])
    defparam i53733_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2101 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[23] [7]), 
            .O(n58889));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2101.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2102 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [0]), 
            .O(n58890));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2102.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51594_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n67768));
    defparam i51594_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1779_3_lut (.I0(n2616), 
            .I1(n2683), .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1782_3_lut (.I0(n2619), 
            .I1(n2686), .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5845));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_17_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1849_3_lut (.I0(n2718), 
            .I1(n2785), .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i2_3_lut (.I0(encoder0_position_scaled_23__N_319[1]), 
            .I1(n32_adj_5937), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1846_3_lut (.I0(n2715), 
            .I1(n2782), .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1850_3_lut (.I0(n2719), 
            .I1(n2786), .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1917_3_lut (.I0(n2818), 
            .I1(n2885), .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30204_2_lut (.I0(duty[22]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5434));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30204_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i54517_1_lut_4_lut (.I0(current[15]), .I1(duty[23]), .I2(n61445), 
            .I3(n61440), .O(n70691));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54517_1_lut_4_lut.LUT_INIT = 16'h4c5d;
    SB_LUT4 i1_4_lut_4_lut_adj_2103 (.I0(current[15]), .I1(duty[23]), .I2(n61445), 
            .I3(n61440), .O(n209));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i1_4_lut_4_lut_adj_2103.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2104 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [1]), 
            .O(n58891));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2104.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2105 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [2]), 
            .O(n58892));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2105.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1916_3_lut (.I0(n2817), 
            .I1(n2884), .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i7_3_lut (.I0(encoder0_position_scaled_23__N_319[6]), 
            .I1(n27), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n952));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2106 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [3]), 
            .O(n58893));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2106.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i6_3_lut (.I0(encoder0_position_scaled_23__N_319[5]), 
            .I1(n28), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n953));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2107 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [4]), 
            .O(n58894));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2107.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20577_4_lut_4_lut (.I0(current[1]), .I1(duty[2]), .I2(current[2]), 
            .I3(duty[1]), .O(n4_adj_5907));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i20577_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51568_2_lut_4_lut (.I0(current[7]), .I1(duty[7]), .I2(current[3]), 
            .I3(duty[3]), .O(n67742));
    defparam i51568_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[3]), .I1(duty[7]), .I2(current[7]), 
            .I3(GND_net), .O(n6_adj_5905));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2108 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [5]), 
            .O(n29283));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2108.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2109 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [6]), 
            .O(n58895));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2109.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2110 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[24] [7]), 
            .O(n58824));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2110.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2111 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [0]), 
            .O(n29256));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2111.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1932_3_lut (.I0(n2833), 
            .I1(n2900), .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30228_2_lut (.I0(n356), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5409));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30228_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i5_3_lut (.I0(encoder0_position_scaled_23__N_319[4]), 
            .I1(n29), .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), 
            .O(n954));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i20_3_lut (.I0(encoder0_position_scaled_23__N_319[19]), 
            .I1(n14_adj_5950), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15376_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n78), .I3(GND_net), .O(n29783));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533_adj_5993));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2112 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [1]), 
            .O(n29255));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2112.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1048_3_lut (.I0(n1533_adj_5993), 
            .I1(n1600), .I2(n1554_adj_5994), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2113 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [2]), 
            .O(n29254));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2113.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2114 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [3]), 
            .O(n58896));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2114.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1115_3_lut (.I0(n1632), 
            .I1(n1699), .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2115 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [4]), 
            .O(n29251));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2115.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2116 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [5]), 
            .O(n58897));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2116.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2117 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [6]), 
            .O(n58898));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2117.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_adj_2118 (.I0(n2_adj_5962), .I1(n3_adj_5961), 
            .I2(encoder0_position_scaled_23__N_319[31]), .I3(GND_net), .O(n63466));
    defparam i1_2_lut_3_lut_adj_2118.LUT_INIT = 16'h8080;
    SB_LUT4 i43757_2_lut_3_lut (.I0(n2_adj_5962), .I1(n3_adj_5961), .I2(n5_adj_6069), 
            .I3(GND_net), .O(n59878));
    defparam i43757_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1182_3_lut (.I0(n1731), 
            .I1(n1798), .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1249_3_lut (.I0(n1830), 
            .I1(n1897), .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1316_3_lut (.I0(n1929), 
            .I1(n1996), .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2119 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [7]), 
            .O(n58828));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2119.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1383_3_lut (.I0(n2028), 
            .I1(n2095), .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1450_3_lut (.I0(n2127), 
            .I1(n2194), .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5917));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2120 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [1]), 
            .O(n58976));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2120.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1517_3_lut (.I0(n2226), 
            .I1(n2293), .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1584_3_lut (.I0(n2325), 
            .I1(n2392), .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1651_3_lut (.I0(n2424), 
            .I1(n2491), .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1718_3_lut (.I0(n2523), 
            .I1(n2590), .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1785_3_lut (.I0(n2622), 
            .I1(n2689), .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30469_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n44773));
    defparam i30469_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2121 (.I0(n1324), .I1(n1323), .I2(n1327), .I3(n1328), 
            .O(n60859));
    defparam i1_4_lut_adj_2121.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2122 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [2]), 
            .O(n58975));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2122.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2123 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [3]), 
            .O(n58974));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2123.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2124 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[6] [4]), 
            .O(n58973));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2124.LUT_INIT = 16'h2300;
    SB_LUT4 i15134_2_lut_3_lut (.I0(n23298), .I1(dti), .I2(n15_adj_5909), 
            .I3(GND_net), .O(n29536));
    defparam i15134_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_2_lut_3_lut_adj_2125 (.I0(n23298), .I1(dti), .I2(n15_adj_5909), 
            .I3(GND_net), .O(n28182));
    defparam i1_2_lut_3_lut_adj_2125.LUT_INIT = 16'hf8f8;
    SB_LUT4 i6615_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_513));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6615_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i1_4_lut_adj_2126 (.I0(n1329), .I1(n44773), .I2(n1330), .I3(n1331), 
            .O(n60700));
    defparam i1_4_lut_adj_2126.LUT_INIT = 16'ha080;
    SB_LUT4 i6613_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_504));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6613_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2127 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [4]), 
            .O(n58965));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2127.LUT_INIT = 16'h2300;
    SB_LUT4 i54457_4_lut (.I0(n60700), .I1(n60859), .I2(n1325), .I3(n1326), 
            .O(n1356));
    defparam i54457_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5918));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_mux_3_i21_3_lut (.I0(encoder0_position_scaled_23__N_319[20]), 
            .I1(n13_adj_5951), .I2(encoder0_position_scaled_23__N_319[31]), 
            .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_2128 (.I0(n1428), .I1(n1427), .I2(GND_net), .I3(GND_net), 
            .O(n63350));
    defparam i1_2_lut_adj_2128.LUT_INIT = 16'heeee;
    SB_LUT4 i15426_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n42166), .I3(n8_adj_5843), .O(n29833));   // verilog/coms.v(130[12] 305[6])
    defparam i15426_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2129 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [5]), 
            .O(n59004));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2129.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2130 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_6083));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2130.LUT_INIT = 16'h7bde;
    \quadrature_decoder(1)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n2270(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .b_prev(b_prev_adj_5931), 
            .n30060(n30060), .n2275(n2275), .position_31__N_3956(position_31__N_3956_adj_5932), 
            .encoder1_position({encoder1_position}), .GND_net(GND_net), 
            .\a_new[1] (a_new_adj_6125[1]), .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[49] 318[6])
    TLI4970 tli (.\data[12] (data_adj_6147[12]), .GND_net(GND_net), .clk16MHz(clk16MHz), 
            .n30250(n30250), .\data[15] (data_adj_6147[15]), .n30249(n30249), 
            .n30248(n30248), .\data[11] (data_adj_6147[11]), .n30247(n30247), 
            .\data[10] (data_adj_6147[10]), .n30246(n30246), .\data[9] (data_adj_6147[9]), 
            .n30245(n30245), .\data[8] (data_adj_6147[8]), .n30244(n30244), 
            .\data[7] (data_adj_6147[7]), .n30243(n30243), .\data[6] (data_adj_6147[6]), 
            .n30242(n30242), .\data[5] (data_adj_6147[5]), .n30241(n30241), 
            .\data[4] (data_adj_6147[4]), .n30240(n30240), .\data[3] (data_adj_6147[3]), 
            .n30239(n30239), .\data[2] (data_adj_6147[2]), .n30238(n30238), 
            .\data[1] (data_adj_6147[1]), .\state[0] (state_adj_6149[0]), 
            .n15(n15_adj_5916), .clk_out(clk_out), .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), 
            .VCC_net(VCC_net), .n6(n6_adj_5883), .\state[1] (state_adj_6149[1]), 
            .n9(n9_adj_6085), .n30025(n30025), .n30023(n30023), .\current[0] (current[0]), 
            .n6_adj_26(n6_adj_5915), .n6_adj_27(n6_adj_5914), .state_7__N_4446(state_7__N_4446), 
            .n43986(n43986), .n30855(n30855), .\data[0] (data_adj_6147[0]), 
            .n30759(n30759), .\current[1] (current[1]), .n30758(n30758), 
            .\current[2] (current[2]), .n30757(n30757), .\current[3] (current[3]), 
            .n30756(n30756), .\current[4] (current[4]), .n30755(n30755), 
            .\current[5] (current[5]), .n30754(n30754), .\current[6] (current[6]), 
            .n30753(n30753), .\current[7] (current[7]), .n30752(n30752), 
            .\current[8] (current[8]), .n30751(n30751), .\current[9] (current[9]), 
            .n30750(n30750), .\current[10] (current[10]), .n30749(n30749), 
            .\current[11] (current[11]), .n28109(n28109), .\current[15] (current[15]), 
            .n11(n11_adj_5928), .n25959(n25959), .n25966(n25966), .n25977(n25977), 
            .n25971(n25971)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(416[11] 422[4])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2131 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [6]), 
            .O(n58964));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2131.LUT_INIT = 16'h2300;
    SB_LUT4 i30467_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n44771));
    defparam i30467_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5919));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2136_3_lut (.I0(n3133), 
            .I1(n3200), .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2132 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n63350), 
            .O(n63356));
    defparam i1_4_lut_adj_2132.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2133 (.I0(commutation_state[0]), .I1(n4_adj_6083), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5909));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut_adj_2133.LUT_INIT = 16'hdede;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2134 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[7] [7]), 
            .O(n58963));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2134.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2135 (.I0(n1429), .I1(n44771), .I2(n1430), .I3(n1431), 
            .O(n60713));
    defparam i1_4_lut_adj_2135.LUT_INIT = 16'ha080;
    SB_LUT4 i30210_2_lut (.I0(duty[16]), .I1(n296), .I2(GND_net), .I3(GND_net), 
            .O(n5440));   // verilog/TinyFPGA_B.v(123[17] 125[11])
    defparam i30210_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [5]), .I3(\data_in_frame[16] [7]), .O(n7_adj_6064));   // verilog/coms.v(99[12:25])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_6082));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_2136 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_6081));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_2136.LUT_INIT = 16'hfffe;
    SB_LUT4 i54398_4_lut (.I0(n60713), .I1(n1422), .I2(n1423), .I3(n63356), 
            .O(n1455));
    defparam i54398_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i7_4_lut_adj_2137 (.I0(dti_counter[0]), .I1(n14_adj_6081), .I2(n10_adj_6082), 
            .I3(dti_counter[3]), .O(n23298));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_2137.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30523_4_lut (.I0(n940), .I1(n1531_adj_5991), .I2(n1532_adj_5992), 
            .I3(n1533_adj_5993), .O(n44827));
    defparam i30523_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2138 (.I0(n1525), .I1(n1527), .I2(n1528), .I3(GND_net), 
            .O(n63326));
    defparam i1_3_lut_adj_2138.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2139 (.I0(n1529), .I1(n63326), .I2(n44827), .I3(n1530), 
            .O(n63328));
    defparam i1_4_lut_adj_2139.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_2140 (.I0(n1522), .I1(n1524), .I2(n1526), .I3(GND_net), 
            .O(n63272));
    defparam i1_3_lut_adj_2140.LUT_INIT = 16'hfefe;
    SB_LUT4 i54376_4_lut (.I0(n63272), .I1(n1521), .I2(n63328), .I3(n1523), 
            .O(n1554_adj_5994));
    defparam i54376_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54381_2_lut (.I0(n23298), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_517));
    defparam i54381_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15406_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n59067), .I3(state_7__N_4237[0]), 
            .O(n29813));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15406_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2141 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [0]), 
            .O(n58962));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2141.LUT_INIT = 16'h2300;
    SB_LUT4 i15502_3_lut_4_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n42166), .I3(n8_adj_5973), .O(n29909));   // verilog/coms.v(130[12] 305[6])
    defparam i15502_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15505_3_lut_4_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n42166), .I3(n8_adj_5973), .O(n29912));   // verilog/coms.v(130[12] 305[6])
    defparam i15505_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i1941_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1642), .I3(n43842), .O(n7082));   // verilog/TinyFPGA_B.v(373[5] 399[12])
    defparam i1941_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i15570_3_lut_4_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(reset), .I3(n51), .O(n29977));   // verilog/coms.v(130[12] 305[6])
    defparam i15570_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n51), .I2(GND_net), .I3(GND_net), 
            .O(n28768));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5920));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2135_3_lut (.I0(n3132), 
            .I1(n3199), .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532_adj_5992));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2142 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [1]), 
            .O(n58961));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2142.LUT_INIT = 16'h2300;
    SB_LUT4 mux_282_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i1_3_lut (.I0(encoder0_position_scaled[0]), .I1(motor_state_23__N_115[0]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5921));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_4_lut_adj_2143 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_522), .I3(n3305), .O(n25_adj_6071));   // verilog/TinyFPGA_B.v(388[7:11])
    defparam i1_4_lut_4_lut_adj_2143.LUT_INIT = 16'h5450;
    SB_LUT4 i1_3_lut_adj_2144 (.I0(n1627), .I1(n1628), .I2(n1626), .I3(GND_net), 
            .O(n63422));
    defparam i1_3_lut_adj_2144.LUT_INIT = 16'hfefe;
    SB_LUT4 i51791_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n40932), 
            .I2(start), .I3(state[0]), .O(n67080));   // verilog/neopixel.v(34[12] 116[6])
    defparam i51791_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2145 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[8] [2]), 
            .O(n58960));   // verilog/TinyFPGA_B.v(370[10] 400[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2145.LUT_INIT = 16'h2300;
    SB_LUT4 i30519_4_lut (.I0(n941), .I1(n1631), .I2(n1632), .I3(n1633), 
            .O(n44823));
    defparam i30519_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2146 (.I0(n1623), .I1(n1624), .I2(n63422), .I3(n1625), 
            .O(n63428));
    defparam i1_4_lut_adj_2146.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2147 (.I0(n1629), .I1(n63428), .I2(n44823), .I3(n1630), 
            .O(n63430));
    defparam i1_4_lut_adj_2147.LUT_INIT = 16'heccc;
    SB_LUT4 i10_1_lut_adj_2148 (.I0(duty[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_setpoint_23__N_255));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i10_1_lut_adj_2148.LUT_INIT = 16'h5555;
    SB_LUT4 i54355_4_lut (.I0(n1621), .I1(n1620), .I2(n63430), .I3(n1622), 
            .O(n1653));
    defparam i54355_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1047_3_lut (.I0(n1532_adj_5992), 
            .I1(n1599), .I2(n1554_adj_5994), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2149 (.I0(n1728), .I1(n1727), .I2(GND_net), .I3(GND_net), 
            .O(n63000));
    defparam i1_2_lut_adj_2149.LUT_INIT = 16'heeee;
    SB_LUT4 i30451_3_lut (.I0(n942), .I1(n1732), .I2(n1733), .I3(GND_net), 
            .O(n44755));
    defparam i30451_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_2150 (.I0(n1724), .I1(n1725), .I2(n63000), .I3(n1726), 
            .O(n63006));
    defparam i1_4_lut_adj_2150.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2151 (.I0(n1729), .I1(n44755), .I2(n1730), .I3(n1731), 
            .O(n60718));
    defparam i1_4_lut_adj_2151.LUT_INIT = 16'ha080;
    SB_LUT4 i48278_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64452));
    defparam i48278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48279_4_lut (.I0(n64452), .I1(n28507), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1] [0]), .O(n64453));
    defparam i48279_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i48277_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64451));
    defparam i48277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2152 (.I0(n1722), .I1(n1723), .I2(n60718), .I3(n63006), 
            .O(n63012));
    defparam i1_4_lut_adj_2152.LUT_INIT = 16'hfffe;
    SB_LUT4 i54333_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n63012), 
            .O(n1752));
    defparam i54333_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i29534_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i29534_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1114_3_lut (.I0(n1631), 
            .I1(n1698), .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2153 (.I0(n1827), .I1(n1826), .I2(n1825), .I3(n1828), 
            .O(n63440));
    defparam i1_4_lut_adj_2153.LUT_INIT = 16'hfffe;
    SB_LUT4 i30473_4_lut (.I0(n943), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n44777));
    defparam i30473_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2154 (.I0(n1822), .I1(n1823), .I2(n63440), .I3(n1824), 
            .O(n63446));
    defparam i1_4_lut_adj_2154.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2155 (.I0(n1829), .I1(n1830), .I2(GND_net), .I3(GND_net), 
            .O(n63470));
    defparam i1_2_lut_adj_2155.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5922));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2156 (.I0(n63470), .I1(n1821), .I2(n63446), .I3(n44777), 
            .O(n63450));
    defparam i1_4_lut_adj_2156.LUT_INIT = 16'hfefc;
    coms neopxl_color_23__I_0 (.VCC_net(VCC_net), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .clk16MHz(clk16MHz), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[1] ({\data_in_frame[1] [7:2], Open_0, Open_1}), 
         .n3358(n3358), .\data_out_frame[6] ({\data_out_frame[6] }), .n58972(n58972), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .IntegralLimit({IntegralLimit}), 
         .n58971(n58971), .GND_net(GND_net), .\data_in_frame[0] ({\data_in_frame[0] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\FRAME_MATCHER.i_31__N_2638 (\FRAME_MATCHER.i_31__N_2638 ), 
         .control_mode({control_mode}), .n58970(n58970), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .n58969(n58969), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .displacement({displacement}), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .ID({ID}), .\data_in_frame[16] ({\data_in_frame[16] [7], Open_2, 
         Open_3, Open_4, Open_5, Open_6, Open_7, Open_8}), .deadband({deadband}), 
         .byte_transmit_counter({Open_9, Open_10, Open_11, Open_12, 
         Open_13, Open_14, Open_15, byte_transmit_counter[0]}), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\byte_transmit_counter[1] (byte_transmit_counter[1]), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n28(n28_adj_6009), .n379(n379_adj_5927), .n405(n405), .n4(n4_adj_6000), 
         .encoder0_position_scaled({encoder0_position_scaled}), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), 
         .n8(n8_adj_5908), .\data_in_frame[14] ({\data_in_frame[14] }), 
         .n58968(n58968), .n58967(n58967), .n58966(n58966), .n58965(n58965), 
         .n59004(n59004), .n58964(n58964), .reset(reset), .setpoint({setpoint}), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n58963(n58963), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .n58962(n58962), .n58961(n58961), 
         .n58960(n58960), .n58959(n58959), .n58958(n58958), .n58957(n58957), 
         .n58825(n58825), .n58956(n58956), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .n58955(n58955), .n58954(n58954), .n58953(n58953), .n58952(n58952), 
         .n58951(n58951), .n30260(n30260), .n30257(n30257), .n149(n149), 
         .n11(n11_adj_5999), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .n70864(n70864), 
         .\data_out_frame[1][7] (\data_out_frame[1] [7]), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n28507(n28507), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n58950(n58950), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .n58949(n58949), 
         .n58948(n58948), .n58947(n58947), .n58946(n58946), .n58945(n58945), 
         .n58944(n58944), .n58943(n58943), .n58942(n58942), .n58941(n58941), 
         .n58940(n58940), .n60(n60), .n51(n51), .n58939(n58939), .n58938(n58938), 
         .n58937(n58937), .n58936(n58936), .n28717(n28717), .n28774(n28774), 
         .rx_data({rx_data}), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n30228(n30228), .n30225(n30225), .n58935(n58935), .n30222(n30222), 
         .n30219(n30219), .n30216(n30216), .n30208(n30208), .n30207(n30207), 
         .neopxl_color({neopxl_color}), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .\data_in_frame[20][7] (\data_in_frame[20] [7]), 
         .\data_in_frame[17] ({Open_16, Open_17, \data_in_frame[17] [5:1], 
         Open_18}), .\data_in_frame[20][1] (\data_in_frame[20] [1]), .\data_in_frame[20][5] (\data_in_frame[20] [5]), 
         .\data_in_frame[8] ({Open_19, \data_in_frame[8] [6], Open_20, 
         Open_21, Open_22, Open_23, Open_24, Open_25}), .n25605(n25605), 
         .n59499(n59499), .n61411(n61411), .encoder1_position_scaled({encoder1_position_scaled}), 
         .\data_in_frame[6] ({Open_26, Open_27, Open_28, Open_29, Open_30, 
         Open_31, Open_32, \data_in_frame[6] [0]}), .\motor_state_23__N_115[13] (motor_state_23__N_115[13]), 
         .n15(n15_adj_5929), .n10(n10), .n58934(n58934), .n58933(n58933), 
         .n58932(n58932), .n58931(n58931), .n58930(n58930), .n58929(n58929), 
         .n58928(n58928), .n58927(n58927), .n58926(n58926), .\Kp[1] (Kp[1]), 
         .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .n58925(n58925), .\Kp[4] (Kp[4]), 
         .n58924(n58924), .n58826(n58826), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
         .\Kp[7] (Kp[7]), .n58923(n58923), .n58922(n58922), .n58921(n58921), 
         .\Kp[8] (Kp[8]), .n58920(n58920), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
         .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .n58919(n58919), .n58918(n58918), 
         .n58917(n58917), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), 
         .n58916(n58916), .n58915(n58915), .\Ki[1] (Ki[1]), .n58914(n58914), 
         .n58913(n58913), .n58912(n58912), .\Ki[2] (Ki[2]), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
         .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
         .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .n26902(n26902), 
         .n58911(n58911), .n58910(n58910), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
         .n30130(n30130), .current_limit({current_limit}), .n30129(n30129), 
         .n30128(n30128), .n30127(n30127), .n58909(n58909), .n58908(n58908), 
         .n58907(n58907), .n58906(n58906), .n30126(n30126), .n30125(n30125), 
         .n30124(n30124), .n30123(n30123), .n30121(n30121), .PWMLimit({PWMLimit}), 
         .n58905(n58905), .n58904(n58904), .n58903(n58903), .n58902(n58902), 
         .n58901(n58901), .\data_in_frame[20][0] (\data_in_frame[20] [0]), 
         .n59138(n59138), .n30090(n30090), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n59971(n59971), .n30075(n30075), .n30074(n30074), .n59994(n59994), 
         .\data_in_frame[8][7] (\data_in_frame[8] [7]), .n58900(n58900), 
         .n28801(n28801), .\data_in_frame[6][2] (\data_in_frame[6] [2]), 
         .n30073(n30073), .n30072(n30072), .n30068(n30068), .n30067(n30067), 
         .n30066(n30066), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n30062(n30062), .n30061(n30061), .n30059(n30059), .n30057(n30057), 
         .n30010(n30010), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n58899(n58899), 
         .n58829(n58829), .n58832(n58832), .n58833(n58833), .n58834(n58834), 
         .n58835(n58835), .n58836(n58836), .n58841(n58841), .n58843(n58843), 
         .n58847(n58847), .n58848(n58848), .n58849(n58849), .n58850(n58850), 
         .n58844(n58844), .n58851(n58851), .n58852(n58852), .n58846(n58846), 
         .n58853(n58853), .n58854(n58854), .n58855(n58855), .n58856(n58856), 
         .n58857(n58857), .n58858(n58858), .n58859(n58859), .n58827(n58827), 
         .\data_in_frame[17][7] (\data_in_frame[17] [7]), .\data_in_frame[17][6] (\data_in_frame[17] [6]), 
         .n58860(n58860), .n58861(n58861), .n58862(n58862), .n58863(n58863), 
         .n58864(n58864), .DE_c(DE_c), .tx_active(tx_active), .LED_c(LED_c), 
         .n58845(n58845), .n59003(n59003), .n58865(n58865), .\data_in_frame[7][7] (\data_in_frame[7] [7]), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n59002(n59002), .\data_in_frame[7][2] (\data_in_frame[7] [2]), 
         .\data_in_frame[6][7] (\data_in_frame[6] [7]), .n58866(n58866), 
         .\data_out_frame[1][0] (\data_out_frame[1] [0]), .n59001(n59001), 
         .n28780(n28780), .\data_in_frame[7][0] (\data_in_frame[7] [0]), 
         .\data_out_frame[1][1] (\data_out_frame[1] [1]), .n59000(n59000), 
         .n58999(n58999), .n31074(n31074), .n29319(n29319), .n31075(n31075), 
         .n29318(n29318), .n58998(n58998), .\data_in_frame[8][4] (\data_in_frame[8] [4]), 
         .\data_in_frame[7][4] (\data_in_frame[7] [4]), .\data_in_frame[8][5] (\data_in_frame[8] [5]), 
         .\data_in_frame[6][3] (\data_in_frame[6] [3]), .\data_in_frame[7][3] (\data_in_frame[7] [3]), 
         .\data_in_frame[7][5] (\data_in_frame[7] [5]), .n30842(n30842), 
         .n30828(n30828), .n23230(n23230), .n30773(n30773), .n30763(n30763), 
         .n30761(n30761), .n30760(n30760), .n30744(n30744), .n30742(n30742), 
         .\data_in_frame[6][1] (\data_in_frame[6] [1]), .n30710(n30710), 
         .n30707(n30707), .n30706(n30706), .n30705(n30705), .n30703(n30703), 
         .n30702(n30702), .n58296(n58296), .n29833(n29833), .n30693(n30693), 
         .n30690(n30690), .n58294(n58294), .n58290(n58290), .n58286(n58286), 
         .n58282(n58282), .n58278(n58278), .n58274(n58274), .n58272(n58272), 
         .n58268(n58268), .n29861(n29861), .n58264(n58264), .n29867(n29867), 
         .n58260(n58260), .n30677(n30677), .n30674(n30674), .n58256(n58256), 
         .n30672(n30672), .n30669(n30669), .n30664(n30664), .n30338(n30338), 
         .n30342(n30342), .n30348(n30348), .n30352(n30352), .\data_in_frame[6][4] (\data_in_frame[6] [4]), 
         .n30361(n30361), .n30365(n30365), .n30368(n30368), .\data_in_frame[7][1] (\data_in_frame[7] [1]), 
         .n30371(n30371), .n30375(n30375), .n30378(n30378), .n30381(n30381), 
         .n30387(n30387), .n30399(n30399), .\data_in_frame[8][3] (\data_in_frame[8] [3]), 
         .n30403(n30403), .n30639(n30639), .n30638(n30638), .n30406(n30406), 
         .n30409(n30409), .n30413(n30413), .n30466(n30466), .n30469(n30469), 
         .n30616(n30616), .n30475(n30475), .n30479(n30479), .n30482(n30482), 
         .n30485(n30485), .n30489(n30489), .n30492(n30492), .n30495(n30495), 
         .n30499(n30499), .n58384(n58384), .n58398(n58398), .n30509(n30509), 
         .n30512(n30512), .n30515(n30515), .n30550(n30550), .n30554(n30554), 
         .n30558(n30558), .n30562(n30562), .n30566(n30566), .n30587(n30587), 
         .n58252(n58252), .n58248(n58248), .n58244(n58244), .\data_in_frame[20][2] (\data_in_frame[20] [2]), 
         .n29909(n29909), .\data_in_frame[20][3] (\data_in_frame[20] [3]), 
         .n29912(n29912), .\data_in_frame[20][4] (\data_in_frame[20] [4]), 
         .n58238(n58238), .n58234(n58234), .n58230(n58230), .n58228(n58228), 
         .n58226(n58226), .n58224(n58224), .n58220(n58220), .n58216(n58216), 
         .n58212(n58212), .n58208(n58208), .n29949(n29949), .\data_in_frame[22] ({\data_in_frame[22] }), 
         .n29952(n29952), .n58202(n58202), .n29958(n29958), .n29961(n29961), 
         .n29964(n29964), .n29968(n29968), .n58198(n58198), .n30539(n30539), 
         .n29977(n29977), .\data_in_frame[23] ({\data_in_frame[23] }), .n29980(n29980), 
         .n29983(n29983), .n29986(n29986), .n29989(n29989), .n29992(n29992), 
         .n29995(n29995), .n30465(n30465), .n30003(n30003), .n30016(n30016), 
         .n30028(n30028), .n30031(n30031), .n30035(n30035), .n58340(n58340), 
         .n58997(n58997), .n58996(n58996), .n58995(n58995), .n58994(n58994), 
         .n58842(n58842), .n31082(n31082), .n29317(n29317), .n58993(n58993), 
         .n58992(n58992), .n58991(n58991), .n58990(n58990), .\data_in_frame[1][1] (\data_in_frame[1] [1]), 
         .n58989(n58989), .n58988(n58988), .rx_data_ready(rx_data_ready), 
         .n59967(n59967), .n58867(n58867), .n58868(n58868), .n58987(n58987), 
         .n58986(n58986), .n58985(n58985), .n58984(n58984), .n58869(n58869), 
         .n58840(n58840), .n58839(n58839), .n58983(n58983), .n58982(n58982), 
         .n58981(n58981), .n58870(n58870), .n42166(n42166), .n28770(n28770), 
         .n58871(n58871), .n59086(n59086), .n29311(n29311), .n58872(n58872), 
         .n58873(n58873), .n58874(n58874), .n58875(n58875), .n58876(n58876), 
         .n58877(n58877), .n58878(n58878), .n8_adj_10(n8_adj_5843), .n28725(n28725), 
         .n58879(n58879), .n58838(n58838), .n58880(n58880), .n58837(n58837), 
         .n58881(n58881), .n58882(n58882), .n8_adj_11(n8_adj_5973), .n8_adj_12(n8_adj_5936), 
         .n28733(n28733), .n58980(n58980), .n58979(n58979), .n58883(n58883), 
         .n58978(n58978), .n58977(n58977), .n58884(n58884), .n58885(n58885), 
         .n58831(n58831), .n58830(n58830), .n58886(n58886), .n58887(n58887), 
         .n58888(n58888), .n58889(n58889), .n58890(n58890), .n58891(n58891), 
         .n58892(n58892), .n58893(n58893), .n58894(n58894), .n29283(n29283), 
         .\data_out_frame[27][6] (\data_out_frame[27] [6]), .\data_out_frame[26][6] (\data_out_frame[26] [6]), 
         .n58895(n58895), .n58824(n58824), .n31162(n31162), .n29256(n29256), 
         .n31163(n31163), .n29255(n29255), .n31164(n31164), .n29254(n29254), 
         .n58896(n58896), .n31166(n31166), .n29251(n29251), .n58897(n58897), 
         .n58898(n58898), .n58828(n58828), .n58976(n58976), .n59079(n59079), 
         .n58975(n58975), .n58974(n58974), .n58973(n58973), .n69908(n69908), 
         .n28778(n28778), .n69906(n69906), .n26087(n26087), .n59593(n59593), 
         .n26490(n26490), .n54003(n54003), .pwm_setpoint({pwm_setpoint}), 
         .n23164(n23164), .n44625(n44625), .n64453(n64453), .n64451(n64451), 
         .n59093(n59093), .n28719(n28719), .n28723(n28723), .n35592(n35592), 
         .n15_adj_13(n15_adj_5933), .n54986(n54986), .n59975(n59975), 
         .n28791(n28791), .\current[7] (current[7]), .\current[6] (current[6]), 
         .\current[5] (current[5]), .\current[4] (current[4]), .\current[3] (current[3]), 
         .\current[2] (current[2]), .\current[1] (current[1]), .\current[0] (current[0]), 
         .\current[15] (current[15]), .\current[11] (current[11]), .\current[10] (current[10]), 
         .\current[9] (current[9]), .\current[8] (current[8]), .\o_Rx_DV_N_3617[24] (o_Rx_DV_N_3617[24]), 
         .r_SM_Main({r_SM_Main_adj_6161}), .n27(n27_adj_5989), .n62584(n62584), 
         .n28320(n28320), .n60079(n60079), .n1(n1), .tx_o(tx_o), .r_Clock_Count({r_Clock_Count_adj_6162}), 
         .n30034(n30034), .n71131(n71131), .n30847(n30847), .\r_Bit_Index[0] (r_Bit_Index_adj_6163[0]), 
         .n6(n6_adj_6068), .tx_enable(tx_enable), .\o_Rx_DV_N_3617[12] (o_Rx_DV_N_3617[12]), 
         .n5254(n5254), .\o_Rx_DV_N_3617[8] (o_Rx_DV_N_3617[8]), .r_Rx_Data(r_Rx_Data), 
         .n29(n29_adj_5988), .n23(n23_adj_5990), .\r_SM_Main[1]_adj_14 (r_SM_Main[1]), 
         .baudrate({baudrate}), .n28324(n28324), .n60053(n60053), .\r_SM_Main[2]_adj_15 (r_SM_Main[2]), 
         .RX_N_2(RX_N_2), .r_Clock_Count_adj_25({r_Clock_Count}), .n30256(n30256), 
         .n30255(n30255), .n30254(n30254), .n30253(n30253), .n30252(n30252), 
         .n25975(n25975), .\o_Rx_DV_N_3617[7] (o_Rx_DV_N_3617[7]), .\o_Rx_DV_N_3617[6] (o_Rx_DV_N_3617[6]), 
         .\o_Rx_DV_N_3617[5] (o_Rx_DV_N_3617[5]), .\o_Rx_DV_N_3617[4] (o_Rx_DV_N_3617[4]), 
         .\o_Rx_DV_N_3617[3] (o_Rx_DV_N_3617[3]), .\o_Rx_DV_N_3617[2] (o_Rx_DV_N_3617[2]), 
         .\o_Rx_DV_N_3617[1] (o_Rx_DV_N_3617[1]), .\o_Rx_DV_N_3617[0] (o_Rx_DV_N_3617[0]), 
         .\r_Bit_Index[0]_adj_24 (r_Bit_Index[0]), .n62864(n62864), .n29921(n29921), 
         .n59011(n59011), .n62764(n62764), .n62780(n62780), .n62748(n62748), 
         .n62828(n62828), .n62812(n62812), .n30854(n30854), .n55126(n55126), 
         .n30850(n30850), .n5257(n5257), .n29791(n29791), .n28127(n28127), 
         .n62796(n62796), .n62846(n62846)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i54139_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n63450), 
            .O(n1851));
    defparam i54139_4_lut.LUT_INIT = 16'h0001;
    EEPROM eeprom (.enable_slow_N_4340(enable_slow_N_4340), .ready_prev(ready_prev), 
           .clk16MHz(clk16MHz), .n6195({n6196}), .\state[2] (state_adj_6139[2]), 
           .GND_net(GND_net), .n30024(n30024), .rw(rw), .n58524(n58524), 
           .data_ready(data_ready), .n30015(n30015), .ID({ID}), .\state[0] (state_adj_6139[0]), 
           .\state[1] (state_adj_6139[1]), .n58352(n58352), .n30804(n30804), 
           .n30803(n30803), .n30802(n30802), .n30801(n30801), .n30800(n30800), 
           .n30799(n30799), .n30798(n30798), .n30797(n30797), .baudrate({baudrate}), 
           .n30796(n30796), .n30795(n30795), .n30794(n30794), .n30793(n30793), 
           .n30792(n30792), .n30791(n30791), .n30790(n30790), .n30772(n30772), 
           .n30771(n30771), .n30770(n30770), .n30769(n30769), .n30768(n30768), 
           .n30767(n30767), .n30766(n30766), .n30765(n30765), .n3(n3_adj_6054), 
           .n6878(n6878), .n11(n11_adj_5913), .\state[2]_adj_5 (state_adj_6170[2]), 
           .\state[3] (state_adj_6170[3]), .n6(n6_adj_6075), .\state_7__N_4253[3] (state_7__N_4253[3]), 
           .\state_7__N_4045[0] (state_7__N_4045[0]), .\state[1]_adj_6 (state_adj_6170[1]), 
           .\state[0]_adj_7 (state_adj_6170[0]), .n59067(n59067), .n61238(n61238), 
           .n59065(n59065), .n5(n5_adj_6076), .n25956(n25956), .data({data_adj_6138}), 
           .n4(n4_adj_5911), .n49984(n49984), .n62253(n62253), .VCC_net(VCC_net), 
           .sda_enable(sda_enable), .sda_out(sda_out), .scl_enable(scl_enable), 
           .n62(n62), .\state_7__N_4237[0] (state_7__N_4237[0]), .\saved_addr[0] (saved_addr[0]), 
           .n30054(n30054), .n30049(n30049), .n30047(n30047), .n30042(n30042), 
           .n30041(n30041), .n11_adj_8(n11_adj_5912), .n30841(n30841), 
           .n8(n8_adj_6087), .n29813(n29813), .n10(n10_adj_6065), .n4_adj_9(n4_adj_5910), 
           .n44006(n44006), .n25984(n25984), .scl(scl)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(402[10] 414[6])
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i1181_3_lut (.I0(n1730), 
            .I1(n1797), .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5923));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30475_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n44779));
    defparam i30475_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_277_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_115[1]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5924));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20583_3_lut (.I0(current[0]), .I1(n2092), .I2(n209), .I3(GND_net), 
            .O(n270));
    defparam i20583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5925));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_228_i2134_3_lut (.I0(n3131), 
            .I1(n3198), .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(324[33:71])
    defparam encoder0_position_scaled_23__I_0_228_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_282_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_115[2]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5926));   // verilog/TinyFPGA_B.v(326[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_282_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5933), .I3(n61039), .O(motor_state_23__N_115[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_282_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_277_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_115[3]), 
            .I2(n15_adj_5929), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_277_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16675_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[20] [3]), 
            .O(n31082));   // verilog/coms.v(130[12] 305[6])
    defparam i16675_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16759_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [4]), 
            .O(n31166));   // verilog/coms.v(130[12] 305[6])
    defparam i16759_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16757_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [2]), 
            .O(n31164));   // verilog/coms.v(130[12] 305[6])
    defparam i16757_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16756_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[25] [1]), 
            .O(n31163));   // verilog/coms.v(130[12] 305[6])
    defparam i16756_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    motorControl control (.\Ki[14] (Ki[14]), .\PID_CONTROLLER.integral_23__N_3844[1] (\PID_CONTROLLER.integral_23__N_3844 [1]), 
            .GND_net(GND_net), .\Ki[15] (Ki[15]), .\Ki[6] (Ki[6]), .\PID_CONTROLLER.integral_23__N_3844[7] (\PID_CONTROLLER.integral_23__N_3844 [7]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Kp[11] (Kp[11]), 
            .\Ki[10] (Ki[10]), .\Ki[1] (Ki[1]), .\PID_CONTROLLER.integral_23__N_3844[0] (\PID_CONTROLLER.integral_23__N_3844 [0]), 
            .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[11] (Ki[11]), .\Ki[3] (Ki[3]), 
            .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Kp[12] (Kp[12]), .\Ki[4] (Ki[4]), 
            .\Kp[13] (Kp[13]), .\Ki[5] (Ki[5]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .deadband({deadband}), .\Kp[6] (Kp[6]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .n379(n379_adj_5927), .\PID_CONTROLLER.integral_23__N_3844[6] (\PID_CONTROLLER.integral_23__N_3844 [6]), 
            .n4(n4_adj_6000), .control_update(control_update), .\PID_CONTROLLER.integral_23__N_3844[5] (\PID_CONTROLLER.integral_23__N_3844 [5]), 
            .n181(n181), .IntegralLimit({IntegralLimit}), .n155(n155), 
            .\PID_CONTROLLER.integral_23__N_3844[15] (\PID_CONTROLLER.integral_23__N_3844 [15]), 
            .\PID_CONTROLLER.integral_23__N_3844[14] (\PID_CONTROLLER.integral_23__N_3844 [14]), 
            .clk16MHz(clk16MHz), .\PID_CONTROLLER.integral_23__N_3844[16] (\PID_CONTROLLER.integral_23__N_3844 [16]), 
            .VCC_net(VCC_net), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .\Kp[9] (Kp[9]), .\PID_CONTROLLER.integral_23__N_3844[4] (\PID_CONTROLLER.integral_23__N_3844 [4]), 
            .PWMLimit({PWMLimit}), .duty({duty}), .reset(reset), .n149(n149), 
            .n136(n136), .\PID_CONTROLLER.integral_23__N_3844[22] (\PID_CONTROLLER.integral_23__N_3844 [22]), 
            .\PID_CONTROLLER.integral_23__N_3844[21] (\PID_CONTROLLER.integral_23__N_3844 [21]), 
            .n11(n11_adj_5999), .\PID_CONTROLLER.integral_23__N_3844[3] (\PID_CONTROLLER.integral_23__N_3844 [3]), 
            .\Kp[10] (Kp[10]), .\PID_CONTROLLER.integral_23__N_3844[20] (\PID_CONTROLLER.integral_23__N_3844 [20]), 
            .setpoint({setpoint}), .\motor_state[23] (motor_state[23]), 
            .\PID_CONTROLLER.integral_23__N_3844[19] (\PID_CONTROLLER.integral_23__N_3844 [19]), 
            .\PID_CONTROLLER.integral_23__N_3844[17] (\PID_CONTROLLER.integral_23__N_3844 [17]), 
            .n6(n6_adj_6052), .n37023(n37023), .\PID_CONTROLLER.integral_23__N_3844[13] (\PID_CONTROLLER.integral_23__N_3844 [13]), 
            .\motor_state[22] (motor_state[22]), .\PID_CONTROLLER.integral_23__N_3844[23] (\PID_CONTROLLER.integral_23__N_3844 [23]), 
            .n20625(n20625), .n37(n37), .n20626(n20626), .\motor_state[21] (motor_state[21]), 
            .\PID_CONTROLLER.integral_23__N_3844[12] (\PID_CONTROLLER.integral_23__N_3844 [12]), 
            .n188(n188), .\motor_state[20] (motor_state[20]), .\PID_CONTROLLER.integral_23__N_3844[11] (\PID_CONTROLLER.integral_23__N_3844 [11]), 
            .\motor_state[19] (motor_state[19]), .\motor_state[18] (motor_state[18]), 
            .\motor_state[17] (motor_state[17]), .\PID_CONTROLLER.integral_23__N_3844[2] (\PID_CONTROLLER.integral_23__N_3844 [2]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .n10(n10), .\motor_state[12] (motor_state[12]), 
            .n51273(n51273), .\motor_state[11] (motor_state[11]), .\motor_state[10] (motor_state[10]), 
            .\motor_state[9] (motor_state[9]), .\motor_state[8] (motor_state[8]), 
            .\motor_state[7] (motor_state[7]), .\motor_state[6] (motor_state[6]), 
            .\motor_state[5] (motor_state[5]), .\PID_CONTROLLER.integral_23__N_3844[10] (\PID_CONTROLLER.integral_23__N_3844 [10]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .\motor_state[1] (motor_state[1]), 
            .n34987(n34987), .\motor_state[0] (motor_state[0]), .\PID_CONTROLLER.integral_23__N_3844[9] (\PID_CONTROLLER.integral_23__N_3844 [9]), 
            .\PID_CONTROLLER.integral_23__N_3844[8] (\PID_CONTROLLER.integral_23__N_3844 [8]), 
            .n30012(n30012), .n30827(n30827), .n30826(n30826), .n30825(n30825), 
            .n30824(n30824), .n30823(n30823), .n30822(n30822), .n30821(n30821), 
            .n30820(n30820), .n30819(n30819), .n30818(n30818), .n30817(n30817), 
            .n30816(n30816), .n30815(n30815), .n30814(n30814), .n30813(n30813), 
            .n30812(n30812), .n30811(n30811), .n30810(n30810), .n30809(n30809), 
            .n30808(n30808), .n30807(n30807), .n30806(n30806), .n30805(n30805), 
            .n219(n219), .n405(n405), .n38(n38), .n28(n28_adj_6009), 
            .n110(n110), .n20576(n20576), .n20577(n20577), .n56(n56)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    pwm PWM (.GND_net(GND_net), .n3358(n3358), .pwm_out(pwm_out), .clk32MHz(clk32MHz), 
        .VCC_net(VCC_net), .reset(reset), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (n29783, \neo_pixel_transmitter.t0 , 
            clk16MHz, \neo_pixel_transmitter.done , GND_net, n40932, 
            neopxl_color, timer, n30237, n30236, n30235, n30234, 
            n30233, n30232, VCC_net, n30231, \state[0] , \state[1] , 
            n43, n30014, n30013, n57856, start, n29784, NEOPXL_c, 
            LED_c, n78) /* synthesis syn_module_defined=1 */ ;
    input n29783;
    output [10:0]\neo_pixel_transmitter.t0 ;
    input clk16MHz;
    output \neo_pixel_transmitter.done ;
    input GND_net;
    output n40932;
    input [23:0]neopxl_color;
    output [10:0]timer;
    input n30237;
    input n30236;
    input n30235;
    input n30234;
    input n30233;
    input n30232;
    input VCC_net;
    input n30231;
    output \state[0] ;
    output \state[1] ;
    output n43;
    input n30014;
    input n30013;
    input n57856;
    output start;
    input n29784;
    output NEOPXL_c;
    input LED_c;
    output n78;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire \neo_pixel_transmitter.done_N_645 , n59025;
    wire [10:0]n1;
    wire [10:0]one_wire_N_609;
    
    wire n40933;
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    
    wire n64544, n64545, n64566, n64565;
    wire [10:0]n49;
    
    wire n52641, n52640, n52639, n52638, n52637, n52636, n52635, 
        n52634, n52633, n52632, n19, n4, n68686, n67085, n35229, 
        n60065, n68687, n60097, \neo_pixel_transmitter.done_N_651 , 
        n67077, n59983, n29225, n25, n7_adj_5835, n64497, n64496, 
        n70804, n53961, n53940, n64498;
    wire [5:0]color_bit_N_631;
    
    wire n64500, n51422, n51421, n70708, n70702, n64499, n70696, 
        n64501, n57_adj_5836, n65606;
    wire [3:0]state_3__N_560;
    
    wire n51420, n57810, n51419, n35244, n35253;
    wire [4:0]n13;
    
    wire n51418, n70693, n70699, n70705, n51417, n62274, n51416, 
        n51415, n51414, n4_adj_5838, n51413, n44641, n44751, n51094, 
        n59023, n8_adj_5839, n38, n12_adj_5840, n8_adj_5841, n67074, 
        n93, n64189, n64077, n70801;
    
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n29783));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n59025), .D(\neo_pixel_transmitter.done_N_645 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut (.I0(one_wire_N_609[10]), .I1(one_wire_N_609[9]), .I2(one_wire_N_609[8]), 
            .I3(GND_net), .O(n40932));   // verilog/neopixel.v(52[15:25])
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(n40932), .I2(GND_net), 
            .I3(GND_net), .O(n40933));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48370_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64544));
    defparam i48370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48371_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64545));
    defparam i48371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48392_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64566));
    defparam i48392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48391_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64565));
    defparam i48391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2048_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n52641), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2048_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n52640), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n30237));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2048_add_4_11 (.CI(n52640), .I0(GND_net), .I1(timer[9]), 
            .CO(n52641));
    SB_LUT4 timer_2048_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n52639), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_10 (.CI(n52639), .I0(GND_net), .I1(timer[8]), 
            .CO(n52640));
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n30236));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 timer_2048_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n52638), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n30235));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n30234));   // verilog/neopixel.v(34[12] 116[6])
    SB_CARRY timer_2048_add_4_9 (.CI(n52638), .I0(GND_net), .I1(timer[7]), 
            .CO(n52639));
    SB_LUT4 timer_2048_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n52637), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_8 (.CI(n52637), .I0(GND_net), .I1(timer[6]), 
            .CO(n52638));
    SB_LUT4 timer_2048_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n52636), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_7 (.CI(n52636), .I0(GND_net), .I1(timer[5]), 
            .CO(n52637));
    SB_LUT4 timer_2048_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n52635), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_6 (.CI(n52635), .I0(GND_net), .I1(timer[4]), 
            .CO(n52636));
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n30233));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 timer_2048_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n52634), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_5 (.CI(n52634), .I0(GND_net), .I1(timer[3]), 
            .CO(n52635));
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n30232));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 timer_2048_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n52633), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_4 (.CI(n52633), .I0(GND_net), .I1(timer[2]), 
            .CO(n52634));
    SB_LUT4 timer_2048_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n52632), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_3 (.CI(n52632), .I0(GND_net), .I1(timer[1]), 
            .CO(n52633));
    SB_LUT4 timer_2048_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2048_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2048_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n52632));
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n30231));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i52893_4_lut (.I0(n19), .I1(n4), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n68686));
    defparam i52893_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i52_4_lut (.I0(n67085), .I1(n40932), .I2(\state[1] ), .I3(n35229), 
            .O(n60065));
    defparam i52_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i51_4_lut (.I0(n60065), .I1(n68687), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n60097));
    defparam i51_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i47_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_651 ));
    defparam i47_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut (.I0(n67077), .I1(n59983), .I2(\neo_pixel_transmitter.done ), 
            .I3(n43), .O(n29225));   // verilog/neopixel.v(16[11:16])
    defparam i13_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n40933), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n7_adj_5835));
    defparam i15_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i48323_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64497));
    defparam i48323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48322_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64496));
    defparam i48322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48324_4_lut (.I0(n64497), .I1(n70804), .I2(n53961), .I3(n53940), 
            .O(n64498));
    defparam i48324_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48326_4_lut (.I0(n64498), .I1(n64496), .I2(n53961), .I3(color_bit_N_631[1]), 
            .O(n64500));
    defparam i48326_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n51422), .O(one_wire_N_609[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n51421), .O(one_wire_N_609[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48325_3_lut (.I0(n70708), .I1(n70702), .I2(color_bit_N_631[2]), 
            .I3(GND_net), .O(n64499));
    defparam i48325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48327_4_lut (.I0(n64500), .I1(n70696), .I2(n53961), .I3(color_bit_N_631[2]), 
            .O(n64501));
    defparam i48327_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i29552_4_lut (.I0(n64501), .I1(n57_adj_5836), .I2(n64499), 
            .I3(n65606), .O(state_3__N_560[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i29552_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY sub_14_add_2_11 (.CI(n51421), .I0(timer[9]), .I1(n1[9]), 
            .CO(n51422));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n51420), .O(one_wire_N_609[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n51420), .I0(timer[8]), .I1(n1[8]), 
            .CO(n51421));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(VCC_net), .D(n57810));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n51419), .O(one_wire_N_609[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_2047__i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(n35244), 
            .D(color_bit_N_631[1]), .R(n35253));   // verilog/neopixel.v(68[23:32])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n30014));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n30013));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_2047__i2 (.Q(bit_ctr[2]), .C(clk16MHz), .E(n35244), 
            .D(n13[2]), .R(n35253));   // verilog/neopixel.v(68[23:32])
    SB_DFFESR bit_ctr_2047__i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n35244), 
            .D(n13[3]), .R(n35253));   // verilog/neopixel.v(68[23:32])
    SB_DFF timer_2048__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY sub_14_add_2_9 (.CI(n51419), .I0(timer[7]), .I1(n1[7]), .CO(n51420));
    SB_DFFESR bit_ctr_2047__i4 (.Q(bit_ctr[4]), .C(clk16MHz), .E(n35244), 
            .D(n13[4]), .R(n35253));   // verilog/neopixel.v(68[23:32])
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n51418), .O(one_wire_N_609[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_2047__i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n35244), 
            .D(n13[0]), .R(n35253));   // verilog/neopixel.v(68[23:32])
    SB_DFF timer_2048__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2048__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY sub_14_add_2_8 (.CI(n51418), .I0(timer[6]), .I1(n1[6]), .CO(n51419));
    SB_LUT4 bit_ctr_0__bdd_4_lut_54526_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n70693));
    defparam bit_ctr_0__bdd_4_lut_54526_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_54531_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n70699));
    defparam bit_ctr_0__bdd_4_lut_54531_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n70705));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_DFF start_103 (.Q(start), .C(clk16MHz), .D(n57856));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n51417), .O(one_wire_N_609[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n40932), 
            .I3(\neo_pixel_transmitter.done ), .O(n62274));   // verilog/neopixel.v(16[11:16])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0002;
    SB_CARRY sub_14_add_2_7 (.CI(n51417), .I0(timer[5]), .I1(n1[5]), .CO(n51418));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk16MHz), .E(n7_adj_5835), 
            .D(state_3__N_560[0]), .S(n29225));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n51416), .O(one_wire_N_609[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n29784));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk16MHz), .E(n60097), .D(\neo_pixel_transmitter.done_N_651 ), 
            .R(n62274));   // verilog/neopixel.v(34[12] 116[6])
    SB_CARRY sub_14_add_2_6 (.CI(n51416), .I0(timer[4]), .I1(n1[4]), .CO(n51417));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n51415), .O(one_wire_N_609[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n51415), .I0(timer[3]), .I1(n1[3]), .CO(n51416));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n51414), .O(one_wire_N_609[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n51414), .I0(timer[2]), .I1(n1[2]), .CO(n51415));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_609[2]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n51413), .O(n4_adj_5838)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_3 (.CI(n51413), .I0(timer[1]), .I1(n1[1]), .CO(n51414));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n51413));
    SB_LUT4 i2_2_lut_4_lut (.I0(LED_c), .I1(n57_adj_5836), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n35253));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i30447_2_lut_3_lut (.I0(bit_ctr[3]), .I1(n44641), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n44751));
    defparam i30447_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[3]), .I1(n44641), .I2(bit_ctr[4]), 
            .I3(GND_net), .O(n53961));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_2_lut_3_lut_adj_1740 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_631[2]));
    defparam i1_2_lut_3_lut_adj_1740.LUT_INIT = 16'h1e1e;
    SB_LUT4 i30341_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n44641));
    defparam i30341_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i36812_1_lut (.I0(bit_ctr[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(68[23:32])
    defparam i36812_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36817_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n51094));   // verilog/neopixel.v(68[23:32])
    defparam i36817_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36828_2_lut_3_lut_4_lut (.I0(bit_ctr[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(bit_ctr[3]), .O(n13[3]));   // verilog/neopixel.v(68[23:32])
    defparam i36828_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i43857_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n59983));
    defparam i43857_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26619_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_645 ));   // verilog/neopixel.v(16[11:16])
    defparam i26619_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i36835_3_lut_4_lut (.I0(bit_ctr[2]), .I1(n51094), .I2(bit_ctr[3]), 
            .I3(bit_ctr[4]), .O(n13[4]));   // verilog/neopixel.v(68[23:32])
    defparam i36835_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i54504_2_lut_3_lut (.I0(start), .I1(\state[1] ), .I2(n59023), 
            .I3(GND_net), .O(n59025));
    defparam i54504_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i36821_2_lut_3_lut (.I0(bit_ctr[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(68[23:32])
    defparam i36821_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_3_lut (.I0(color_bit_N_631[2]), .I1(n53961), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n8_adj_5839));
    defparam i3_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1095_4_lut (.I0(color_bit_N_631[1]), .I1(n44751), .I2(n8_adj_5839), 
            .I3(n53940), .O(n57_adj_5836));   // verilog/neopixel.v(21[26:38])
    defparam i1095_4_lut.LUT_INIT = 16'h3233;
    SB_LUT4 i2_3_lut (.I0(LED_c), .I1(n57_adj_5836), .I2(\state[0] ), 
            .I3(GND_net), .O(n38));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i20852_3_lut (.I0(n25), .I1(n38), .I2(\state[1] ), .I3(GND_net), 
            .O(n35244));   // verilog/neopixel.v(16[11:16])
    defparam i20852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(one_wire_N_609[10]), .I1(one_wire_N_609[8]), .I2(one_wire_N_609[6]), 
            .I3(one_wire_N_609[7]), .O(n12_adj_5840));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_609[4]), .I1(n12_adj_5840), .I2(one_wire_N_609[9]), 
            .I3(one_wire_N_609[5]), .O(n35229));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i59_4_lut (.I0(n35229), .I1(n19), .I2(n4), .I3(\state[0] ), 
            .O(n43));   // verilog/neopixel.v(16[11:16])
    defparam i59_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i2_3_lut_adj_1741 (.I0(n43), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n25));   // verilog/neopixel.v(16[11:16])
    defparam i2_3_lut_adj_1741.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_1742 (.I0(bit_ctr[3]), .I1(n44641), .I2(GND_net), 
            .I3(GND_net), .O(n53940));
    defparam i1_2_lut_adj_1742.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1743 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_631[1]));
    defparam i1_2_lut_adj_1743.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1744 (.I0(color_bit_N_631[2]), .I1(n53961), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n8_adj_5841));
    defparam i3_3_lut_adj_1744.LUT_INIT = 16'h0404;
    SB_LUT4 i51182_4_lut (.I0(color_bit_N_631[1]), .I1(\state[0] ), .I2(n8_adj_5841), 
            .I3(n53940), .O(n67074));   // verilog/neopixel.v(16[11:16])
    defparam i51182_4_lut.LUT_INIT = 16'h7333;
    SB_LUT4 i26_4_lut (.I0(n25), .I1(n67074), .I2(\state[1] ), .I3(n44751), 
            .O(n57810));   // verilog/neopixel.v(16[11:16])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_609[3]), .I1(n4_adj_5838), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/neopixel.v(6[16:24])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1745 (.I0(one_wire_N_609[3]), .I1(one_wire_N_609[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/neopixel.v(52[15:25])
    defparam i1_2_lut_adj_1745.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(n4), .I1(n19), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n93));
    defparam i1_4_lut.LUT_INIT = 16'h5775;
    SB_LUT4 i48024_4_lut (.I0(one_wire_N_609[5]), .I1(one_wire_N_609[4]), 
            .I2(one_wire_N_609[6]), .I3(one_wire_N_609[8]), .O(n64189));
    defparam i48024_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47913_2_lut (.I0(one_wire_N_609[7]), .I1(one_wire_N_609[10]), 
            .I2(GND_net), .I3(GND_net), .O(n64077));
    defparam i47913_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut (.I0(n64077), .I1(n64189), .I2(one_wire_N_609[9]), 
            .I3(n93), .O(n59023));
    defparam i7_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_adj_1746 (.I0(\state[1] ), .I1(start), .I2(n59023), 
            .I3(GND_net), .O(n78));
    defparam i1_3_lut_adj_1746.LUT_INIT = 16'hbaba;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50967_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n40932), 
            .I3(GND_net), .O(n67077));   // verilog/neopixel.v(16[11:16])
    defparam i50967_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(52[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49432_2_lut_3_lut (.I0(n53961), .I1(bit_ctr[3]), .I2(n44641), 
            .I3(GND_net), .O(n65606));   // verilog/neopixel.v(21[26:38])
    defparam i49432_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 color_bit_N_631_1__bdd_4_lut (.I0(color_bit_N_631[1]), .I1(n64565), 
            .I2(n64566), .I3(color_bit_N_631[2]), .O(n70801));
    defparam color_bit_N_631_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n70801_bdd_4_lut (.I0(n70801), .I1(n64545), .I2(n64544), .I3(color_bit_N_631[2]), 
            .O(n70804));
    defparam n70801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i52512_3_lut_4_lut (.I0(start), .I1(\state[1] ), .I2(n68686), 
            .I3(n35229), .O(n68687));
    defparam i52512_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51526_2_lut_3_lut (.I0(one_wire_N_609[3]), .I1(one_wire_N_609[2]), 
            .I2(start), .I3(GND_net), .O(n67085));
    defparam i51526_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n70705_bdd_4_lut (.I0(n70705), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(color_bit_N_631[1]), .O(n70708));
    defparam n70705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70699_bdd_4_lut (.I0(n70699), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(color_bit_N_631[1]), .O(n70702));
    defparam n70699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n70693_bdd_4_lut (.I0(n70693), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_631[1]), .O(n70696));
    defparam n70693_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (ENCODER0_B_N_keep, n2270, ENCODER0_A_N_keep, 
            encoder0_position, GND_net, VCC_net, b_prev, \a_new[1] , 
            n30058, n2234, position_31__N_3956) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n2270;
    input ENCODER0_A_N_keep;
    output [31:0]encoder0_position;
    input GND_net;
    input VCC_net;
    output b_prev;
    output \a_new[1] ;
    input n30058;
    output n2234;
    output position_31__N_3956;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3964, debounce_cnt;
    wire [31:0]n133;
    
    wire direction_N_3961, n52808, n52807, n52806, n52805, n52804, 
        n52803, n52802, n52801, n52800, n52799, n52798, n52797, 
        n52796, n52795, n52794, n52793, n52792, n52791, n52790, 
        n52789, n52788, n52787, n52786, n52785, n52784, n52783, 
        n52782, n52781, n52780, n52779, n52778, n30098, a_prev, 
        n30091, position_31__N_3959;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2270), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n2270), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2270), .D(a_prev_N_3964));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2060_add_4_33_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[31]), .I3(n52808), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2060_add_4_32_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[30]), .I3(n52807), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_32 (.CI(n52807), .I0(direction_N_3961), 
            .I1(encoder0_position[30]), .CO(n52808));
    SB_LUT4 position_2060_add_4_31_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[29]), .I3(n52806), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_31 (.CI(n52806), .I0(direction_N_3961), 
            .I1(encoder0_position[29]), .CO(n52807));
    SB_LUT4 position_2060_add_4_30_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[28]), .I3(n52805), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_30 (.CI(n52805), .I0(direction_N_3961), 
            .I1(encoder0_position[28]), .CO(n52806));
    SB_LUT4 position_2060_add_4_29_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[27]), .I3(n52804), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_29 (.CI(n52804), .I0(direction_N_3961), 
            .I1(encoder0_position[27]), .CO(n52805));
    SB_LUT4 position_2060_add_4_28_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[26]), .I3(n52803), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_28 (.CI(n52803), .I0(direction_N_3961), 
            .I1(encoder0_position[26]), .CO(n52804));
    SB_LUT4 position_2060_add_4_27_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[25]), .I3(n52802), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_27 (.CI(n52802), .I0(direction_N_3961), 
            .I1(encoder0_position[25]), .CO(n52803));
    SB_LUT4 position_2060_add_4_26_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[24]), .I3(n52801), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_26 (.CI(n52801), .I0(direction_N_3961), 
            .I1(encoder0_position[24]), .CO(n52802));
    SB_LUT4 position_2060_add_4_25_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[23]), .I3(n52800), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_25 (.CI(n52800), .I0(direction_N_3961), 
            .I1(encoder0_position[23]), .CO(n52801));
    SB_LUT4 position_2060_add_4_24_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[22]), .I3(n52799), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_24 (.CI(n52799), .I0(direction_N_3961), 
            .I1(encoder0_position[22]), .CO(n52800));
    SB_LUT4 position_2060_add_4_23_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[21]), .I3(n52798), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_23 (.CI(n52798), .I0(direction_N_3961), 
            .I1(encoder0_position[21]), .CO(n52799));
    SB_LUT4 position_2060_add_4_22_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[20]), .I3(n52797), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_22 (.CI(n52797), .I0(direction_N_3961), 
            .I1(encoder0_position[20]), .CO(n52798));
    SB_LUT4 position_2060_add_4_21_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[19]), .I3(n52796), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_21 (.CI(n52796), .I0(direction_N_3961), 
            .I1(encoder0_position[19]), .CO(n52797));
    SB_LUT4 position_2060_add_4_20_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[18]), .I3(n52795), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_20 (.CI(n52795), .I0(direction_N_3961), 
            .I1(encoder0_position[18]), .CO(n52796));
    SB_LUT4 position_2060_add_4_19_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[17]), .I3(n52794), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_19 (.CI(n52794), .I0(direction_N_3961), 
            .I1(encoder0_position[17]), .CO(n52795));
    SB_LUT4 position_2060_add_4_18_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[16]), .I3(n52793), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_18 (.CI(n52793), .I0(direction_N_3961), 
            .I1(encoder0_position[16]), .CO(n52794));
    SB_LUT4 position_2060_add_4_17_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[15]), .I3(n52792), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_17 (.CI(n52792), .I0(direction_N_3961), 
            .I1(encoder0_position[15]), .CO(n52793));
    SB_LUT4 position_2060_add_4_16_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[14]), .I3(n52791), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_16 (.CI(n52791), .I0(direction_N_3961), 
            .I1(encoder0_position[14]), .CO(n52792));
    SB_LUT4 position_2060_add_4_15_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[13]), .I3(n52790), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_15 (.CI(n52790), .I0(direction_N_3961), 
            .I1(encoder0_position[13]), .CO(n52791));
    SB_LUT4 position_2060_add_4_14_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[12]), .I3(n52789), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_14 (.CI(n52789), .I0(direction_N_3961), 
            .I1(encoder0_position[12]), .CO(n52790));
    SB_LUT4 position_2060_add_4_13_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[11]), .I3(n52788), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_13 (.CI(n52788), .I0(direction_N_3961), 
            .I1(encoder0_position[11]), .CO(n52789));
    SB_LUT4 position_2060_add_4_12_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[10]), .I3(n52787), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_12 (.CI(n52787), .I0(direction_N_3961), 
            .I1(encoder0_position[10]), .CO(n52788));
    SB_LUT4 position_2060_add_4_11_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[9]), .I3(n52786), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_11 (.CI(n52786), .I0(direction_N_3961), 
            .I1(encoder0_position[9]), .CO(n52787));
    SB_LUT4 position_2060_add_4_10_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[8]), .I3(n52785), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_10 (.CI(n52785), .I0(direction_N_3961), 
            .I1(encoder0_position[8]), .CO(n52786));
    SB_LUT4 position_2060_add_4_9_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[7]), .I3(n52784), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_9 (.CI(n52784), .I0(direction_N_3961), 
            .I1(encoder0_position[7]), .CO(n52785));
    SB_LUT4 position_2060_add_4_8_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[6]), .I3(n52783), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_8 (.CI(n52783), .I0(direction_N_3961), 
            .I1(encoder0_position[6]), .CO(n52784));
    SB_LUT4 position_2060_add_4_7_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[5]), .I3(n52782), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_7 (.CI(n52782), .I0(direction_N_3961), 
            .I1(encoder0_position[5]), .CO(n52783));
    SB_LUT4 position_2060_add_4_6_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[4]), .I3(n52781), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_6 (.CI(n52781), .I0(direction_N_3961), 
            .I1(encoder0_position[4]), .CO(n52782));
    SB_LUT4 position_2060_add_4_5_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[3]), .I3(n52780), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_5 (.CI(n52780), .I0(direction_N_3961), 
            .I1(encoder0_position[3]), .CO(n52781));
    SB_LUT4 position_2060_add_4_4_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[2]), .I3(n52779), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_4 (.CI(n52779), .I0(direction_N_3961), 
            .I1(encoder0_position[2]), .CO(n52780));
    SB_LUT4 position_2060_add_4_3_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder0_position[1]), .I3(n52778), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_3 (.CI(n52778), .I0(direction_N_3961), 
            .I1(encoder0_position[1]), .CO(n52779));
    SB_LUT4 position_2060_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2060_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2060_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n52778));
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2270), .D(n30098));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3961));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2270), .D(n30091));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n2234), .C(n2270), .D(n30058));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2060__i0 (.Q(encoder0_position[0]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i31 (.Q(encoder0_position[31]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i30 (.Q(encoder0_position[30]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i29 (.Q(encoder0_position[29]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i28 (.Q(encoder0_position[28]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i27 (.Q(encoder0_position[27]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i26 (.Q(encoder0_position[26]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i25 (.Q(encoder0_position[25]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i24 (.Q(encoder0_position[24]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i23 (.Q(encoder0_position[23]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i22 (.Q(encoder0_position[22]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i21 (.Q(encoder0_position[21]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i20 (.Q(encoder0_position[20]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i19 (.Q(encoder0_position[19]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i18 (.Q(encoder0_position[18]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i17 (.Q(encoder0_position[17]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i16 (.Q(encoder0_position[16]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i15 (.Q(encoder0_position[15]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i14 (.Q(encoder0_position[14]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i13 (.Q(encoder0_position[13]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i12 (.Q(encoder0_position[12]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i11 (.Q(encoder0_position[11]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i10 (.Q(encoder0_position[10]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i9 (.Q(encoder0_position[9]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i8 (.Q(encoder0_position[8]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i7 (.Q(encoder0_position[7]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i6 (.Q(encoder0_position[6]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i5 (.Q(encoder0_position[5]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i4 (.Q(encoder0_position[4]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i3 (.Q(encoder0_position[3]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i2 (.Q(encoder0_position[2]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2060__i1 (.Q(encoder0_position[1]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 i53778_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3964));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i53778_4_lut.LUT_INIT = 16'h8421;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n2270), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2270), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15691_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3964), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n30098));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15691_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15684_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3964), .I2(b_new[1]), 
            .I3(b_prev), .O(n30091));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3959));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3959), 
            .I3(\a_new[1] ), .O(position_31__N_3956));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (ENCODER1_B_N_keep, n2270, ENCODER1_A_N_keep, 
            b_prev, n30060, n2275, position_31__N_3956, encoder1_position, 
            GND_net, \a_new[1] , VCC_net) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n2270;
    input ENCODER1_A_N_keep;
    output b_prev;
    input n30060;
    output n2275;
    output position_31__N_3956;
    output [31:0]encoder1_position;
    input GND_net;
    output \a_new[1] ;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3964, debounce_cnt, n30100, n30099, a_prev;
    wire [31:0]n133;
    
    wire direction_N_3961, n52764, n52763, n52762, n52761, n52760, 
        n52759, n52758, n52757, n52756, n52755, n52754, n52753, 
        n52752, n52751, n52750, n52749, n52748, n52747, n52746, 
        n52745, n52744, n52743, n52742, n52741, n52740, n52739, 
        n52738, n52737, n52736, n52735, n52734, position_31__N_3959;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n2270), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n2270), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n2270), .D(a_prev_N_3964));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n2270), .D(n30100));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n2270), .D(n30099));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n2275), .C(n2270), .D(n30060));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i0 (.Q(encoder1_position[0]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i31 (.Q(encoder1_position[31]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(encoder1_position[30]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(encoder1_position[29]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(encoder1_position[28]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(encoder1_position[27]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(encoder1_position[26]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(encoder1_position[25]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(encoder1_position[24]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(encoder1_position[23]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(encoder1_position[22]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(encoder1_position[21]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(encoder1_position[20]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(encoder1_position[19]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(encoder1_position[18]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(encoder1_position[17]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(encoder1_position[16]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(encoder1_position[15]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(encoder1_position[14]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(encoder1_position[13]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(encoder1_position[12]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(encoder1_position[11]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(encoder1_position[10]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(encoder1_position[9]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(encoder1_position[8]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(encoder1_position[7]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(encoder1_position[6]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(encoder1_position[5]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(encoder1_position[4]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(encoder1_position[3]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(encoder1_position[2]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(encoder1_position[1]), .C(n2270), .E(position_31__N_3956), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[31]), .I3(n52764), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[30]), .I3(n52763), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n52763), .I0(direction_N_3961), 
            .I1(encoder1_position[30]), .CO(n52764));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[29]), .I3(n52762), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n52762), .I0(direction_N_3961), 
            .I1(encoder1_position[29]), .CO(n52763));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[28]), .I3(n52761), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n52761), .I0(direction_N_3961), 
            .I1(encoder1_position[28]), .CO(n52762));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[27]), .I3(n52760), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n52760), .I0(direction_N_3961), 
            .I1(encoder1_position[27]), .CO(n52761));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[26]), .I3(n52759), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n52759), .I0(direction_N_3961), 
            .I1(encoder1_position[26]), .CO(n52760));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[25]), .I3(n52758), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n52758), .I0(direction_N_3961), 
            .I1(encoder1_position[25]), .CO(n52759));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[24]), .I3(n52757), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n52757), .I0(direction_N_3961), 
            .I1(encoder1_position[24]), .CO(n52758));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[23]), .I3(n52756), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n52756), .I0(direction_N_3961), 
            .I1(encoder1_position[23]), .CO(n52757));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[22]), .I3(n52755), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n52755), .I0(direction_N_3961), 
            .I1(encoder1_position[22]), .CO(n52756));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[21]), .I3(n52754), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n52754), .I0(direction_N_3961), 
            .I1(encoder1_position[21]), .CO(n52755));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[20]), .I3(n52753), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n52753), .I0(direction_N_3961), 
            .I1(encoder1_position[20]), .CO(n52754));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[19]), .I3(n52752), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n52752), .I0(direction_N_3961), 
            .I1(encoder1_position[19]), .CO(n52753));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[18]), .I3(n52751), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n52751), .I0(direction_N_3961), 
            .I1(encoder1_position[18]), .CO(n52752));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[17]), .I3(n52750), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n52750), .I0(direction_N_3961), 
            .I1(encoder1_position[17]), .CO(n52751));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[16]), .I3(n52749), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n52749), .I0(direction_N_3961), 
            .I1(encoder1_position[16]), .CO(n52750));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[15]), .I3(n52748), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n52748), .I0(direction_N_3961), 
            .I1(encoder1_position[15]), .CO(n52749));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[14]), .I3(n52747), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n52747), .I0(direction_N_3961), 
            .I1(encoder1_position[14]), .CO(n52748));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[13]), .I3(n52746), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n52746), .I0(direction_N_3961), 
            .I1(encoder1_position[13]), .CO(n52747));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[12]), .I3(n52745), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n52745), .I0(direction_N_3961), 
            .I1(encoder1_position[12]), .CO(n52746));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[11]), .I3(n52744), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n52744), .I0(direction_N_3961), 
            .I1(encoder1_position[11]), .CO(n52745));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[10]), .I3(n52743), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n52743), .I0(direction_N_3961), 
            .I1(encoder1_position[10]), .CO(n52744));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[9]), .I3(n52742), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n52742), .I0(direction_N_3961), 
            .I1(encoder1_position[9]), .CO(n52743));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[8]), .I3(n52741), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n52741), .I0(direction_N_3961), 
            .I1(encoder1_position[8]), .CO(n52742));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[7]), .I3(n52740), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n52740), .I0(direction_N_3961), 
            .I1(encoder1_position[7]), .CO(n52741));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[6]), .I3(n52739), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n52739), .I0(direction_N_3961), 
            .I1(encoder1_position[6]), .CO(n52740));
    SB_LUT4 i53781_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3964));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i53781_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[5]), .I3(n52738), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n52738), .I0(direction_N_3961), 
            .I1(encoder1_position[5]), .CO(n52739));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[4]), .I3(n52737), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n2270), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_2054_add_4_6 (.CI(n52737), .I0(direction_N_3961), 
            .I1(encoder1_position[4]), .CO(n52738));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[3]), .I3(n52736), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n52736), .I0(direction_N_3961), 
            .I1(encoder1_position[3]), .CO(n52737));
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n2270), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[2]), .I3(n52735), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n52735), .I0(direction_N_3961), 
            .I1(encoder1_position[2]), .CO(n52736));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3961), 
            .I2(encoder1_position[1]), .I3(n52734), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n52734), .I0(direction_N_3961), 
            .I1(encoder1_position[1]), .CO(n52735));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n52734));
    SB_LUT4 i15693_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3964), .I2(b_new[1]), 
            .I3(b_prev), .O(n30100));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15693_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15692_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3964), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n30099));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15692_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3959));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3959), 
            .I3(\a_new[1] ), .O(position_31__N_3956));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3961));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\data[12] , GND_net, clk16MHz, n30250, \data[15] , 
            n30249, n30248, \data[11] , n30247, \data[10] , n30246, 
            \data[9] , n30245, \data[8] , n30244, \data[7] , n30243, 
            \data[6] , n30242, \data[5] , n30241, \data[4] , n30240, 
            \data[3] , n30239, \data[2] , n30238, \data[1] , \state[0] , 
            n15, clk_out, CS_c, CS_CLK_c, VCC_net, n6, \state[1] , 
            n9, n30025, n30023, \current[0] , n6_adj_26, n6_adj_27, 
            state_7__N_4446, n43986, n30855, \data[0] , n30759, \current[1] , 
            n30758, \current[2] , n30757, \current[3] , n30756, \current[4] , 
            n30755, \current[5] , n30754, \current[6] , n30753, \current[7] , 
            n30752, \current[8] , n30751, \current[9] , n30750, \current[10] , 
            n30749, \current[11] , n28109, \current[15] , n11, n25959, 
            n25966, n25977, n25971) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \data[12] ;
    input GND_net;
    input clk16MHz;
    input n30250;
    output \data[15] ;
    input n30249;
    input n30248;
    output \data[11] ;
    input n30247;
    output \data[10] ;
    input n30246;
    output \data[9] ;
    input n30245;
    output \data[8] ;
    input n30244;
    output \data[7] ;
    input n30243;
    output \data[6] ;
    input n30242;
    output \data[5] ;
    input n30241;
    output \data[4] ;
    input n30240;
    output \data[3] ;
    input n30239;
    output \data[2] ;
    input n30238;
    output \data[1] ;
    output \state[0] ;
    output n15;
    output clk_out;
    output CS_c;
    output CS_CLK_c;
    input VCC_net;
    output n6;
    output \state[1] ;
    input n9;
    input n30025;
    input n30023;
    output \current[0] ;
    output n6_adj_26;
    output n6_adj_27;
    output state_7__N_4446;
    output n43986;
    input n30855;
    output \data[0] ;
    input n30759;
    output \current[1] ;
    input n30758;
    output \current[2] ;
    input n30757;
    output \current[3] ;
    input n30756;
    output \current[4] ;
    input n30755;
    output \current[5] ;
    input n30754;
    output \current[6] ;
    input n30753;
    output \current[7] ;
    input n30752;
    output \current[8] ;
    input n30751;
    output \current[9] ;
    input n30750;
    output \current[10] ;
    input n30749;
    output \current[11] ;
    output n28109;
    output \current[15] ;
    output n11;
    output n25959;
    output n25966;
    output n25977;
    output n25971;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [13:0]n241;
    
    wire clk_slow_N_4359, n7225, n44482;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n52777, n52776;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n12596, n28347, n29231;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n52775, n52774, n52773, n52772, n52771, n52770, n52769, 
        n23048, n28164;
    wire [7:0]n37;
    
    wire n29529, delay_counter_15__N_4441, clk_slow_N_4360, n52768, 
        n52767, n52766, n52765, n23050, n23052, n23054, n52671, 
        n52670, n52669, n52668, n67003, n52667, n66920, n52666, 
        n66939, n52665, n66948, n6_adj_5834, n8, n12, n10;
    
    SB_LUT4 i2202_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2202_1_lut.LUT_INIT = 16'h5555;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4359));   // verilog/tli4970.v(13[10] 19[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n30250));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n30249));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n30248));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n30247));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n30246));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n30245));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n30244));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n30243));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n30242));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n30241));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n30240));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n30239));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n30238));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i6091_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n7225));   // verilog/tli4970.v(43[5] 67[12])
    defparam i6091_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53788_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n44482));
    defparam i53788_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 counter_2058_2059_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52777), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2058_2059_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2058_2059_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52776), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2058_2059_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2058_2059_add_4_3 (.CI(n52776), .I0(GND_net), .I1(counter[1]), 
            .CO(n52777));
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 counter_2058_2059_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2058_2059_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2058_2059_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52776));
    SB_LUT4 equal_374_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_374_i6_2_lut.LUT_INIT = 16'heeee;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28347), .D(n12596), 
            .R(n29231));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n30025));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n30023));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 delay_counter_2056_2057_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n52775), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2056_2057_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n52774), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_12 (.CI(n52774), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n52775));
    SB_LUT4 delay_counter_2056_2057_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n52773), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_11 (.CI(n52773), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n52774));
    SB_LUT4 delay_counter_2056_2057_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n52772), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_372_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_26));   // verilog/tli4970.v(54[9:26])
    defparam equal_372_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_CARRY delay_counter_2056_2057_add_4_10 (.CI(n52772), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n52773));
    SB_LUT4 delay_counter_2056_2057_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n52771), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_9 (.CI(n52771), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n52772));
    SB_LUT4 delay_counter_2056_2057_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n52770), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_8 (.CI(n52770), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n52771));
    SB_LUT4 delay_counter_2056_2057_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n52769), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFNE bit_counter_2050__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28164), 
            .D(n23048));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2050__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28164), 
            .D(n37[4]), .R(n29529));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2056_2057__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2058_2059__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4360));   // verilog/tli4970.v(14[16:27])
    SB_CARRY delay_counter_2056_2057_add_4_7 (.CI(n52769), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n52770));
    SB_LUT4 delay_counter_2056_2057_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n52768), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_6 (.CI(n52768), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n52769));
    SB_DFFSR counter_2058_2059__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4360));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2058_2059__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4360));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 delay_counter_2056_2057_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n52767), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_5 (.CI(n52767), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n52768));
    SB_LUT4 delay_counter_2056_2057_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n52766), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_4 (.CI(n52766), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n52767));
    SB_LUT4 delay_counter_2056_2057_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n52765), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2056_2057_add_4_3 (.CI(n52765), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n52766));
    SB_LUT4 delay_counter_2056_2057_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2056_2057_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFNSR delay_counter_2056_2057__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2056_2057__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4441));   // verilog/tli4970.v(40[24:39])
    SB_LUT4 equal_367_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_27));   // verilog/tli4970.v(54[9:26])
    defparam equal_367_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4446));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i29691_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n43986));
    defparam i29691_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNESR bit_counter_2050__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28164), 
            .D(n37[5]), .R(n29529));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2050__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28164), 
            .D(n37[6]), .R(n29529));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2050__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28164), 
            .D(n37[7]), .R(n29529));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2050__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28164), 
            .D(n23050));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2050__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28164), 
            .D(n23052));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2050__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28164), 
            .D(n23054));   // verilog/tli4970.v(55[24:39])
    SB_CARRY delay_counter_2056_2057_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n52765));
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30855));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30759));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30758));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30757));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30756));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30755));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30754));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30753));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30752));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30751));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30750));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30749));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28109), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 equal_302_i11_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_302_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n25959));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1737 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[1]), .I3(bit_counter[0]), .O(n25966));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1737.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1738 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[1]), .I3(bit_counter[0]), .O(n25977));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1738.LUT_INIT = 16'hffbf;
    SB_LUT4 i2174_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4360));
    defparam i2174_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4360), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4359));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28347), .D(n44482), 
            .S(n29231));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 bit_counter_2050_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n52671), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2050_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n52670), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2050_add_4_8 (.CI(n52670), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n52671));
    SB_LUT4 bit_counter_2050_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n52669), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2050_add_4_7 (.CI(n52669), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n52670));
    SB_LUT4 bit_counter_2050_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n52668), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2050_add_4_6 (.CI(n52668), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n52669));
    SB_LUT4 bit_counter_2050_add_4_5_lut (.I0(n7225), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n52667), .O(n67003)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2050_add_4_5 (.CI(n52667), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n52668));
    SB_LUT4 bit_counter_2050_add_4_4_lut (.I0(n7225), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n52666), .O(n66920)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2050_add_4_4 (.CI(n52666), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n52667));
    SB_LUT4 bit_counter_2050_add_4_3_lut (.I0(n7225), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n52665), .O(n66939)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2050_add_4_3 (.CI(n52665), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n52666));
    SB_LUT4 bit_counter_2050_add_4_2_lut (.I0(n7225), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n66948)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2050_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2050_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n52665));
    SB_LUT4 i8895_3_lut (.I0(\state[0] ), .I1(n66939), .I2(\state[1] ), 
            .I3(GND_net), .O(n23054));   // verilog/tli4970.v(55[24:39])
    defparam i8895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8893_3_lut (.I0(\state[0] ), .I1(n66920), .I2(\state[1] ), 
            .I3(GND_net), .O(n23052));   // verilog/tli4970.v(55[24:39])
    defparam i8893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8891_3_lut (.I0(\state[0] ), .I1(n67003), .I2(\state[1] ), 
            .I3(GND_net), .O(n23050));   // verilog/tli4970.v(55[24:39])
    defparam i8891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4441), .O(n28347));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i14824_2_lut_4_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(delay_counter_15__N_4441), .O(n29231));
    defparam i14824_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_LUT4 i13984_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28164));
    defparam i13984_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8889_3_lut (.I0(\state[0] ), .I1(n66948), .I2(\state[1] ), 
            .I3(GND_net), .O(n23048));   // verilog/tli4970.v(55[24:39])
    defparam i8889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53763_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n28109));
    defparam i53763_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i15123_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29529));   // verilog/tli4970.v(55[24:39])
    defparam i15123_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5834));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_5834), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2175_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2175_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_1739 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_1739.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4441));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2142_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n12596));
    defparam mux_2142_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n25971));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    
endmodule
//
// Verilog Description of module coms
//

module coms (VCC_net, \data_in_frame[4] , clk16MHz, \data_in_frame[2] , 
            \data_in_frame[1] , n3358, \data_out_frame[6] , n58972, 
            \data_in_frame[11] , IntegralLimit, n58971, GND_net, \data_in_frame[0] , 
            \data_out_frame[5] , \FRAME_MATCHER.i_31__N_2638 , control_mode, 
            n58970, \data_in_frame[12] , \data_out_frame[7] , n58969, 
            \data_out_frame[20] , displacement, \data_out_frame[4] , ID, 
            \data_in_frame[16] , deadband, byte_transmit_counter, \data_out_frame[0][2] , 
            \data_out_frame[18] , \data_out_frame[19] , \data_out_frame[16] , 
            \data_out_frame[17] , \byte_transmit_counter[1] , \byte_transmit_counter[2] , 
            n28, n379, n405, n4, encoder0_position_scaled, \FRAME_MATCHER.state[3] , 
            \FRAME_MATCHER.i[3] , \FRAME_MATCHER.i[4] , n8, \data_in_frame[14] , 
            n58968, n58967, n58966, n58965, n59004, n58964, reset, 
            setpoint, \data_out_frame[3][7] , n58963, \data_out_frame[8] , 
            n58962, n58961, n58960, n58959, n58958, n58957, n58825, 
            n58956, \data_out_frame[9] , n58955, n58954, n58953, n58952, 
            n58951, n30260, n30257, n149, n11, \data_out_frame[12] , 
            \data_out_frame[13] , \data_out_frame[14] , \data_out_frame[15] , 
            \data_out_frame[3][6] , \data_out_frame[1][6] , n70864, \data_out_frame[1][7] , 
            \data_out_frame[3][4] , \data_out_frame[3][3] , \data_out_frame[10] , 
            \data_out_frame[11] , \data_out_frame[3][1] , n28507, \data_out_frame[1][5] , 
            n58950, \data_out_frame[0][3] , \data_out_frame[1][3] , n58949, 
            n58948, n58947, n58946, n58945, n58944, n58943, n58942, 
            n58941, n58940, n60, n51, n58939, n58938, n58937, 
            n58936, n28717, n28774, rx_data, \data_out_frame[22] , 
            \data_out_frame[23] , \data_out_frame[21] , n30228, n30225, 
            n58935, n30222, n30219, n30216, n30208, n30207, neopxl_color, 
            \data_in_frame[18] , \data_in_frame[21] , \data_in_frame[20][7] , 
            \data_in_frame[17] , \data_in_frame[20][1] , \data_in_frame[20][5] , 
            \data_in_frame[8] , n25605, n59499, n61411, encoder1_position_scaled, 
            \data_in_frame[6] , \motor_state_23__N_115[13] , n15, n10, 
            n58934, n58933, n58932, n58931, n58930, n58929, n58928, 
            n58927, n58926, \Kp[1] , \Kp[2] , \Kp[3] , n58925, \Kp[4] , 
            n58924, n58826, \Kp[5] , \Kp[6] , \Kp[7] , n58923, n58922, 
            n58921, \Kp[8] , n58920, \Kp[9] , \Kp[10] , \Kp[11] , 
            \Kp[12] , n58919, n58918, n58917, \Kp[13] , \Kp[14] , 
            \Kp[15] , n58916, n58915, \Ki[1] , n58914, n58913, n58912, 
            \Ki[2] , \data_out_frame[24] , \Ki[3] , \Ki[4] , \Ki[5] , 
            \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , 
            \Ki[12] , \Ki[13] , n26902, n58911, n58910, \Ki[14] , 
            \Ki[15] , n30130, current_limit, n30129, n30128, n30127, 
            n58909, n58908, n58907, n58906, n30126, n30125, n30124, 
            n30123, n30121, PWMLimit, n58905, n58904, n58903, n58902, 
            n58901, \data_in_frame[20][0] , n59138, n30090, \FRAME_MATCHER.rx_data_ready_prev , 
            n59971, n30075, n30074, n59994, \data_in_frame[8][7] , 
            n58900, n28801, \data_in_frame[6][2] , n30073, n30072, 
            n30068, n30067, n30066, \data_out_frame[25] , n30062, 
            n30061, n30059, n30057, n30010, \Ki[0] , \Kp[0] , n58899, 
            n58829, n58832, n58833, n58834, n58835, n58836, n58841, 
            n58843, n58847, n58848, n58849, n58850, n58844, n58851, 
            n58852, n58846, n58853, n58854, n58855, n58856, n58857, 
            n58858, n58859, n58827, \data_in_frame[17][7] , \data_in_frame[17][6] , 
            n58860, n58861, n58862, n58863, n58864, DE_c, tx_active, 
            LED_c, n58845, n59003, n58865, \data_in_frame[7][7] , 
            \data_in_frame[5] , \data_out_frame[0][4] , n59002, \data_in_frame[7][2] , 
            \data_in_frame[6][7] , n58866, \data_out_frame[1][0] , n59001, 
            n28780, \data_in_frame[7][0] , \data_out_frame[1][1] , n59000, 
            n58999, n31074, n29319, n31075, n29318, n58998, \data_in_frame[8][4] , 
            \data_in_frame[7][4] , \data_in_frame[8][5] , \data_in_frame[6][3] , 
            \data_in_frame[7][3] , \data_in_frame[7][5] , n30842, n30828, 
            n23230, n30773, n30763, n30761, n30760, n30744, n30742, 
            \data_in_frame[6][1] , n30710, n30707, n30706, n30705, 
            n30703, n30702, n58296, n29833, n30693, n30690, n58294, 
            n58290, n58286, n58282, n58278, n58274, n58272, n58268, 
            n29861, n58264, n29867, n58260, n30677, n30674, n58256, 
            n30672, n30669, n30664, n30338, n30342, n30348, n30352, 
            \data_in_frame[6][4] , n30361, n30365, n30368, \data_in_frame[7][1] , 
            n30371, n30375, n30378, n30381, n30387, n30399, \data_in_frame[8][3] , 
            n30403, n30639, n30638, n30406, n30409, n30413, n30466, 
            n30469, n30616, n30475, n30479, n30482, n30485, n30489, 
            n30492, n30495, n30499, n58384, n58398, n30509, n30512, 
            n30515, n30550, n30554, n30558, n30562, n30566, n30587, 
            n58252, n58248, n58244, \data_in_frame[20][2] , n29909, 
            \data_in_frame[20][3] , n29912, \data_in_frame[20][4] , n58238, 
            n58234, n58230, n58228, n58226, n58224, n58220, n58216, 
            n58212, n58208, n29949, \data_in_frame[22] , n29952, n58202, 
            n29958, n29961, n29964, n29968, n58198, n30539, n29977, 
            \data_in_frame[23] , n29980, n29983, n29986, n29989, n29992, 
            n29995, n30465, n30003, n30016, n30028, n30031, n30035, 
            n58340, n58997, n58996, n58995, n58994, n58842, n31082, 
            n29317, n58993, n58992, n58991, n58990, \data_in_frame[1][1] , 
            n58989, n58988, rx_data_ready, n59967, n58867, n58868, 
            n58987, n58986, n58985, n58984, n58869, n58840, n58839, 
            n58983, n58982, n58981, n58870, n42166, n28770, n58871, 
            n59086, n29311, n58872, n58873, n58874, n58875, n58876, 
            n58877, n58878, n8_adj_10, n28725, n58879, n58838, n58880, 
            n58837, n58881, n58882, n8_adj_11, n8_adj_12, n28733, 
            n58980, n58979, n58883, n58978, n58977, n58884, n58885, 
            n58831, n58830, n58886, n58887, n58888, n58889, n58890, 
            n58891, n58892, n58893, n58894, n29283, \data_out_frame[27][6] , 
            \data_out_frame[26][6] , n58895, n58824, n31162, n29256, 
            n31163, n29255, n31164, n29254, n58896, n31166, n29251, 
            n58897, n58898, n58828, n58976, n59079, n58975, n58974, 
            n58973, n69908, n28778, n69906, n26087, n59593, n26490, 
            n54003, pwm_setpoint, n23164, n44625, n64453, n64451, 
            n59093, n28719, n28723, n35592, n15_adj_13, n54986, 
            n59975, n28791, \current[7] , \current[6] , \current[5] , 
            \current[4] , \current[3] , \current[2] , \current[1] , 
            \current[0] , \current[15] , \current[11] , \current[10] , 
            \current[9] , \current[8] , \o_Rx_DV_N_3617[24] , r_SM_Main, 
            n27, n62584, n28320, n60079, n1, tx_o, r_Clock_Count, 
            n30034, n71131, n30847, \r_Bit_Index[0] , n6, tx_enable, 
            \o_Rx_DV_N_3617[12] , n5254, \o_Rx_DV_N_3617[8] , r_Rx_Data, 
            n29, n23, \r_SM_Main[1]_adj_14 , baudrate, n28324, n60053, 
            \r_SM_Main[2]_adj_15 , RX_N_2, r_Clock_Count_adj_25, n30256, 
            n30255, n30254, n30253, n30252, n25975, \o_Rx_DV_N_3617[7] , 
            \o_Rx_DV_N_3617[6] , \o_Rx_DV_N_3617[5] , \o_Rx_DV_N_3617[4] , 
            \o_Rx_DV_N_3617[3] , \o_Rx_DV_N_3617[2] , \o_Rx_DV_N_3617[1] , 
            \o_Rx_DV_N_3617[0] , \r_Bit_Index[0]_adj_24 , n62864, n29921, 
            n59011, n62764, n62780, n62748, n62828, n62812, n30854, 
            n55126, n30850, n5257, n29791, n28127, n62796, n62846) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    output [7:0]\data_in_frame[4] ;
    input clk16MHz;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[1] ;
    input n3358;
    output [7:0]\data_out_frame[6] ;
    input n58972;
    output [7:0]\data_in_frame[11] ;
    output [23:0]IntegralLimit;
    input n58971;
    input GND_net;
    output [7:0]\data_in_frame[0] ;
    output [7:0]\data_out_frame[5] ;
    output \FRAME_MATCHER.i_31__N_2638 ;
    output [7:0]control_mode;
    input n58970;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_out_frame[7] ;
    input n58969;
    output [7:0]\data_out_frame[20] ;
    input [23:0]displacement;
    output [7:0]\data_out_frame[4] ;
    input [7:0]ID;
    output [7:0]\data_in_frame[16] ;
    output [23:0]deadband;
    output [7:0]byte_transmit_counter;
    output \data_out_frame[0][2] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output \byte_transmit_counter[1] ;
    output \byte_transmit_counter[2] ;
    input n28;
    input n379;
    input n405;
    output n4;
    input [23:0]encoder0_position_scaled;
    output \FRAME_MATCHER.state[3] ;
    output \FRAME_MATCHER.i[3] ;
    output \FRAME_MATCHER.i[4] ;
    output n8;
    output [7:0]\data_in_frame[14] ;
    input n58968;
    input n58967;
    input n58966;
    input n58965;
    input n59004;
    input n58964;
    input reset;
    output [23:0]setpoint;
    output \data_out_frame[3][7] ;
    input n58963;
    output [7:0]\data_out_frame[8] ;
    input n58962;
    input n58961;
    input n58960;
    input n58959;
    input n58958;
    input n58957;
    input n58825;
    input n58956;
    output [7:0]\data_out_frame[9] ;
    input n58955;
    input n58954;
    input n58953;
    input n58952;
    input n58951;
    input n30260;
    input n30257;
    input n149;
    output n11;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output \data_out_frame[3][6] ;
    output \data_out_frame[1][6] ;
    input n70864;
    output \data_out_frame[1][7] ;
    output \data_out_frame[3][4] ;
    output \data_out_frame[3][3] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    output \data_out_frame[3][1] ;
    output n28507;
    output \data_out_frame[1][5] ;
    input n58950;
    output \data_out_frame[0][3] ;
    output \data_out_frame[1][3] ;
    input n58949;
    input n58948;
    input n58947;
    input n58946;
    input n58945;
    input n58944;
    input n58943;
    input n58942;
    input n58941;
    input n58940;
    output n60;
    output n51;
    input n58939;
    input n58938;
    input n58937;
    input n58936;
    output n28717;
    input n28774;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[21] ;
    input n30228;
    input n30225;
    input n58935;
    input n30222;
    input n30219;
    input n30216;
    input n30208;
    input n30207;
    output [23:0]neopxl_color;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[21] ;
    output \data_in_frame[20][7] ;
    output [7:0]\data_in_frame[17] ;
    output \data_in_frame[20][1] ;
    output \data_in_frame[20][5] ;
    output [7:0]\data_in_frame[8] ;
    input n25605;
    output n59499;
    input n61411;
    input [23:0]encoder1_position_scaled;
    output [7:0]\data_in_frame[6] ;
    input \motor_state_23__N_115[13] ;
    output n15;
    output n10;
    input n58934;
    input n58933;
    input n58932;
    input n58931;
    input n58930;
    input n58929;
    input n58928;
    input n58927;
    input n58926;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    input n58925;
    output \Kp[4] ;
    input n58924;
    input n58826;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    input n58923;
    input n58922;
    input n58921;
    output \Kp[8] ;
    input n58920;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    input n58919;
    input n58918;
    input n58917;
    output \Kp[13] ;
    output \Kp[14] ;
    output \Kp[15] ;
    input n58916;
    input n58915;
    output \Ki[1] ;
    input n58914;
    input n58913;
    input n58912;
    output \Ki[2] ;
    output [7:0]\data_out_frame[24] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output n26902;
    input n58911;
    input n58910;
    output \Ki[14] ;
    output \Ki[15] ;
    input n30130;
    output [15:0]current_limit;
    input n30129;
    input n30128;
    input n30127;
    input n58909;
    input n58908;
    input n58907;
    input n58906;
    input n30126;
    input n30125;
    input n30124;
    input n30123;
    input n30121;
    output [23:0]PWMLimit;
    input n58905;
    input n58904;
    input n58903;
    input n58902;
    input n58901;
    output \data_in_frame[20][0] ;
    input n59138;
    input n30090;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output n59971;
    input n30075;
    input n30074;
    output n59994;
    output \data_in_frame[8][7] ;
    input n58900;
    output n28801;
    output \data_in_frame[6][2] ;
    input n30073;
    input n30072;
    input n30068;
    input n30067;
    input n30066;
    output [7:0]\data_out_frame[25] ;
    input n30062;
    input n30061;
    input n30059;
    input n30057;
    input n30010;
    output \Ki[0] ;
    output \Kp[0] ;
    input n58899;
    input n58829;
    input n58832;
    input n58833;
    input n58834;
    input n58835;
    input n58836;
    input n58841;
    input n58843;
    input n58847;
    input n58848;
    input n58849;
    input n58850;
    input n58844;
    input n58851;
    input n58852;
    input n58846;
    input n58853;
    input n58854;
    input n58855;
    input n58856;
    input n58857;
    input n58858;
    input n58859;
    input n58827;
    output \data_in_frame[17][7] ;
    output \data_in_frame[17][6] ;
    input n58860;
    input n58861;
    input n58862;
    input n58863;
    input n58864;
    output DE_c;
    output tx_active;
    output LED_c;
    input n58845;
    input n59003;
    input n58865;
    output \data_in_frame[7][7] ;
    output [7:0]\data_in_frame[5] ;
    output \data_out_frame[0][4] ;
    input n59002;
    output \data_in_frame[7][2] ;
    output \data_in_frame[6][7] ;
    input n58866;
    output \data_out_frame[1][0] ;
    input n59001;
    input n28780;
    output \data_in_frame[7][0] ;
    output \data_out_frame[1][1] ;
    input n59000;
    input n58999;
    input n31074;
    input n29319;
    input n31075;
    input n29318;
    input n58998;
    output \data_in_frame[8][4] ;
    output \data_in_frame[7][4] ;
    output \data_in_frame[8][5] ;
    output \data_in_frame[6][3] ;
    output \data_in_frame[7][3] ;
    output \data_in_frame[7][5] ;
    input n30842;
    input n30828;
    output n23230;
    input n30773;
    input n30763;
    input n30761;
    input n30760;
    input n30744;
    input n30742;
    output \data_in_frame[6][1] ;
    input n30710;
    input n30707;
    input n30706;
    input n30705;
    input n30703;
    input n30702;
    input n58296;
    input n29833;
    input n30693;
    input n30690;
    input n58294;
    input n58290;
    input n58286;
    input n58282;
    input n58278;
    input n58274;
    input n58272;
    input n58268;
    input n29861;
    input n58264;
    input n29867;
    input n58260;
    input n30677;
    input n30674;
    input n58256;
    input n30672;
    input n30669;
    input n30664;
    input n30338;
    input n30342;
    input n30348;
    input n30352;
    output \data_in_frame[6][4] ;
    input n30361;
    input n30365;
    input n30368;
    output \data_in_frame[7][1] ;
    input n30371;
    input n30375;
    input n30378;
    input n30381;
    input n30387;
    input n30399;
    output \data_in_frame[8][3] ;
    input n30403;
    input n30639;
    input n30638;
    input n30406;
    input n30409;
    input n30413;
    input n30466;
    input n30469;
    input n30616;
    input n30475;
    input n30479;
    input n30482;
    input n30485;
    input n30489;
    input n30492;
    input n30495;
    input n30499;
    input n58384;
    input n58398;
    input n30509;
    input n30512;
    input n30515;
    input n30550;
    input n30554;
    input n30558;
    input n30562;
    input n30566;
    input n30587;
    input n58252;
    input n58248;
    input n58244;
    output \data_in_frame[20][2] ;
    input n29909;
    output \data_in_frame[20][3] ;
    input n29912;
    output \data_in_frame[20][4] ;
    input n58238;
    input n58234;
    input n58230;
    input n58228;
    input n58226;
    input n58224;
    input n58220;
    input n58216;
    input n58212;
    input n58208;
    input n29949;
    output [7:0]\data_in_frame[22] ;
    input n29952;
    input n58202;
    input n29958;
    input n29961;
    input n29964;
    input n29968;
    input n58198;
    input n30539;
    input n29977;
    output [7:0]\data_in_frame[23] ;
    input n29980;
    input n29983;
    input n29986;
    input n29989;
    input n29992;
    input n29995;
    input n30465;
    input n30003;
    input n30016;
    input n30028;
    input n30031;
    input n30035;
    input n58340;
    input n58997;
    input n58996;
    input n58995;
    input n58994;
    input n58842;
    input n31082;
    input n29317;
    input n58993;
    input n58992;
    input n58991;
    input n58990;
    output \data_in_frame[1][1] ;
    input n58989;
    input n58988;
    output rx_data_ready;
    output n59967;
    input n58867;
    input n58868;
    input n58987;
    input n58986;
    input n58985;
    input n58984;
    input n58869;
    input n58840;
    input n58839;
    input n58983;
    input n58982;
    input n58981;
    input n58870;
    output n42166;
    output n28770;
    input n58871;
    output n59086;
    input n29311;
    input n58872;
    input n58873;
    input n58874;
    input n58875;
    input n58876;
    input n58877;
    input n58878;
    output n8_adj_10;
    output n28725;
    input n58879;
    input n58838;
    input n58880;
    input n58837;
    input n58881;
    input n58882;
    output n8_adj_11;
    output n8_adj_12;
    output n28733;
    input n58980;
    input n58979;
    input n58883;
    input n58978;
    input n58977;
    input n58884;
    input n58885;
    input n58831;
    input n58830;
    input n58886;
    input n58887;
    input n58888;
    input n58889;
    input n58890;
    input n58891;
    input n58892;
    input n58893;
    input n58894;
    input n29283;
    output \data_out_frame[27][6] ;
    output \data_out_frame[26][6] ;
    input n58895;
    input n58824;
    input n31162;
    input n29256;
    input n31163;
    input n29255;
    input n31164;
    input n29254;
    input n58896;
    input n31166;
    input n29251;
    input n58897;
    input n58898;
    input n58828;
    input n58976;
    output n59079;
    input n58975;
    input n58974;
    input n58973;
    input n69908;
    output n28778;
    input n69906;
    input n26087;
    output n59593;
    input n26490;
    output n54003;
    input [23:0]pwm_setpoint;
    output n23164;
    output n44625;
    input n64453;
    input n64451;
    output n59093;
    output n28719;
    output n28723;
    input n35592;
    output n15_adj_13;
    output n54986;
    output n59975;
    output n28791;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    output \o_Rx_DV_N_3617[24] ;
    output [2:0]r_SM_Main;
    output n27;
    input n62584;
    output n28320;
    output n60079;
    output n1;
    output tx_o;
    output [8:0]r_Clock_Count;
    input n30034;
    input n71131;
    input n30847;
    output \r_Bit_Index[0] ;
    output n6;
    output tx_enable;
    output \o_Rx_DV_N_3617[12] ;
    input n5254;
    output \o_Rx_DV_N_3617[8] ;
    output r_Rx_Data;
    output n29;
    output n23;
    output \r_SM_Main[1]_adj_14 ;
    input [31:0]baudrate;
    output n28324;
    output n60053;
    output \r_SM_Main[2]_adj_15 ;
    input RX_N_2;
    output [7:0]r_Clock_Count_adj_25;
    input n30256;
    input n30255;
    input n30254;
    input n30253;
    input n30252;
    output n25975;
    output \o_Rx_DV_N_3617[7] ;
    output \o_Rx_DV_N_3617[6] ;
    output \o_Rx_DV_N_3617[5] ;
    output \o_Rx_DV_N_3617[4] ;
    output \o_Rx_DV_N_3617[3] ;
    output \o_Rx_DV_N_3617[2] ;
    output \o_Rx_DV_N_3617[1] ;
    output \o_Rx_DV_N_3617[0] ;
    output \r_Bit_Index[0]_adj_24 ;
    output n62864;
    input n29921;
    input n59011;
    output n62764;
    output n62780;
    output n62748;
    output n62828;
    output n62812;
    input n30854;
    input n55126;
    input n30850;
    input n5257;
    input n29791;
    output n28127;
    output n62796;
    output n62846;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n30310, n30307, n10_c, n59245, n26, n2, Kp_23__N_741, 
        Kp_23__N_1877, n30167, n2_adj_5401, n30168;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.i_31__N_2636 , n66925, n5, n24, n59127, n29_c, 
        n66932;
    wire [31:0]\FRAME_MATCHER.state_31__N_2741 ;
    
    wire n2_adj_5402, n2_adj_5403, n2_adj_5404, n27_c, n53451, n22, 
        n26786, n31, n30169, n2_adj_5405, n30050, n30170, n2_adj_5406, 
        n2_adj_5407, n30303, n2_adj_5408, n2_adj_5409, n66937, n2_adj_5410, 
        n2_adj_5411, n2_adj_5412, n2_adj_5413, n2_adj_5414, n2_adj_5415, 
        n30200, n67005, n64437, n66938, n64436;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n64438, n70762, n70816, n64392, n64391, n64393, n71086;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n66940;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n30199, n70912, n70822, n69082, n30198, n66943, n70828, 
        n30197, n64058, n30196, n30195, n30194, n30193, n66944, 
        n2_adj_5416, n30192;
    wire [7:0]\data_in_frame[16]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30201, n2_adj_5417, n30300, \FRAME_MATCHER.i_31__N_2643 , 
        n2436, n61096, n4452, n20805, n71065, n71068, n37386, 
        n23149, n4_adj_5418, n28024, n69079, n67088, n71053, n30205, 
        n30297, n30294, n30291, n3303, \FRAME_MATCHER.i_31__N_2641 , 
        n2545, n70774, n7, n30288, n30285;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n30282, n30279, n30276, n30063, n30272, n2439, n2442, 
        n63987, n30269, n61848, n58084, n66945, n2440, n25927, 
        n20798, n2534, n771, \FRAME_MATCHER.i_31__N_2637 , n2533, 
        n5_adj_5419, n66946, n25998, n25869, n27431, n61244, n66947, 
        n25935, n27436;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n10_adj_5420;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n14, n66982, n25950, n20, n25866;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n19, n64191, n67000, n3942, n28716, n26008, n18, n26005, 
        n20_adj_5421, n15_c, n4_adj_5422, n4_adj_5423, n44648, n10_adj_5424, 
        n14_adj_5425, n15_adj_5426, n16, n30203, n17, n30204, n16_adj_5427, 
        n17_adj_5428, n30202, \FRAME_MATCHER.i_31__N_2642 , n59074, 
        n6_c;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [23:0]n5169;
    
    wire n61010, n71150, n30191, n30190, n30189, n30188, n30187, 
        n30186, n30185, n30184, n2_adj_5429, n2_adj_5430;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n30183, n30182, n2_adj_5431, n2_adj_5432, n30181, n2_adj_5433, 
        n2_adj_5434, n2553, n2_adj_5435, n30180, n28140, n30179, 
        n30178, n2_adj_5436, n30177, n2_adj_5437, n30266, n30176, 
        n30263, n2_adj_5438, n2_adj_5439, n30175, n30174, n2_adj_5440, 
        n2_adj_5441, n2_adj_5442, n2_adj_5443, n2_adj_5444, n2_adj_5445, 
        n2_adj_5446, n2_adj_5447, n2_adj_5448, n2_adj_5449, n2_adj_5450, 
        n30173, n30171, n2_adj_5451, n30172, n67090, n67089, n2_adj_5452, 
        n28472, n64419, n64420, n64418, n71116, n70768, n14_adj_5453, 
        n67091, n2_adj_5454, n70972, n69089, n28470, n64416, n64417, 
        n64415, n2_adj_5455, n64568, n2_adj_5456, n64569, n64560, 
        n64559, n64505, n64506, n64512, n2_adj_5457, n64511, n64523, 
        n64524, n2_adj_5458, n64407, n2_adj_5459, n64406, n70852, 
        n66957, n70744, n70780, n69091, n70750, n67132, n64553, 
        n64554, n64563, n64562, n64425, n64426, n64424, n2_adj_5460, 
        n71128, n70720, n14_adj_5461, n70846, n66958, n71122, n70978, 
        n69097, n1_c, n64400, n2_adj_5462, n2_adj_5463, n2_adj_5464, 
        n2_adj_5465, n2_adj_5466, n2_adj_5467, n2_adj_5468, n2_adj_5469, 
        n2_adj_5470, n2_adj_5471, n57, n2_adj_5472, n2_adj_5473, n2_adj_5474, 
        n2_adj_5475;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    
    wire n58298, n70981, n70984, n70975, n70969, n2_adj_5476, n30092, 
        n30095, n30109, n30116, n2_adj_5477, n59517, n54600, n27123, 
        n54920, n59357, Kp_23__N_1004, n59443, n4_adj_5478, n10_adj_5479, 
        n60931, n55033, n59735, n26568, n54732, n61861, n6_adj_5480, 
        n59653, n26806, n5_adj_5481, n61481, n61866, n59711, n26365, 
        n12, n59485, n55007, Kp_23__N_1680, n59341, n59285, n26395, 
        n59331, n59720, n54954, Kp_23__N_1400, n60999, n59461, n59566, 
        n59514, n59107, Kp_23__N_798, n26455, n10_adj_5482, n59392, 
        n54952, n10_adj_5483, n59678, n54914, n14_adj_5484, n33, 
        n54959, n59717, n55098, n59476, n59732, n26447, n59239, 
        n53922, n26389, n59147, n6_adj_5485, n26281, n59657, n10_adj_5486, 
        n10_adj_5487, n54940, n14_adj_5488, n59563, n59110, n59482, 
        n7_adj_5489, n61489, n59553, n54971, n4_adj_5490, n59377;
    wire [7:0]\data_in_frame[17]_c ;   // verilog/coms.v(99[12:25])
    
    wire n10_adj_5491, n59557, n59097, n54016;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    
    wire n59590, n28_adj_5492, n26809, n32, n59773, n54434, n59294, 
        n30, n59174, n53899, n31_adj_5493;
    wire [7:0]\data_in_frame[6]_c ;   // verilog/coms.v(99[12:25])
    
    wire n59281, n59830, n26231, n29_adj_5494, n66899, n2_adj_5495, 
        n66900, n59758, n24160, n59413, n55047, n3, n66901, n2_adj_5498, 
        n66902, n66903, n66904, n66905, n2_adj_5499, n66906, n2_adj_5500, 
        n10_adj_5501, n30166, n30165, n30164, n2_adj_5502, n61452, 
        n59423, n30163, n59755, n2_adj_5503, n2_adj_5504, n2_adj_5505, 
        n2_adj_5506, n30162, n2_adj_5507, n30161, n26598, n6_adj_5508, 
        n60966, n10_adj_5509, n30160, n59821, n30159, n30158, n59729, 
        n42, n2_adj_5510, n58816, n51498, n58814, n58817, n51497, 
        n30157, n2_adj_5511, n2_adj_5512, n30156, n30155, n30154, 
        n2_adj_5513, n2_adj_5514, n2_adj_5515, n30153, n2_adj_5516, 
        n30152, n66907, n30151, n30150, n30149, n2_adj_5517, n2_adj_5518, 
        n2_adj_5519, n30148, n66908, n30147, n30146, n2_adj_5520, 
        n59827, n8_adj_5521, n66909, n2_adj_5522, n30145, n2_adj_5523, 
        n2_adj_5524, n2_adj_5525, n30144, n66912, n59746, n59749, 
        n54411, n12_adj_5526, n66913, n30143, n30142, n30141, n30140, 
        n30139, n30138, n30137, n66917, n66918, n57_adj_5527, n66919, 
        n30136, n30135, n30134, n30133, n55066, n66, n26376, n64, 
        n2_adj_5528, n2_adj_5529, n30132, n30131, n2_adj_5530, Kp_23__N_1518, 
        n38, n65, n2_adj_5531, n58818, n51496, n2_adj_5532, n2_adj_5533, 
        n66921, n3_adj_5534, n30122, n30120, n66922, n26197, n63, 
        n30119, n30115, n2_adj_5535, n2_adj_5536, n30112, n2_adj_5537, 
        n2_adj_5538, n30108, n30107, n30106, n2_adj_5539, n30105, 
        n2_adj_5540, n2_adj_5541, n44, n58819, n51495, n54900, n59824, 
        n59493, n27228, n62, n59818, n61, n72, n59488, n60_adj_5542, 
        n59338, n67, n54957, n59464, n30101, n59309, n54397, n59507, 
        n10_adj_5543, n24389, n26134, n26878, n26189, n6_adj_5544, 
        n59242;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    
    wire n59545, n24393, n59762, n54440, n54943, n61148, n3_adj_5545, 
        Kp_23__N_1214, n59504, n30089, n30088, n30087, n30086, n30085, 
        n30084, n30083, n30082, n30081, n30080, n30079, n27255, 
        n26316, n59699, n30078, n30077, n30076;
    wire [7:0]\data_in_frame[8]_c ;   // verilog/coms.v(99[12:25])
    
    wire n58444, n59578, n6_adj_5546, n30393, tx_transmit_N_3545, 
        \FRAME_MATCHER.i_31__N_2640 , n1_adj_5547, n58438;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n30646, n54659, n26687, n6_adj_5548, n64526, n64527, n70909, 
        n25, n64503, n64502, n33_adj_5549, n2_adj_5550, n38_adj_5551, 
        n27142, n36, n58434, n58428, n58446, n59522, n55073, n4_adj_5552, 
        n54896, n69904, n71077, n30071, n30070, n30069, n54694, 
        n3_adj_5553, n30027, n30011, n30009, n30008, n2_adj_5554, 
        n30007, n30006, n30002, n29998, n2_adj_5555, n2_adj_5556, 
        n2_adj_5557, n2_adj_5558, n2_adj_5559, n2_adj_5560, n2_adj_5561, 
        n2_adj_5562, n2_adj_5563, n2_adj_5564, n2_adj_5565, n2_adj_5566, 
        n2_adj_5567, n2_adj_5568, n2_adj_5569, n2_adj_5570, n2_adj_5571, 
        n2_adj_5572, n2_adj_5573, n2_adj_5574, n2_adj_5575, n2_adj_5576, 
        n2_adj_5577, n2_adj_5578, n2_adj_5579, n2_adj_5580, n2_adj_5581, 
        n2_adj_5582, n64493, n64494, n70903, n54030, n22_adj_5583, 
        n37, n58820, n51494, n59638, n35, n2_adj_5584, n26719, 
        n59714, n59446, n12_adj_5585, n59741, n8_adj_5586, n10_adj_5587, 
        n59524, n59726, n12_adj_5588, n2_adj_5589, n58821, n51493, 
        n2_adj_5590, n16_adj_5591, n6_adj_5592, n28405, n59171, Kp_23__N_1007, 
        n59276, n10_adj_5593, n26357, n59650, n26296, n6_adj_5594, 
        n59764, n2_adj_5595, n2_adj_5596, n2_adj_5597, n2_adj_5598, 
        n28407, n28409, n28411, n28413, n28415, n28417, n28419, 
        n28421, n28423, n28425, n28427, n28429, n28431, n28433, 
        n28435, n28437, n28439, n28441, n28443, n28445, n28447, 
        n28449, n28451, n28453, n28455, n28457, n28459, n28461, 
        n28463, n28465, n28467, n2_adj_5599, n2_adj_5600, n2_adj_5601, 
        n59300, n6_adj_5602, n59060, n27340;
    wire [2:0]r_SM_Main_2__N_3674;
    
    wire n2_adj_5603, Kp_23__N_1209, n8_adj_5604, n12_adj_5605, n59395, 
        n59191, n10_adj_5606, n16_adj_5607, n59312, LED_N_3537, LED_N_3536, 
        n27759, n29263, n59799, n54912, n15_adj_5608, n14_adj_5609, 
        n6_adj_5610, n60988, n53918, n3_adj_5611, n58822, n51492, 
        n55118, n2_adj_5612, n59510, n25579, n59533, n5_adj_5613, 
        n2_adj_5614, n2_adj_5615, n24221, n59569, n53905, n59632, 
        n59212, n12_adj_5616, n2_adj_5617, n8_adj_5618, n59644, n64509, 
        n64508, n70906, n26707, n2_adj_5619, n2_adj_5620, n58184, 
        n26844, n59573, n59130, n55014, n59141, n54996, n18_adj_5621, 
        n2_adj_5622, n2_adj_5623, n26753, n2_adj_5624, n54889, n61790, 
        n59723, n20_adj_5625, n28_adj_5626, n4_adj_5627, n15_adj_5628, 
        n61719, n26756, n6_adj_5629, n2_adj_5630, n2_adj_5631, n26330, 
        Kp_23__N_1001, Kp_23__N_998, n26173, n26333, n59420, n59365, 
        n2329, n3_adj_5632, Kp_23__N_901, n26339, n6_adj_5633, n61557, 
        n59796, n27074, n26760, n29785, n59264, n30858, n59479, 
        n59839, n10_adj_5634, n29788, n6_adj_5635, n59681, n26617, 
        n12_adj_5636, n29792, n29795, n29798, n29801, n29804, n29807, 
        n29810, n59407, n53959, n59602, n59315, n3_adj_5637, n29815, 
        n29818, n30313, Kp_23__N_928, n6_adj_5638, n30745, n29821, 
        n30741, n53944, n30740, n30739, n30738, n30737, n30736, 
        n30735, n30734, n30733, n30732, n30731, n30730, n30729, 
        n30728, n30727, n30726, n30725, n30724, n30723, n30722, 
        n30721, n6_adj_5639, n30720, n30719, n30718, n30717, n30716, 
        n30715, n30714, n30713, n30712, n30711, n29824, n30316, 
        n30699, n6_adj_5640, n30319, n30322, n30326, n3_adj_5641, 
        n59251, n29876, n29879, n29882, n29885, n30329, n30332, 
        n30335, n30416, n26848, n59527, n59705, n12_adj_5642, n26302, 
        n30419, n30422, n30425, n30428, n30431, n30434, n8_adj_5643, 
        n3_adj_5644, n30437, n30440, n58460, n30446, n30449, n30453, 
        n30456, n30459, n30462, n30519, n30522, n30525, n30529, 
        n30532, n30536, n30541, n30545, n29888, n29891, n29894, 
        n29897, n59805, n59144, n10_adj_5645, n6_adj_5646, n59473, 
        n3_adj_5647, n59585, n59165, n27181, n59354, n59672, n26750, 
        n59291, n18_adj_5648, n30_adj_5649, n6_adj_5650, n59560, Kp_23__N_877, 
        n28_adj_5651, n29_adj_5652, n27_adj_5653, n59273, n54966, 
        n61480, n30019;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    
    wire n59470, n59104, n61255, n59205, n26123, n59539, n14_adj_5654, 
        n59168, n13, n7_adj_5655, n64209, n27305, n14_adj_5656, 
        n59761, n64242, n28_adj_5657, n29_adj_5658, n59363, n13_adj_5659, 
        n7_adj_5660, n27_adj_5661, n10_adj_5662, n55120, n20_adj_5663, 
        n59440, n13_adj_5664, n59845, n22_adj_5665, n59542, n21, 
        n59842, n61385, n59814, n59583, n10_adj_5666, n59647, n10_adj_5667, 
        n59744, n55038, n3_adj_5668, n61318, n61138, n14_adj_5669, 
        n59437, n15_adj_5670, n10_adj_5671, n61218, n59449, n54753, 
        n59383, n59660, n26523, n30043, n23_c, n14_adj_5672, n13_adj_5673, 
        n60916, n18_adj_5674, n64044, n61145, n29_adj_5675, n8_adj_5676, 
        n7_adj_5677, n64048, n61289, n22_adj_5678, n64046, n61159, 
        n32_adj_5679, n27_adj_5680, n44_adj_5681, n26113, n59404, 
        n54669, n59416, n42_adj_5682, n43, n41, n40, n39, n50, 
        n45, n6_adj_5683, n59547, n3_adj_5684, n61040, n26237, n59371, 
        n59254, n25546, n68989, n66942, n70879, n70792, n7_adj_5685, 
        n4_adj_5686, n5_adj_5687, n70873, n67007, n67006, n70876, 
        n70867, n64401, n2_adj_5688, n59693, n59431, n54945, n10_adj_5689, 
        n2_adj_5690, n59083, n2_adj_5691, n2_adj_5692, n2_adj_5693, 
        n2_adj_5694, n2_adj_5695, n2_adj_5696, n7_adj_5697, n2_adj_5698, 
        n2_adj_5699, n28480, n2_adj_5701, n2_adj_5702, n64449, n2_adj_5703, 
        n64450, n2_adj_5704, n2_adj_5705, n64448, n2_adj_5706, n58815, 
        n2_adj_5709, n2_adj_5710, n2_adj_5711, n2_adj_5712, n2_adj_5713, 
        n2_adj_5714, n2_adj_5715, n10_adj_5716, n70756, n53903, n14_adj_5717, 
        n2_adj_5718, n2_adj_5719, n2_adj_5720, n2_adj_5721, n2_adj_5722, 
        n59550, n2_adj_5723, n2_adj_5724, n2_adj_5725, n2_adj_5726, 
        n2_adj_5727, n2_adj_5728, n2_adj_5729, n1_adj_5730, n1_adj_5731, 
        n1_adj_5732, n1_adj_5733, n1_adj_5734, n1_adj_5735, n1_adj_5736, 
        n3_adj_5737;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n58798, n3_adj_5738, n58799, n3_adj_5739, n58800, n3_adj_5740, 
        n58796, n3_adj_5741, n58801, n58802, n58803, n58804;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n58805, n58806, n58807, n58797, n29261, n58808, n29241, 
        n70732, n58809, n59077, n1_adj_5742, n58810, n58795, n7_adj_5743, 
        n26970, n59318, n25517, n6_adj_5744, n52702, n52701, n52700, 
        n52699, n52698, n52697, n52696, n52695, n52694, n52693, 
        n52692, n52691, n52690, n66924, n52689, n52688, n59833, 
        n59185, n10_adj_5745, n52687, n52686, n52685, n52684, n52683, 
        n52682, n26094, n6_adj_5746, n61754, n52681, n59690, n18_adj_5747, 
        n54222, n16_adj_5748, n20_adj_5749, n52680, n70855, n55026, 
        n70858, n70849, n52679, n52678, n52677, n52676, n52675, 
        n52674, n52673, n52672;
    wire [31:0]n133;
    
    wire n161, n6_adj_5750, n54991, n6_adj_5751, n59121, n59225, 
        n54962, n59663, n10_adj_5752, n54916, n59360, n54161, n42164, 
        n59100, n26509, n59261, n54982, n59361, n59784, n30_adj_5753, 
        n34, n59811, n59635, n32_adj_5754, n33_adj_5755, n26137, 
        n31_adj_5756, n59625, n6_adj_5757, n10_adj_5758, n10_adj_5759, 
        n1519, n1516, n59347, n10_adj_5760, n54734, n59157, n43937, 
        n59235, n59196, n59150, n22_adj_5761, n54994, n16_adj_5762, 
        n24_adj_5763, n70843, n1312, n26693, n20_adj_5764, n59606, 
        n59455, n59629, n59114, n54935, n59368, n26651, n59675, 
        n59641, n26504, n54383, n59793, n54908, n6_adj_5765, n10_adj_5766, 
        n6_adj_5767, n59458, n59188, n10_adj_5768, n59598, n59708, 
        n59781, n54750, n59616, n59619, n59767, n10_adj_5769, n54698, 
        n59270, n27113, n53893, n59808, n11_adj_5770, n59776, n27029, 
        n13_adj_5771, n10_adj_5772, n59222, n32_adj_5773, n61823, 
        n59162, n6_adj_5774, n59669, n6_adj_5775, n61686, n59327, 
        n59401, n1835, n1130, n26660, n12_adj_5776, n59350, n10_adj_5777, 
        n59267, n24_adj_5778, n59154, n26_adj_5779, n59202, n25_adj_5780, 
        n59181, n26516, n14_adj_5781, n27_adj_5782, n9, n6_adj_5783, 
        n1191, n14_adj_5784, n59666, n14_adj_5785, n13_adj_5786, n27086, 
        n59218, n26768, n10_adj_5787, n59153, n59344, n26681, n59324, 
        n14_adj_5788, n15_adj_5789, n44_adj_5790, n59836, n42_adj_5791, 
        n43_adj_5792, n41_adj_5793, n40_adj_5794, n45_adj_5795, n50_adj_5796, 
        n49, n59374, n59610, n8_adj_5797, n7_adj_5798, n59118, n59047, 
        n64549, n59232, n12_adj_5799, n12_adj_5800, n7_adj_5801, n7_adj_5802, 
        n7_adj_5803, n8_adj_5804, n26954, n14_adj_5805, n12_adj_5806, 
        n70837, n70840, n28745, n59790, n59398, n59613, n70831, 
        n59787, n70834, n22_adj_5807, n70714, n70825, n23_adj_5808, 
        n71125, n59687, n71119, n10_adj_5810, n70819, n59410, n71113, 
        n70813, n71107, n70807, n70810, n71101, n70786, n70795, 
        n71095, n70798, n70789, n70783, n70777, n70771, n70765, 
        n70759, n70753, n70747, n70741, n70729, n70723, n70726, 
        n70717, n70711, n71089, n6_adj_5811, n5_adj_5812, n6_adj_5813, 
        n7_adj_5814, n59135, n71083, n62490;
    wire [2:0]r_SM_Main_2__N_3665;
    
    wire n60937, n60609;
    
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30310));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30307));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut (.I0(\data_in_frame[2] [0]), .I1(n10_c), .I2(n59245), 
            .I3(\data_in_frame[1] [5]), .O(n26));
    defparam i9_4_lut.LUT_INIT = 16'h2100;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2), .S(n58972));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15760_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n30167));
    defparam i15760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5401), .S(n58971));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15761_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n30168));
    defparam i15761_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51373_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66925));   // verilog/coms.v(158[12:15])
    defparam i51373_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(n5), .I1(n24), .I2(\data_in_frame[0] [7]), 
            .I3(n59127), .O(n29_c));
    defparam i12_4_lut.LUT_INIT = 16'h0440;
    SB_LUT4 i51846_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66932));   // verilog/coms.v(158[12:15])
    defparam i51846_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_810_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5403), .S(n58970));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_4_lut (.I0(n27_c), .I1(n53451), .I2(n22), .I3(n26786), 
            .O(n31));
    defparam i14_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i15762_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n30169));
    defparam i15762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5405), .S(n58969));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
           .D(n30050));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15763_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n30170));
    defparam i15763_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_810_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[5] [1]), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30303));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1108 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[5] [0]), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1108.LUT_INIT = 16'ha088;
    SB_LUT4 select_810_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51096_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66937));   // verilog/coms.v(158[12:15])
    defparam i51096_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_810_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15793_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n30200));
    defparam i15793_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51153_2_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67005));
    defparam i51153_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i48263_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64437));
    defparam i48263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51099_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66938));   // verilog/coms.v(158[12:15])
    defparam i51099_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48262_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64436));
    defparam i48262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48264_4_lut (.I0(n64437), .I1(n67005), .I2(byte_transmit_counter_c[4]), 
            .I3(\byte_transmit_counter[1] ), .O(n64438));
    defparam i48264_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i48218_3_lut (.I0(n70762), .I1(n70816), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n64392));
    defparam i48218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48217_4_lut (.I0(n64438), .I1(n64436), .I2(byte_transmit_counter_c[4]), 
            .I3(\byte_transmit_counter[1] ), .O(n64391));
    defparam i48217_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i48219_3_lut (.I0(n64391), .I1(n64392), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n64393));
    defparam i48219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(n64393), .I1(n71086), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(tx_data[2]));   // verilog/coms.v(105[12:33])
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51105_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66940));   // verilog/coms.v(158[12:15])
    defparam i51105_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15792_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n30199));
    defparam i15792_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i52907_4_lut (.I0(n70912), .I1(n70822), .I2(byte_transmit_counter_c[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n69082));
    defparam i52907_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i21864_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n30198));
    defparam i21864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51208_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66943));   // verilog/coms.v(158[12:15])
    defparam i51208_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48399_3_lut (.I0(n70828), .I1(n69082), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i48399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15790_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n30197));
    defparam i15790_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut (.I0(n31), .I1(n29_c), .I2(n64058), .I3(n26), 
            .O(\FRAME_MATCHER.state_31__N_2741 [3]));
    defparam i16_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i15789_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n30196));
    defparam i15789_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15788_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n30195));
    defparam i15788_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15787_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n30194));
    defparam i15787_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23004_3_lut (.I0(n28), .I1(n379), .I2(n405), .I3(GND_net), 
            .O(n4));
    defparam i23004_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i15786_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n30193));
    defparam i15786_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51116_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66944));   // verilog/coms.v(158[12:15])
    defparam i51116_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_810_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15785_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n30192));
    defparam i15785_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15794_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [6]), 
            .I3(deadband[6]), .O(n30201));
    defparam i15794_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_810_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30300));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6726_4_lut (.I0(\FRAME_MATCHER.i_31__N_2643 ), .I1(n2436), 
            .I2(n61096), .I3(n4452), .O(n20805));   // verilog/coms.v(148[4] 304[11])
    defparam i6726_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54834 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n71065));
    defparam byte_transmit_counter_0__bdd_4_lut_54834.LUT_INIT = 16'he4aa;
    SB_LUT4 n71065_bdd_4_lut (.I0(n71065), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n71068));
    defparam n71065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i23026_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [1]), 
            .I3(deadband[1]), .O(n37386));
    defparam i23026_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1109 (.I0(n20805), .I1(n2436), .I2(n23149), .I3(n4_adj_5418), 
            .O(n28024));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1109.LUT_INIT = 16'hbbba;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54839 (.I0(byte_transmit_counter_c[3]), 
            .I1(n69079), .I2(n67088), .I3(byte_transmit_counter_c[4]), 
            .O(n71053));
    defparam byte_transmit_counter_3__bdd_4_lut_54839.LUT_INIT = 16'he4aa;
    SB_LUT4 i15798_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [2]), 
            .I3(deadband[2]), .O(n30205));
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30294));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30291));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i495_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2641 ), .I2(GND_net), 
            .I3(GND_net), .O(n2545));   // verilog/coms.v(148[4] 304[11])
    defparam i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71053_bdd_4_lut (.I0(n71053), .I1(n70774), .I2(n7), .I3(byte_transmit_counter_c[4]), 
            .O(tx_data[1]));
    defparam n71053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30285));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30282));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30279));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30276));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
           .D(n30063));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30272));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47824_4_lut (.I0(n2436), .I1(n2439), .I2(n3303), .I3(n2442), 
            .O(n63987));   // verilog/coms.v(139[4] 141[7])
    defparam i47824_4_lut.LUT_INIT = 16'h0a02;
    SB_DFFE data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30269));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1110 (.I0(\FRAME_MATCHER.i_31__N_2641 ), .I1(n2439), 
            .I2(n63987), .I3(n61848), .O(n58084));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1110.LUT_INIT = 16'hb3a0;
    SB_LUT4 i51117_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66945));   // verilog/coms.v(158[12:15])
    defparam i51117_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6719_4_lut (.I0(n2440), .I1(\FRAME_MATCHER.state[3] ), .I2(n2442), 
            .I3(n25927), .O(n20798));   // verilog/coms.v(148[4] 304[11])
    defparam i6719_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i484_2_lut (.I0(\FRAME_MATCHER.state_31__N_2741 [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(GND_net), .I3(GND_net), .O(n2534));   // verilog/coms.v(148[4] 304[11])
    defparam i484_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i483_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2637 ), .I2(GND_net), 
            .I3(GND_net), .O(n2533));   // verilog/coms.v(148[4] 304[11])
    defparam i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29739_4_lut (.I0(n5_adj_5419), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i29739_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i51118_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66946));   // verilog/coms.v(158[12:15])
    defparam i51118_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(n25998), .I2(GND_net), 
            .I3(GND_net), .O(n25869));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29741_4_lut (.I0(n8), .I1(\FRAME_MATCHER.i [31]), .I2(n25869), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i29741_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2641 ), .I2(GND_net), 
            .I3(GND_net), .O(n23149));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_2_lut (.I0(n25927), .I1(\FRAME_MATCHER.i_31__N_2636 ), .I2(GND_net), 
            .I3(GND_net), .O(n27431));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(n4452), .I1(n27431), .I2(\FRAME_MATCHER.i_31__N_2643 ), 
            .I3(n23149), .O(n61244));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i51119_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66947));   // verilog/coms.v(158[12:15])
    defparam i51119_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1111 (.I0(n25935), .I1(n2442), .I2(n2440), .I3(n61244), 
            .O(n27436));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1111.LUT_INIT = 16'hbaaa;
    SB_LUT4 i2_2_lut_adj_1112 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5420));
    defparam i2_2_lut_adj_1112.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), .I2(\data_in[3] [1]), 
            .I3(\data_in[0] [7]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51021_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66982));   // verilog/coms.v(158[12:15])
    defparam i51021_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut (.I0(\data_in[3] [6]), .I1(n14), .I2(n10_adj_5420), 
            .I3(\data_in[2] [1]), .O(n25950));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), .I2(n25950), 
            .I3(\data_in[0] [5]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1113 (.I0(n25866), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19));
    defparam i7_4_lut_adj_1113.LUT_INIT = 16'hfeff;
    SB_LUT4 i48026_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [3]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n64191));
    defparam i48026_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i51173_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n67000));   // verilog/coms.v(158[12:15])
    defparam i51173_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14310_1_lut (.I0(n3942), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28716));   // verilog/coms.v(148[4] 304[11])
    defparam i14310_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_3_lut (.I0(n64191), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n2436));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1114 (.I0(\data_in[2] [4]), .I1(n25950), .I2(\data_in[1] [5]), 
            .I3(n26008), .O(n18));
    defparam i7_4_lut_adj_1114.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1115 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n26005), .O(n20_adj_5421));
    defparam i9_4_lut_adj_1115.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_c));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_c), .I1(n20_adj_5421), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n2439));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5422));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter[0]), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[1] ), 
            .O(n4_adj_5423));
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'ha8a0;
    SB_LUT4 i30348_4_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5423), .I3(n4_adj_5422), .O(n44648));
    defparam i30348_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i4_4_lut (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [4]), .O(n10_adj_5424));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut (.I0(\data_in[3] [4]), .I1(n10_adj_5424), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n26008));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i5_3_lut_adj_1118 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5425));
    defparam i5_3_lut_adj_1118.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1119 (.I0(\data_in[0] [6]), .I1(n26008), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5426));
    defparam i6_4_lut_adj_1119.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1120 (.I0(n15_adj_5426), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5425), .I3(\data_in[0] [3]), .O(n25866));
    defparam i8_4_lut_adj_1120.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1121 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut_adj_1121.LUT_INIT = 16'hfffe;
    SB_LUT4 i15796_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [4]), 
            .I3(deadband[4]), .O(n30203));
    defparam i15796_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1122 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_1122.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1123 (.I0(n17), .I1(\data_in[1] [6]), .I2(n16), 
            .I3(\data_in[3] [7]), .O(n26005));
    defparam i9_4_lut_adj_1123.LUT_INIT = 16'hfbff;
    SB_LUT4 i15797_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [3]), 
            .I3(deadband[3]), .O(n30204));
    defparam i15797_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1124 (.I0(n26005), .I1(\data_in[3] [3]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_5427));
    defparam i6_4_lut_adj_1124.LUT_INIT = 16'hffbf;
    SB_LUT4 i7_4_lut_adj_1125 (.I0(\data_in[2] [3]), .I1(n25866), .I2(\data_in[3] [5]), 
            .I3(\data_in[0] [7]), .O(n17_adj_5428));
    defparam i7_4_lut_adj_1125.LUT_INIT = 16'hffdf;
    SB_LUT4 i15795_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [5]), 
            .I3(deadband[5]), .O(n30202));
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_4_lut_adj_1126 (.I0(n17_adj_5428), .I1(\data_in[0] [2]), 
            .I2(n16_adj_5427), .I3(\data_in[3] [1]), .O(n2442));
    defparam i9_4_lut_adj_1126.LUT_INIT = 16'hfbff;
    SB_LUT4 i401_2_lut (.I0(n2439), .I1(n2436), .I2(GND_net), .I3(GND_net), 
            .O(n2440));   // verilog/coms.v(142[4] 144[7])
    defparam i401_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\FRAME_MATCHER.i_31__N_2642 ), .I1(Kp_23__N_1877), 
            .I2(GND_net), .I3(GND_net), .O(n59074));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1128 (.I0(n59074), .I1(n2440), .I2(n2442), .I3(\FRAME_MATCHER.i_31__N_2636 ), 
            .O(n6_c));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1128.LUT_INIT = 16'heaaa;
    SB_LUT4 mux_1084_i1_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n5169[0]));
    defparam mux_1084_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i3_4_lut (.I0(n61010), .I1(n6_c), .I2(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2638 ), .O(n71150));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut.LUT_INIT = 16'hefee;
    SB_LUT4 i15784_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n30191));
    defparam i15784_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15783_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n30190));
    defparam i15783_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15782_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n30189));
    defparam i15782_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15781_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n30188));
    defparam i15781_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15780_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n30187));
    defparam i15780_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15779_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n30186));
    defparam i15779_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15778_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n30185));
    defparam i15778_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15777_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n30184));
    defparam i15777_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5429), .S(n58968));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5430), .S(n58967));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15776_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n30183));
    defparam i15776_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15775_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n30182));
    defparam i15775_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5431), .S(n58966));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5432), .S(n58965));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15774_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n30181));
    defparam i15774_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5433), .S(n59004));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5434), .S(n58964));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1877), .C(clk16MHz), 
            .D(n2553), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 select_810_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15773_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n30180));
    defparam i15773_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n28140), 
            .D(n5169[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i21865_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n30179));
    defparam i21865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15771_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n30178));
    defparam i15771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_810_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), .O(n2_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15770_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n30177));
    defparam i15770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_810_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30266));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15769_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n30176));
    defparam i15769_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30263));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5438), .S(n58963));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5439), .S(n58962));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15768_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n30175));
    defparam i15768_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15767_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n30174));
    defparam i15767_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5440), .S(n58961));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5441), .S(n58960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5442), .S(n58959));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5443), .S(n58958));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5444), .S(n58957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5445), .S(n58825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5446), .S(n58956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5447), .S(n58955));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5448), .S(n58954));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5449), .S(n58953));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5450), .S(n58952));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22309_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n30173));
    defparam i22309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15764_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n30171));
    defparam i15764_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5451), .S(n58951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30260));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i22310_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n30172));
    defparam i22310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30257));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23_2_lut (.I0(n149), .I1(IntegralLimit[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(248[22:35])
    defparam i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51425_4_lut (.I0(\data_out_frame[12] [2]), .I1(byte_transmit_counter_c[4]), 
            .I2(\data_out_frame[13] [2]), .I3(byte_transmit_counter[0]), 
            .O(n67090));
    defparam i51425_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51234_4_lut (.I0(\data_out_frame[14] [2]), .I1(byte_transmit_counter_c[4]), 
            .I2(\data_out_frame[15] [2]), .I3(byte_transmit_counter[0]), 
            .O(n67089));
    defparam i51234_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 select_810_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14066_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28472));   // verilog/coms.v(109[34:55])
    defparam i14066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48245_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64419));
    defparam i48245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48246_4_lut (.I0(n64419), .I1(n28472), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n64420));
    defparam i48246_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48244_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64418));
    defparam i48244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30768125_i1_3_lut (.I0(n71116), .I1(n70768), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5453));
    defparam i30768125_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51424_2_lut (.I0(n70864), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67091));
    defparam i51424_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_810_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i52914_3_lut (.I0(n71068), .I1(n70972), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69089));
    defparam i52914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14064_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28470));   // verilog/coms.v(109[34:55])
    defparam i14064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48242_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64416));
    defparam i48242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48243_4_lut (.I0(n64416), .I1(n28470), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n64417));
    defparam i48243_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48241_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64415));
    defparam i48241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .I2(\data_out_frame[3][4] ), .I3(GND_net), .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i48394_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64568));
    defparam i48394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i48395_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64569));
    defparam i48395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48386_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64560));
    defparam i48386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48385_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64559));
    defparam i48385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48331_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64505));
    defparam i48331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48332_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64506));
    defparam i48332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48338_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64512));
    defparam i48338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i48337_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64511));
    defparam i48337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48349_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64523));
    defparam i48349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48350_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64524));
    defparam i48350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i48233_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64407));
    defparam i48233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i48232_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64406));
    defparam i48232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51123_2_lut (.I0(n70852), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66957));
    defparam i51123_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i52916_3_lut (.I0(n70744), .I1(n70780), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69091));
    defparam i52916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51248_2_lut (.I0(n70750), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67132));
    defparam i51248_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48379_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64553));
    defparam i48379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48380_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64554));
    defparam i48380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48389_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64563));
    defparam i48389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48388_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64562));
    defparam i48388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48251_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64425));
    defparam i48251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48252_4_lut (.I0(n64425), .I1(n28507), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][5] ), .O(n64426));
    defparam i48252_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i48250_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64424));
    defparam i48250_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5460), .S(n58950));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i30756119_i1_3_lut (.I0(n71128), .I1(n70720), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_5461));
    defparam i30756119_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51221_2_lut (.I0(n70846), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66958));
    defparam i51221_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i52922_3_lut (.I0(n71122), .I1(n70978), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69097));
    defparam i52922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_c));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48226_4_lut (.I0(n1_c), .I1(\data_out_frame[3][3] ), .I2(\byte_transmit_counter[1] ), 
            .I3(byte_transmit_counter[0]), .O(n64400));
    defparam i48226_4_lut.LUT_INIT = 16'hca0a;
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5462), .S(n58949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5463), .S(n58948));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5464), .S(n58947));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5465), .S(n58946));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5466), .S(n58945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5467), .S(n58944));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5468), .S(n58943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5469), .S(n58942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5470), .S(n58941));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5471), .S(n58940));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut (.I0(n3942), .I1(n60), .I2(n57), .I3(GND_net), 
            .O(n51));
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5472), .S(n58939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5473), .S(n58938));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5474), .S(n58937));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5475), .S(n58936));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut_adj_1129 (.I0(\data_in_frame[20] [6]), .I1(n28717), 
            .I2(n28774), .I3(rx_data[6]), .O(n58298));
    defparam i12_4_lut_adj_1129.LUT_INIT = 16'h3a0a;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54824 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70981));
    defparam byte_transmit_counter_0__bdd_4_lut_54824.LUT_INIT = 16'he4aa;
    SB_LUT4 n70981_bdd_4_lut (.I0(n70981), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70984));
    defparam n70981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54754 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n70975));
    defparam byte_transmit_counter_0__bdd_4_lut_54754.LUT_INIT = 16'he4aa;
    SB_LUT4 n70975_bdd_4_lut (.I0(n70975), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n70978));
    defparam n70975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54749 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n70969));
    defparam byte_transmit_counter_0__bdd_4_lut_54749.LUT_INIT = 16'he4aa;
    SB_LUT4 n70969_bdd_4_lut (.I0(n70969), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n70972));
    defparam n70969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30228));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30225));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5476), .S(n58935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30222));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30219));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30216));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n30092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n30095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n30109));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n30116));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30208));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n30207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n37386), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n30205), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n30204), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n30203), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n30202), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1130 (.I0(\data_in_frame[18] [0]), .I1(n59517), 
            .I2(n54600), .I3(n27123), .O(n54920));
    defparam i3_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n30201), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[4] [2]), .I1(n59357), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[1] [6]), .O(Kp_23__N_1004));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n30200), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1131 (.I0(n59443), .I1(\data_in_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5478));
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1132 (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[21] [0]), 
            .I2(\data_in_frame[18] [6]), .I3(\data_in_frame[20][7] ), .O(n10_adj_5479));
    defparam i4_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n60931), .I1(n10_adj_5479), .I2(n55033), .I3(n4_adj_5478), 
            .O(n59735));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1133 (.I0(n26568), .I1(n54732), .I2(\data_in_frame[19] [4]), 
            .I3(GND_net), .O(n61861));
    defparam i2_3_lut_adj_1133.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5480));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1135 (.I0(n59653), .I1(n26806), .I2(n5_adj_5481), 
            .I3(n6_adj_5480), .O(n61481));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1136 (.I0(\data_in_frame[15] [3]), .I1(n61866), 
            .I2(n59711), .I3(n26365), .O(n12));
    defparam i5_4_lut_adj_1136.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1137 (.I0(n59485), .I1(n12), .I2(n61481), .I3(\data_in_frame[17] [5]), 
            .O(n54600));
    defparam i6_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(n55007), .I1(n54600), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1680));
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1139 (.I0(\data_in_frame[20][1] ), .I1(n59341), 
            .I2(\data_in_frame[18] [1]), .I3(GND_net), .O(n59285));
    defparam i2_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1140 (.I0(\data_in_frame[16]_c [2]), .I1(n26395), 
            .I2(\data_in_frame[14] [0]), .I3(n59331), .O(n59720));
    defparam i3_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1141 (.I0(\data_in_frame[16]_c [3]), .I1(n59720), 
            .I2(n54954), .I3(Kp_23__N_1400), .O(n60931));
    defparam i3_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(n60931), .I1(n60999), .I2(GND_net), 
            .I3(GND_net), .O(n27123));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(n27123), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[20][5] ), .I3(\data_in_frame[18] [4]), .O(n59461));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1144 (.I0(\data_in_frame[16]_c [3]), .I1(n59566), 
            .I2(\data_in_frame[18] [5]), .I3(\data_in_frame[20][7] ), .O(n59514));
    defparam i3_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[8] [6]), .I1(n59107), 
            .I2(GND_net), .I3(GND_net), .O(n26806));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1146 (.I0(n59711), .I1(Kp_23__N_798), .I2(n26455), 
            .I3(n5_adj_5481), .O(n10_adj_5482));
    defparam i4_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1147 (.I0(\data_in_frame[15] [3]), .I1(n59392), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n55007));
    defparam i2_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1148 (.I0(n59392), .I1(n54952), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5483));
    defparam i2_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1149 (.I0(n59678), .I1(n54914), .I2(Kp_23__N_1400), 
            .I3(\data_in_frame[14] [7]), .O(n14_adj_5484));
    defparam i6_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1150 (.I0(\data_in_frame[17] [3]), .I1(n14_adj_5484), 
            .I2(n10_adj_5483), .I3(n33), .O(n26568));
    defparam i7_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[17] [1]), .I1(n54732), 
            .I2(GND_net), .I3(GND_net), .O(n54959));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1152 (.I0(\data_in_frame[21] [5]), .I1(n25605), 
            .I2(n54959), .I3(\data_in_frame[19] [3]), .O(n59717));
    defparam i1_4_lut_adj_1152.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(n26568), .I1(n55007), .I2(GND_net), 
            .I3(GND_net), .O(n55098));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1154 (.I0(n55098), .I1(n59717), .I2(\data_in_frame[19] [5]), 
            .I3(\data_in_frame[21] [6]), .O(n59476));
    defparam i3_4_lut_adj_1154.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1155 (.I0(\data_in_frame[16]_c [6]), .I1(\data_in_frame[16]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59732));
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[14] [7]), .I3(n59653), .O(n59499));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1400));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(n26447), .I1(n59239), .I2(\data_in_frame[13] [0]), 
            .I3(GND_net), .O(n53922));
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1158 (.I0(n26389), .I1(\data_in_frame[13] [2]), 
            .I2(n59147), .I3(n6_adj_5485), .O(n59239));   // verilog/coms.v(88[17:63])
    defparam i4_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1159 (.I0(n59239), .I1(n53922), .I2(n26281), 
            .I3(n59657), .O(n10_adj_5486));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1160 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(n10_adj_5486), .I3(\data_in_frame[14] [7]), .O(n10_adj_5487));
    defparam i2_4_lut_adj_1160.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1161 (.I0(n59499), .I1(n26455), .I2(n54940), 
            .I3(\data_in_frame[15] [1]), .O(n14_adj_5488));
    defparam i6_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1162 (.I0(\data_in_frame[17] [2]), .I1(n14_adj_5488), 
            .I2(n10_adj_5487), .I3(\data_in_frame[12] [6]), .O(n54732));
    defparam i7_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1163 (.I0(n59563), .I1(\data_in_frame[19] [2]), 
            .I2(n59110), .I3(GND_net), .O(n59482));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1164 (.I0(n25605), .I1(n59482), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5489));
    defparam i2_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1165 (.I0(n7_adj_5489), .I1(\data_in_frame[17] [1]), 
            .I2(\data_in_frame[21] [3]), .I3(n61489), .O(n59553));
    defparam i4_4_lut_adj_1165.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_in_frame[19] [3]), .I1(n59482), 
            .I2(n54732), .I3(GND_net), .O(n54971));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_in_frame[14] [6]), .I1(n26447), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5490));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1168 (.I0(\data_in_frame[16] [7]), .I1(n59377), 
            .I2(\data_in_frame[17]_c [0]), .I3(n4_adj_5490), .O(n59563));   // verilog/coms.v(81[16:27])
    defparam i2_4_lut_adj_1168.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n30199), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n30198), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1169 (.I0(n59443), .I1(n61411), .I2(\data_in_frame[19] [1]), 
            .I3(n59563), .O(n10_adj_5491));
    defparam i4_4_lut_adj_1169.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n30197), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1170 (.I0(\data_in_frame[12] [2]), .I1(n59557), 
            .I2(n59097), .I3(n54016), .O(n55033));
    defparam i3_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n30196), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut_adj_1171 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[9] [4]), .I3(n59590), .O(n28_adj_5492));
    defparam i10_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(n26809), .I1(n28_adj_5492), .I2(\data_in_frame[12] [0]), 
            .I3(GND_net), .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n30195), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut_adj_1172 (.I0(Kp_23__N_1004), .I1(n59773), .I2(n54434), 
            .I3(n59294), .O(n30));
    defparam i12_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n30194), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_4_lut (.I0(n59174), .I1(\data_in_frame[6] [0]), .I2(\data_in_frame[9] [6]), 
            .I3(n53899), .O(n31_adj_5493));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[6]_c [5]), .I1(n59281), .I2(n59830), 
            .I3(n26231), .O(n29_adj_5494));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n29_adj_5494), .I1(n31_adj_5493), .I2(n30), 
            .I3(n32), .O(n54954));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n30193), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n30192), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51133_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66899));   // verilog/coms.v(158[12:15])
    defparam i51133_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n30191), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51367_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66900));   // verilog/coms.v(158[12:15])
    defparam i51367_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(n61489), .I1(n59110), .I2(GND_net), 
            .I3(GND_net), .O(n59758));
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h9999;
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n30190), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_211_i3_4_lut (.I0(n24160), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59413), .I3(n55047), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n30189), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n30188), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n30187), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i28328_3_lut (.I0(encoder0_position_scaled[13]), .I1(\motor_state_23__N_115[13] ), 
            .I2(n15), .I3(GND_net), .O(n10));
    defparam i28328_3_lut.LUT_INIT = 16'h3535;
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n30186), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1174 (.I0(n61411), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59566));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h9999;
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n30185), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50997_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66901));   // verilog/coms.v(158[12:15])
    defparam i50997_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5498), .S(n58934));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n30184), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n30183), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n30182), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n30181), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i50998_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66902));   // verilog/coms.v(158[12:15])
    defparam i50998_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50999_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66903));   // verilog/coms.v(158[12:15])
    defparam i50999_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51000_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66904));   // verilog/coms.v(158[12:15])
    defparam i51000_2_lut.LUT_INIT = 16'h2222;
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n30180), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n30179), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n30178), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n30177), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n30176), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n30175), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n30174), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n30173), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n30172), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n30171), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n30170), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n30169), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51001_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66905));   // verilog/coms.v(158[12:15])
    defparam i51001_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5499), .S(n58933));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51002_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66906));   // verilog/coms.v(158[12:15])
    defparam i51002_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5500), .S(n58932));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n30168), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n30167), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1175 (.I0(\data_in_frame[21] [2]), .I1(n59566), 
            .I2(\data_in_frame[18] [7]), .I3(n59758), .O(n10_adj_5501));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n30166), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n30165), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n30164), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5502), .S(n58931));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1176 (.I0(n61452), .I1(n10_adj_5501), .I2(\data_in_frame[18] [6]), 
            .I3(GND_net), .O(n59423));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_adj_1176.LUT_INIT = 16'h6969;
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n30163), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1177 (.I0(n54971), .I1(n59553), .I2(\data_in_frame[21] [4]), 
            .I3(GND_net), .O(n59755));
    defparam i2_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5503), .S(n58930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5504), .S(n58929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5505), .S(n58928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5506), .S(n58927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n30162), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5507), .S(n58926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n30161), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1178 (.I0(n26598), .I1(\data_in_frame[18] [7]), 
            .I2(n59514), .I3(n6_adj_5508), .O(n60966));
    defparam i4_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1179 (.I0(n60966), .I1(n59755), .I2(n59423), 
            .I3(\data_in_frame[21] [1]), .O(n10_adj_5509));
    defparam i4_4_lut_adj_1179.LUT_INIT = 16'h9669;
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n30160), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1180 (.I0(n59476), .I1(n10_adj_5509), .I2(\data_in_frame[21] [7]), 
            .I3(GND_net), .O(n59821));
    defparam i5_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n30159), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n30158), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[18] [6]), .I1(n59729), .I2(GND_net), 
            .I3(GND_net), .O(n42));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5510), .S(n58925));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1117_9_lut (.I0(n58814), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n51498), .O(n58816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1117_8_lut (.I0(n58814), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n51497), .O(n58817)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_8_lut.LUT_INIT = 16'h8228;
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n30157), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5511), .S(n58924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5512), .S(n58826));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n30156), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n30155), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n30154), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5513), .S(n58923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5514), .S(n58922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5515), .S(n58921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n30153), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5516), .S(n58920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n30152), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51366_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66907));   // verilog/coms.v(158[12:15])
    defparam i51366_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n30151), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n30150), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n30149), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5517), .S(n58919));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1117_8 (.CI(n51497), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n51498));
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5518), .S(n58918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5519), .S(n58917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n30148), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51124_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66908));   // verilog/coms.v(158[12:15])
    defparam i51124_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n30147), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n30146), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5520), .S(n58916));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1181 (.I0(n59827), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5521));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i51115_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66909));   // verilog/coms.v(158[12:15])
    defparam i51115_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5522), .S(n58915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n30145), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5523), .S(n58914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5524), .S(n58913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5525), .S(n58912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n30144), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51241_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66912));   // verilog/coms.v(158[12:15])
    defparam i51241_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_4_lut_adj_1182 (.I0(n59746), .I1(n59749), .I2(\data_out_frame[24] [0]), 
            .I3(n54411), .O(n12_adj_5526));
    defparam i5_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i51043_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66913));   // verilog/coms.v(158[12:15])
    defparam i51043_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n30143), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n30142), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n30141), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n30140), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n30139), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n30138), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n30137), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51114_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66917));   // verilog/coms.v(158[12:15])
    defparam i51114_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51053_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66918));   // verilog/coms.v(158[12:15])
    defparam i51053_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i20_4_lut (.I0(n59514), .I1(n59758), .I2(\data_in_frame[19] [6]), 
            .I3(n59461), .O(n57_adj_5527));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i51112_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66919));   // verilog/coms.v(158[12:15])
    defparam i51112_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n30136), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n30135), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n30134), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n30133), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i29_4_lut (.I0(n57_adj_5527), .I1(n55066), .I2(n42), .I3(\data_in_frame[20] [6]), 
            .O(n66));
    defparam i29_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut (.I0(n26376), .I1(n61411), .I2(n26902), .I3(\data_in_frame[15] [4]), 
            .O(n64));
    defparam i27_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5528), .S(n58911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5529), .S(n58910));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n30132), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n30131), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n30130));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n30129));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n30128));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n30127));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5530), .S(n58909));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i28_4_lut (.I0(\data_in_frame[15] [2]), .I1(Kp_23__N_1518), 
            .I2(\data_in_frame[16]_c [1]), .I3(n38), .O(n65));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5531), .S(n58908));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1117_7_lut (.I0(n58814), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n51496), .O(n58818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_7_lut.LUT_INIT = 16'h8228;
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5532), .S(n58907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5533), .S(n58906));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n30126));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51120_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66921));   // verilog/coms.v(158[12:15])
    defparam i51120_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1183 (.I0(\FRAME_MATCHER.state[3] ), .I1(\data_out_frame[24] [1]), 
            .I2(n12_adj_5526), .I3(n8_adj_5521), .O(n3_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'h2882;
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n30125));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n30124));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n30123));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n30122));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n30121));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n30120), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51055_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66922));   // verilog/coms.v(158[12:15])
    defparam i51055_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i26_4_lut (.I0(n26197), .I1(n59720), .I2(n59732), .I3(n59653), 
            .O(n63));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30119), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30115), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5535), .S(n58905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5536), .S(n58904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30112), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5538), .S(n58903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30108), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1117_7 (.CI(n51496), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n51497));
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30107), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30106), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30105), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5540), .S(n58902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5541), .S(n58901));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[20][0] ), .I3(GND_net), .O(n44));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_1117_6_lut (.I0(n58814), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n51495), .O(n58819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1184 (.I0(n54900), .I1(n59824), .I2(n59746), 
            .I3(n59493), .O(n24160));
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n59678), .I1(n27228), .I2(n59138), .I3(\data_in_frame[15] [6]), 
            .O(n62));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n54959), .I1(\data_in_frame[15] [3]), .I2(n59517), 
            .I3(n59818), .O(n61));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n63), .I1(n65), .I2(n64), .I3(n66), .O(n72));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n59488), .I1(n60_adj_5542), .I2(n44), .I3(n59338), 
            .O(n67));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i36_4_lut (.I0(n67), .I1(n72), .I2(n61), .I3(n62), .O(n54957));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1117_6 (.CI(n51495), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n51496));
    SB_LUT4 i2_3_lut_adj_1185 (.I0(n61452), .I1(n59735), .I2(\data_in_frame[20] [6]), 
            .I3(GND_net), .O(n59464));
    defparam i2_3_lut_adj_1185.LUT_INIT = 16'h6969;
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30101), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1186 (.I0(n59309), .I1(n24160), .I2(n54397), 
            .I3(n59507), .O(n10_adj_5543));
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1187 (.I0(n26395), .I1(n26376), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n33));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1188 (.I0(n54952), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n59147));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1188.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1189 (.I0(\data_in_frame[11] [6]), .I1(n24389), 
            .I2(n26134), .I3(n26878), .O(n59331));
    defparam i3_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1190 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[15] [6]), 
            .I2(n26189), .I3(n6_adj_5544), .O(n59242));
    defparam i4_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_in_frame[10] [2]), .I1(n59545), 
            .I2(n24393), .I3(n59762), .O(n54440));
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_209_i3_4_lut (.I0(n54943), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5543), .I3(n61148), .O(n3_adj_5545));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(n26902), .I1(n54440), .I2(GND_net), 
            .I3(GND_net), .O(n54940));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1193 (.I0(\data_in_frame[10] [0]), .I1(n24389), 
            .I2(Kp_23__N_1214), .I3(n24393), .O(n54434));
    defparam i2_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1194 (.I0(\data_in_frame[12] [2]), .I1(n54434), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n59504));
    defparam i2_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n30090));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30089), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30088), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30087), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30086), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30085), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_12__7__I_0_4035_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_798));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_12__7__I_0_4035_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30084), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30083), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30082), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30081), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30080), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30079), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1195 (.I0(\data_in_frame[10] [1]), .I1(n27255), 
            .I2(n26316), .I3(GND_net), .O(n59699));
    defparam i2_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1196 (.I0(\data_in_frame[11] [7]), .I1(n59699), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n59557));
    defparam i2_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30078), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30077), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30076), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i53726_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[8]_c [2]), 
            .I2(n59971), .I3(GND_net), .O(n58444));   // verilog/coms.v(94[13:20])
    defparam i53726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1197 (.I0(\data_in_frame[10] [3]), .I1(n26809), 
            .I2(n59578), .I3(n6_adj_5546), .O(n26902));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i15986_3_lut (.I0(\data_in_frame[8]_c [1]), .I1(rx_data[1]), 
            .I2(n59971), .I3(GND_net), .O(n30393));   // verilog/coms.v(130[12] 305[6])
    defparam i15986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(n26455), .I1(n26902), .I2(\data_in_frame[12] [5]), 
            .I3(GND_net), .O(n26447));
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 select_1727_Select_0_i1_2_lut (.I0(tx_transmit_N_3545), .I1(\FRAME_MATCHER.i_31__N_2640 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5547));   // verilog/coms.v(148[4] 304[11])
    defparam select_1727_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n30075));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i53725_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[8]_c [0]), 
            .I2(n59971), .I3(GND_net), .O(n58438));   // verilog/coms.v(94[13:20])
    defparam i53725_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n30074));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23770_3_lut (.I0(n59994), .I1(rx_data[6]), .I2(\data_in_frame[7] [6]), 
            .I3(GND_net), .O(n30646));   // verilog/coms.v(94[13:20])
    defparam i23770_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 select_810_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1199 (.I0(\data_in_frame[9] [0]), .I1(n54659), 
            .I2(n26687), .I3(n6_adj_5548), .O(n59773));
    defparam i4_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n64526), .I2(n64527), .I3(\byte_transmit_counter[2] ), 
            .O(n70909));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_3_lut (.I0(n59557), .I1(\data_in_frame[8][7] ), .I2(\data_in_frame[8] [6]), 
            .I3(GND_net), .O(n25));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 n70909_bdd_4_lut (.I0(n70909), .I1(n64503), .I2(n64502), .I3(\byte_transmit_counter[2] ), 
            .O(n70912));
    defparam n70909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut_adj_1200 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[11] [3]), 
            .I2(n59377), .I3(n59773), .O(n33_adj_5549));
    defparam i12_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5550), .S(n58900));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17_4_lut_adj_1201 (.I0(n33_adj_5549), .I1(n25), .I2(\data_in_frame[9] [5]), 
            .I3(\data_in_frame[11] [2]), .O(n38_adj_5551));
    defparam i17_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n59107), .I1(n59762), .I2(n27142), .I3(n24393), 
            .O(n36));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i53724_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[6]_c [6]), 
            .I2(n28801), .I3(GND_net), .O(n58434));   // verilog/coms.v(94[13:20])
    defparam i53724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53723_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[6]_c [5]), 
            .I2(n28801), .I3(GND_net), .O(n58428));   // verilog/coms.v(94[13:20])
    defparam i53723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_3_lut_adj_1202 (.I0(rx_data[2]), .I1(\data_in_frame[6][2] ), 
            .I2(n28801), .I3(GND_net), .O(n58446));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1202.LUT_INIT = 16'hcaca;
    SB_LUT4 select_810_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i53729_4_lut (.I0(n59522), .I1(n55073), .I2(n4_adj_5552), 
            .I3(n54896), .O(n69904));
    defparam i53729_4_lut.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n30073));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n30072));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54864 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n71077));
    defparam byte_transmit_counter_0__bdd_4_lut_54864.LUT_INIT = 16'he4aa;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n30071));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n30070));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n30069));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n30068));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n30067));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n30066));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_208_i3_4_lut (.I0(n69904), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[25] [6]), .I3(n54694), .O(n3_adj_5553));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n30062));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n30061));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n30059));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n30057));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n30027));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n30011), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n30010));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n30009));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n30008));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1203 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5554));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1203.LUT_INIT = 16'ha088;
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n30007), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n30006), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n30002), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29998), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5555), .S(n58899));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5556));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1204 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[25] [5]), 
            .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5557));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1204.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5558), .S(n58829));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5559), .S(n58832));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5560), .S(n58833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5561), .S(n58834));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5562), .S(n58835));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5563), .S(n58836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5564), .S(n58841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5565), .S(n58843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5566), .S(n58847));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5567), .S(n58848));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5568), .S(n58849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5569), .S(n58850));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5570), .S(n58844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5571), .S(n58851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5572), .S(n58852));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5573), .S(n58846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5574), .S(n58853));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5575), .S(n58854));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5576), .S(n58855));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5577), .S(n58856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5578), .S(n58857));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1205 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[25] [4]), 
            .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5579));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1205.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5580), .S(n58858));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5581), .S(n58859));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5582), .S(n58827));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54694 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64493), .I2(n64494), .I3(\byte_transmit_counter[2] ), 
            .O(n70903));
    defparam byte_transmit_counter_1__bdd_4_lut_54694.LUT_INIT = 16'he4aa;
    SB_LUT4 i16_4_lut_adj_1206 (.I0(\data_in_frame[11] [4]), .I1(Kp_23__N_798), 
            .I2(n54030), .I3(n22_adj_5583), .O(n37));
    defparam i16_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 add_1117_5_lut (.I0(n58814), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n51494), .O(n58820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14_4_lut_adj_1207 (.I0(\data_in_frame[12] [5]), .I1(n59638), 
            .I2(n59657), .I3(n59504), .O(n35));
    defparam i14_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1208 (.I0(n35), .I1(n37), .I2(n36), .I3(n38_adj_5551), 
            .O(n54952));
    defparam i20_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5584));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1209 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n59485));
    defparam i2_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_CARRY add_1117_5 (.CI(n51494), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n51495));
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_in_frame[11] [2]), .I1(n26719), 
            .I2(GND_net), .I3(GND_net), .O(n59714));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1211 (.I0(\data_in_frame[13] [3]), .I1(n59714), 
            .I2(\data_in_frame[11] [0]), .I3(n59446), .O(n12_adj_5585));
    defparam i5_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1212 (.I0(\data_in_frame[9] [1]), .I1(n12_adj_5585), 
            .I2(\data_in_frame[15] [4]), .I3(n59485), .O(n61866));
    defparam i6_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17][7] ), 
            .I1(\data_in_frame[17][6] ), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1518));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[13] [1]), .I1(n54952), .I2(n59741), 
            .I3(GND_net), .O(n8_adj_5586));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_in_frame[14] [0]), .I1(n59331), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5587));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1214 (.I0(n26376), .I1(n59524), .I2(n8_adj_5586), 
            .I3(n59726), .O(n12_adj_5588));
    defparam i3_4_lut_adj_1214.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5589));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1117_4_lut (.I0(n58814), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n51493), .O(n58821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1117_4 (.CI(n51493), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n51494));
    SB_LUT4 select_810_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5590));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1215 (.I0(n59242), .I1(\data_in_frame[16]_c [0]), 
            .I2(\data_in_frame[13] [3]), .I3(n10_adj_5587), .O(n16_adj_5591));
    defparam i7_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1216 (.I0(n59741), .I1(n16_adj_5591), .I2(n12_adj_5588), 
            .I3(n59147), .O(n60999));
    defparam i8_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1217 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[13] [4]), 
            .I2(n59242), .I3(n6_adj_5592), .O(n59341));
    defparam i4_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2052__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n28405), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i4_4_lut_adj_1218 (.I0(n59171), .I1(Kp_23__N_1007), .I2(n26687), 
            .I3(n59276), .O(n10_adj_5593));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1219 (.I0(\data_in_frame[11] [3]), .I1(n26357), 
            .I2(n10_adj_5593), .I3(\data_in_frame[8][7] ), .O(n26376));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n59650));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1221 (.I0(n26296), .I1(\data_in_frame[8]_c [0]), 
            .I2(n26809), .I3(n6_adj_5594), .O(n26316));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_in_frame[8]_c [1]), .I1(\data_in_frame[8]_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59764));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(n26719), .I1(n26878), .I2(GND_net), 
            .I3(GND_net), .O(n27142));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5595));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5596));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26134));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1214));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5597), .S(n58860));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5598), .S(n58861));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_2052__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n28407), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n28409), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i2_3_lut_adj_1225 (.I0(Kp_23__N_1214), .I1(n26134), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n59097));
    defparam i2_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1226 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26687));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_DFFR \FRAME_MATCHER.i_2052__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n28411), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n28413), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n28415), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n28417), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n28419), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n28421), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n28423), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n28425), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28427), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28429), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28431), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28433), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28435), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28437), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28439), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28441), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28443), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28445), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28447), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28449), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28451), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28453), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28455), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28457), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n28459), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n28461), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n28463), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28465), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2052__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28467), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5599), .S(n58862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5600), .S(n58863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5601), .S(n58864));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1227 (.I0(\data_in_frame[9] [1]), .I1(n59300), 
            .I2(GND_net), .I3(GND_net), .O(n26189));
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1228 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(n6_adj_5602), .I3(n59060), .O(n27340));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1228.LUT_INIT = 16'haaa8;
    SB_LUT4 i53806_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3674[0]), 
            .I2(n44648), .I3(GND_net), .O(tx_transmit_N_3545));
    defparam i53806_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 select_810_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5603));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1229 (.I0(Kp_23__N_1209), .I1(n27142), .I2(n8_adj_5604), 
            .I3(n59762), .O(n12_adj_5605));
    defparam i3_4_lut_adj_1229.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1230 (.I0(n59395), .I1(n59191), .I2(n59300), 
            .I3(n10_adj_5606), .O(n16_adj_5607));
    defparam i7_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1231 (.I0(n59764), .I1(n16_adj_5607), .I2(n12_adj_5605), 
            .I3(n59312), .O(n53899));
    defparam i8_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3674[0]), 
            .I2(n44648), .I3(\FRAME_MATCHER.i_31__N_2640 ), .O(n25927));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i29593_2_lut (.I0(LED_c), .I1(LED_N_3537), .I2(GND_net), .I3(GND_net), 
            .O(LED_N_3536));   // verilog/coms.v(253[15] 255[9])
    defparam i29593_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1232 (.I0(\data_in_frame[16]_c [1]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n59524));
    defparam i2_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i14856_4_lut (.I0(n3358), .I1(LED_N_3536), .I2(n27759), .I3(\FRAME_MATCHER.i_31__N_2642 ), 
            .O(n29263));   // verilog/coms.v(130[12] 305[6])
    defparam i14856_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i6_4_lut_adj_1233 (.I0(n59799), .I1(\data_in_frame[14] [1]), 
            .I2(n54912), .I3(n59650), .O(n15_adj_5608));
    defparam i6_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1234 (.I0(n15_adj_5608), .I1(\data_in_frame[11] [7]), 
            .I2(n14_adj_5609), .I3(\data_in_frame[13] [7]), .O(n26598));
    defparam i8_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1235 (.I0(n26598), .I1(\data_in_frame[16]_c [2]), 
            .I2(n59524), .I3(n6_adj_5610), .O(n60988));
    defparam i4_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1236 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n53918), .I3(GND_net), .O(n54016));
    defparam i2_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 select_1725_Select_0_i3_3_lut (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n3_adj_5611));   // verilog/coms.v(148[4] 304[11])
    defparam select_1725_Select_0_i3_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_1117_3_lut (.I0(n58814), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n51492), .O(n58822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26389));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(n26281), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5481));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(\data_in_frame[9] [0]), .I1(n26365), 
            .I2(GND_net), .I3(GND_net), .O(n59446));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_in_frame[18] [3]), .I1(n60988), 
            .I2(GND_net), .I3(GND_net), .O(n55118));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5612), .S(n58845));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1241 (.I0(\data_in_frame[17][7] ), .I1(n59729), 
            .I2(n59510), .I3(\data_in_frame[15] [5]), .O(n25579));
    defparam i3_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1242 (.I0(\data_in_frame[1] [7]), .I1(n59533), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[4] [3]), .O(Kp_23__N_1007));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1243 (.I0(LED_c), .I1(n3_adj_5611), .I2(Kp_23__N_1877), 
            .I3(Kp_23__N_741), .O(n5_adj_5613));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1243.LUT_INIT = 16'hfcec;
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5614), .S(n59003));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5615), .S(n58865));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1244 (.I0(\data_in_frame[7][7] ), .I1(\data_in_frame[5] [5]), 
            .I2(n24221), .I3(GND_net), .O(n26809));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1245 (.I0(tx_active), .I1(r_SM_Main_2__N_3674[0]), 
            .I2(\FRAME_MATCHER.i_31__N_2640 ), .I3(n44648), .O(n61010));
    defparam i2_3_lut_4_lut_adj_1245.LUT_INIT = 16'h1000;
    SB_LUT4 i2_2_lut_adj_1246 (.I0(n59569), .I1(n26809), .I2(GND_net), 
            .I3(GND_net), .O(n59799));   // verilog/coms.v(81[16:27])
    defparam i2_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1247 (.I0(n53905), .I1(n59632), .I2(\data_out_frame[17] [2]), 
            .I3(n59212), .O(n12_adj_5616));
    defparam i5_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5617), .S(n59002));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1248 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[15] [2]), 
            .I2(n12_adj_5616), .I3(n8_adj_5618), .O(n55073));
    defparam i1_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1249 (.I0(\data_in_frame[5] [0]), .I1(n59644), 
            .I2(\data_in_frame[7][2] ), .I3(GND_net), .O(n26878));
    defparam i2_3_lut_adj_1249.LUT_INIT = 16'h9696;
    SB_LUT4 n70903_bdd_4_lut (.I0(n70903), .I1(n64509), .I2(n64508), .I3(\byte_transmit_counter[2] ), 
            .O(n70906));
    defparam n70903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1250 (.I0(\data_in_frame[6][7] ), .I1(n59276), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n26707));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5619), .S(n58866));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5620), .S(n59001));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_4_lut_adj_1251 (.I0(\data_in_frame[17]_c [0]), .I1(rx_data[0]), 
            .I2(n28780), .I3(n3942), .O(n58184));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1251.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[6]_c [6]), .I1(\data_in_frame[7][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n59590));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i20_2_lut (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26844));   // verilog/coms.v(99[12:25])
    defparam i20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1253 (.I0(n26844), .I1(n59573), .I2(n59130), 
            .I3(\data_in_frame[1] [4]), .O(n27255));
    defparam i3_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1254 (.I0(\data_out_frame[22] [1]), .I1(n55014), 
            .I2(n59141), .I3(n54996), .O(n18_adj_5621));
    defparam i7_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5622), .S(n59000));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5623), .S(n58999));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_in_frame[6][7] ), .I1(n26753), 
            .I2(GND_net), .I3(GND_net), .O(n59171));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n31074), .D(n2_adj_5624), .S(n29319));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1256 (.I0(n54889), .I1(n18_adj_5621), .I2(n61790), 
            .I3(n59723), .O(n20_adj_5625));
    defparam i9_4_lut_adj_1256.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1257 (.I0(n27255), .I1(n28_adj_5626), .I2(\data_in_frame[8]_c [2]), 
            .I3(GND_net), .O(n4_adj_5627));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1258 (.I0(n15_adj_5628), .I1(n20_adj_5625), .I2(\data_out_frame[21] [6]), 
            .I3(n61719), .O(n55047));
    defparam i10_4_lut_adj_1258.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n26231));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(n26756), .I1(\data_in_frame[4] [6]), 
            .I2(n59171), .I3(n6_adj_5629), .O(n26719));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n31075), .D(n2_adj_5630), .S(n29318));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5631), .S(n58998));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1260 (.I0(n26330), .I1(Kp_23__N_1001), .I2(Kp_23__N_998), 
            .I3(\data_in_frame[8][4] ), .O(n26365));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1261 (.I0(n26173), .I1(\data_in_frame[7] [6]), 
            .I2(n26333), .I3(GND_net), .O(n24393));
    defparam i2_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1262 (.I0(\data_in_frame[5] [3]), .I1(n59420), 
            .I2(n59365), .I3(\data_in_frame[7][4] ), .O(n59294));
    defparam i3_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(n55047), .I1(n2329), .I2(GND_net), 
            .I3(GND_net), .O(n59507));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_212_i3_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n59507), .I3(\data_out_frame[24] [3]), 
            .O(n3_adj_5632));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_212_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1264 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26756));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1264.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1265 (.I0(Kp_23__N_901), .I1(n26339), .I2(\data_in_frame[0] [0]), 
            .I3(n6_adj_5633), .O(Kp_23__N_1001));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[17] [3]), .I1(n61557), 
            .I2(GND_net), .I3(GND_net), .O(n59796));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[4] [7]), .I1(n59174), 
            .I2(GND_net), .I3(GND_net), .O(n27074));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(n26760), .I1(n59294), .I2(n5), .I3(GND_net), 
            .O(n24389));
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n29785));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1269 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2637 ), 
            .I2(n2436), .I3(n2439), .O(n25935));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1269.LUT_INIT = 16'h4000;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(\data_in_frame[8][5] ), .I1(n59264), 
            .I2(\data_in_frame[6][3] ), .I3(Kp_23__N_1001), .O(n26281));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30858));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1271 (.I0(n2436), .I1(n4452), .I2(n2439), 
            .I3(n2442), .O(n61096));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1271.LUT_INIT = 16'h2000;
    SB_LUT4 i4_4_lut_adj_1272 (.I0(n59796), .I1(n59479), .I2(\data_out_frame[15] [1]), 
            .I3(n59839), .O(n10_adj_5634));
    defparam i4_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n29788));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1273 (.I0(\data_in_frame[7][3] ), .I1(n27074), 
            .I2(n59365), .I3(n6_adj_5635), .O(n53918));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1274 (.I0(n59681), .I1(\data_out_frame[19] [5]), 
            .I2(n10_adj_5634), .I3(\data_out_frame[15] [3]), .O(n54900));
    defparam i1_4_lut_adj_1274.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1275 (.I0(\data_in_frame[3] [1]), .I1(n26617), 
            .I2(\data_in_frame[7][5] ), .I3(\data_in_frame[3] [3]), .O(n12_adj_5636));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n29792));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n29795));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n29798));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16]_c [0]), .C(clk16MHz), 
           .D(n29801));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16]_c [1]), .C(clk16MHz), 
           .D(n29804));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16]_c [2]), .C(clk16MHz), 
           .D(n29807));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16]_c [3]), .C(clk16MHz), 
           .D(n29810));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n30828));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\data_out_frame[20] [5]), .I1(n59407), 
            .I2(n53959), .I3(n61790), .O(n2329));
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1277 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_5636), 
            .I2(n59602), .I3(\data_in_frame[5] [3]), .O(n54659));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(reset), .I3(GND_net), .O(n23230));
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[5] [6]), .I1(n26333), 
            .I2(GND_net), .I3(GND_net), .O(n59573));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_213_i3_4_lut (.I0(n54397), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59315), .I3(n2329), .O(n3_adj_5637));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_213_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n30773));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16]_c [4]), .C(clk16MHz), 
           .D(n29815));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n30763));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16]_c [5]), .C(clk16MHz), 
           .D(n29818));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n30761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n30760));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n30313));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1279 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_928), 
            .I2(n26357), .I3(n6_adj_5638), .O(n59569));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n30744));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16]_c [6]), .C(clk16MHz), 
           .D(n29821));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n30742));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30741));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1280 (.I0(n53944), .I1(\data_in_frame[8]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59395));
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30739));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30737));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30736));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30735));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30733));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30732));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30731));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30730));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30729));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30728));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30727));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30726));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30725));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30724));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30723));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30722));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30721));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1281 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[6][1] ), 
            .I2(\data_in_frame[3] [7]), .I3(n6_adj_5639), .O(n59578));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30720));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30719));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30718));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30717));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30716));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30715));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30714));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30713));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30712));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30711));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n30710));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n29824));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n30316));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n30707));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n30706));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n30705));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17]_c [0]), .C(clk16MHz), 
           .D(n58184));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n30703));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26339));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n30702));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30699));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1283 (.I0(n54397), .I1(\data_out_frame[24] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5640));
    defparam i2_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n58296));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n30319));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n30322));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n29833));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n30326));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n30693));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30690));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n58294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n58290));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n58286));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1284 (.I0(\FRAME_MATCHER.state[3] ), .I1(\data_out_frame[24] [4]), 
            .I2(n6_adj_5640), .I3(n54943), .O(n3_adj_5641));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1284.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17][6] ), .C(clk16MHz), 
           .D(n58282));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17][7] ), .C(clk16MHz), 
           .D(n58278));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n58274));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n58272));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n58268));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29861));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n58264));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29867));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n58260));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n30677));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30674));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n58256));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1285 (.I0(\data_in_frame[1] [6]), .I1(n59251), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_998));   // verilog/coms.v(81[16:27])
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n30672));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30669));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29876));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29879));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29882));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n30664));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n30329));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n30332));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n30335));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n30338));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6][1] ), .C(clk16MHz), 
           .D(n30342));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6][2] ), .C(clk16MHz), 
           .D(n58446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6][3] ), .C(clk16MHz), 
           .D(n30348));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6][4] ), .C(clk16MHz), 
           .D(n30352));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6]_c [5]), .C(clk16MHz), 
           .D(n58428));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6]_c [6]), .C(clk16MHz), 
           .D(n58434));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6][7] ), .C(clk16MHz), 
           .D(n30361));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7][0] ), .C(clk16MHz), 
           .D(n30365));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7][1] ), .C(clk16MHz), 
           .D(n30368));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7][2] ), .C(clk16MHz), 
           .D(n30371));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7][3] ), .C(clk16MHz), 
           .D(n30375));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7][4] ), .C(clk16MHz), 
           .D(n30378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7][5] ), .C(clk16MHz), 
           .D(n30381));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n30646));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7][7] ), .C(clk16MHz), 
           .D(n30387));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8]_c [0]), .C(clk16MHz), 
           .D(n58438));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8]_c [1]), .C(clk16MHz), 
           .D(n30393));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8]_c [2]), .C(clk16MHz), 
           .D(n58444));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8][3] ), .C(clk16MHz), 
           .D(n30399));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8][4] ), .C(clk16MHz), 
           .D(n30403));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n30639));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n30638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8][5] ), .C(clk16MHz), 
           .D(n30406));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
           .D(n30409));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8][7] ), .C(clk16MHz), 
           .D(n30413));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n30416));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_in_frame[6][2] ), .I1(\data_in_frame[8][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n59312));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_4_lut (.I0(n2436), .I1(n4452), .I2(n4_adj_5418), 
            .I3(\FRAME_MATCHER.i_31__N_2643 ), .O(n61848));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i2_3_lut_adj_1287 (.I0(n28_adj_5626), .I1(n59312), .I2(Kp_23__N_998), 
            .I3(GND_net), .O(n26848));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1288 (.I0(n59527), .I1(n59705), .I2(\data_out_frame[25] [0]), 
            .I3(n54943), .O(n12_adj_5642));
    defparam i5_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1289 (.I0(\data_in_frame[0] [6]), .I1(n26302), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n26760));
    defparam i2_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n30419));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n30422));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n30425));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n30428));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n30431));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n30434));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_215_i3_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n12_adj_5642), .I3(n8_adj_5643), 
            .O(n3_adj_5644));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30437));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
           .D(n30440));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
           .D(n58460));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
           .D(n30446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n30449));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n30453));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n30456));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n30459));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n30462));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n30466));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n30469));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n30616));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n30475));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n30479));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n30482));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30485));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30489));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30492));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30495));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n30499));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n58384));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n58398));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n30509));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n30512));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30515));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30519));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30522));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30525));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30529));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n30532));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30536));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n30541));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n30545));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n30550));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n30554));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n30558));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
           .D(n30562));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n30566));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29888));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n29891));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n30587));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29894));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29897));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20][0] ), .C(clk16MHz), 
           .D(n58252));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20][1] ), .C(clk16MHz), 
           .D(n58248));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20][2] ), .C(clk16MHz), 
           .D(n58244));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20][3] ), .C(clk16MHz), 
           .D(n29909));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20][4] ), .C(clk16MHz), 
           .D(n29912));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20][5] ), .C(clk16MHz), 
           .D(n58238));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n58298));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(\FRAME_MATCHER.i [2]), .O(n60));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20][7] ), .C(clk16MHz), 
           .D(n58234));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n58230));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n58228));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n58226));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n58224));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n58220));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n58216));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n58212));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n58208));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29949));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1290 (.I0(n26786), .I1(\data_in_frame[4] [3]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n59357));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29952));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59805));
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(n59281), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[5] [1]), .I3(n59144), .O(n10_adj_5645));   // verilog/coms.v(169[9:87])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n58202));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13_2_lut (.I0(\data_in_frame[6]_c [5]), .I1(\data_in_frame[6]_c [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26357));   // verilog/coms.v(99[12:25])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29958));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_901));   // verilog/coms.v(81[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29961));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26296));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29964));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29968));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n58198));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n30539));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29977));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29980));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_216_i3_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5646), .I3(n59473), 
            .O(n3_adj_5647));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_216_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n29983));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n29986));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1294 (.I0(\data_out_frame[17] [2]), .I1(n59585), 
            .I2(n59165), .I3(n27181), .O(n54411));
    defparam i3_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1295 (.I0(n59602), .I1(\data_in_frame[3] [1]), 
            .I2(n59354), .I3(GND_net), .O(n59672));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n29992));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1296 (.I0(\data_in_frame[5] [4]), .I1(n59420), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n26173));
    defparam i2_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n29995));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_in_frame[5] [0]), .I1(Kp_23__N_928), 
            .I2(GND_net), .I3(GND_net), .O(n26750));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n30465));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1298 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n26333));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_out_frame[19] [3]), .I1(n54411), 
            .I2(GND_net), .I3(GND_net), .O(n54896));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n30003));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n30016));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1300 (.I0(\data_in_frame[3] [3]), .I1(n59354), 
            .I2(n26333), .I3(GND_net), .O(n24221));
    defparam i2_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59291));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1302 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [7]), 
            .I2(n26750), .I3(n18_adj_5648), .O(n30_adj_5649));
    defparam i13_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1303 (.I0(\data_out_frame[20] [0]), .I1(n54996), 
            .I2(\data_out_frame[22] [2]), .I3(n6_adj_5650), .O(n59560));
    defparam i4_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1304 (.I0(Kp_23__N_877), .I1(n26173), .I2(\data_in_frame[5] [3]), 
            .I3(n59672), .O(n28_adj_5651));
    defparam i11_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1305 (.I0(n59533), .I1(\data_in_frame[5] [6]), 
            .I2(n59291), .I3(\data_in_frame[5] [2]), .O(n29_adj_5652));
    defparam i12_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1306 (.I0(n59644), .I1(n59805), .I2(\data_in_frame[1] [3]), 
            .I3(n59357), .O(n27_adj_5653));
    defparam i10_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1307 (.I0(n27_adj_5653), .I1(n29_adj_5652), .I2(n28_adj_5651), 
            .I3(n30_adj_5649), .O(n53944));
    defparam i16_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59315));
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1309 (.I0(\data_out_frame[22] [1]), .I1(n59560), 
            .I2(n59273), .I3(n54966), .O(n61480));
    defparam i3_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1]_c [0]), .C(clk16MHz), 
           .D(n30019));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_in_frame[8]_c [1]), .I1(n53944), 
            .I2(GND_net), .I3(GND_net), .O(n59470));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1311 (.I0(n61480), .I1(n54889), .I2(\data_out_frame[21] [7]), 
            .I3(GND_net), .O(n59407));
    defparam i2_3_lut_adj_1311.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_in_frame[6][3] ), .I1(\data_in_frame[6][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n26330));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1313 (.I0(\data_out_frame[22] [3]), .I1(n59104), 
            .I2(\data_out_frame[22] [4]), .I3(GND_net), .O(n61255));
    defparam i2_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n30028));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1314 (.I0(\data_in_frame[6][4] ), .I1(n59830), 
            .I2(\data_in_frame[6][7] ), .I3(GND_net), .O(n59205));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59130));
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1316 (.I0(n53905), .I1(n26123), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n59681));
    defparam i2_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[22] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59141));
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n30031));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n30035));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n58340));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n59539));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1319 (.I0(n59539), .I1(n59130), .I2(n59205), 
            .I3(\data_in_frame[3] [6]), .O(n14_adj_5654));   // verilog/coms.v(81[16:27])
    defparam i6_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5459), .S(n58997));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59413));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1321 (.I0(n26231), .I1(n59470), .I2(n59168), 
            .I3(n26756), .O(n13));   // verilog/coms.v(81[16:27])
    defparam i5_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1322 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[15] [7]), 
            .I2(\data_in_frame[13] [3]), .I3(\data_in_frame[13] [4]), .O(n59726));
    defparam i1_2_lut_3_lut_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i48044_4_lut (.I0(n13), .I1(n7_adj_5655), .I2(n14_adj_5654), 
            .I3(n26848), .O(n64209));
    defparam i48044_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i6_4_lut_adj_1323 (.I0(n54694), .I1(\data_out_frame[20] [1]), 
            .I2(n27305), .I3(n59413), .O(n14_adj_5656));
    defparam i6_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i48077_4_lut (.I0(n53451), .I1(n64209), .I2(n59395), .I3(n59761), 
            .O(n64242));
    defparam i48077_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i11_4_lut_adj_1324 (.I0(n54659), .I1(n53918), .I2(n26281), 
            .I3(n24389), .O(n28_adj_5657));
    defparam i11_4_lut_adj_1324.LUT_INIT = 16'h0400;
    SB_LUT4 i12_4_lut_adj_1325 (.I0(n24393), .I1(n26365), .I2(n26719), 
            .I3(n4_adj_5627), .O(n29_adj_5658));
    defparam i12_4_lut_adj_1325.LUT_INIT = 16'h0002;
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5458), .S(n58996));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1326 (.I0(n61255), .I1(n59407), .I2(n59315), 
            .I3(n59363), .O(n13_adj_5659));
    defparam i5_4_lut_adj_1326.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1327 (.I0(n59545), .I1(n26707), .I2(n26878), 
            .I3(n7_adj_5660), .O(n27_adj_5661));
    defparam i10_4_lut_adj_1327.LUT_INIT = 16'h0002;
    SB_LUT4 i16_4_lut_adj_1328 (.I0(n27_adj_5661), .I1(n29_adj_5658), .I2(n28_adj_5657), 
            .I3(n64242), .O(LED_N_3537));
    defparam i16_4_lut_adj_1328.LUT_INIT = 16'h0080;
    SB_LUT4 i4_4_lut_adj_1329 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[22] [0]), .I3(\data_in_frame[21] [6]), .O(n10_adj_5662));
    defparam i4_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5457), .S(n58995));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5456), .S(n58994));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5455), .S(n58842));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1330 (.I0(\data_out_frame[24] [6]), .I1(n59749), 
            .I2(\data_out_frame[23] [5]), .I3(n55120), .O(n20_adj_5663));
    defparam i8_4_lut_adj_1330.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n31082), .D(n2_adj_5454), .S(n29317));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1331 (.I0(n13_adj_5659), .I1(n59440), .I2(n14_adj_5656), 
            .I3(GND_net), .O(n13_adj_5664));
    defparam i1_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5452), .S(n58993));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut_adj_1332 (.I0(n13_adj_5664), .I1(n20_adj_5663), .I2(n59845), 
            .I3(\data_out_frame[24] [7]), .O(n22_adj_5665));
    defparam i10_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1333 (.I0(\data_out_frame[24] [5]), .I1(n59824), 
            .I2(\data_out_frame[23] [2]), .I3(n59542), .O(n21));
    defparam i9_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1334 (.I0(\data_out_frame[25] [5]), .I1(n21), .I2(\data_out_frame[25] [6]), 
            .I3(n22_adj_5665), .O(n59842));   // verilog/coms.v(100[12:26])
    defparam i2_4_lut_adj_1334.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5437), .S(n58992));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5436), .S(n58991));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1335 (.I0(\data_in_frame[22] [5]), .I1(n59338), 
            .I2(n25579), .I3(\data_in_frame[18] [1]), .O(n61385));
    defparam i3_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59814));
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(n59814), .I1(n59583), .I2(n59363), 
            .I3(n59842), .O(n10_adj_5666));
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1338 (.I0(n59341), .I1(\data_in_frame[18] [2]), 
            .I2(n60999), .I3(n59647), .O(n10_adj_5667));
    defparam i4_4_lut_adj_1338.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_217_i3_4_lut (.I0(n59744), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5666), .I3(n55038), .O(n3_adj_5668));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_217_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_4_lut_adj_1339 (.I0(n59464), .I1(n54957), .I2(\data_in_frame[23] [0]), 
            .I3(n59821), .O(n61318));
    defparam i2_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1340 (.I0(\data_in_frame[22] [6]), .I1(n59461), 
            .I2(\data_in_frame[20][4] ), .I3(GND_net), .O(n61138));
    defparam i2_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n28140), 
            .D(n5169[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5435), .S(n58990));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1341 (.I0(n25579), .I1(n60988), .I2(\data_in_frame[20][1] ), 
            .I3(GND_net), .O(n14_adj_5669));
    defparam i5_3_lut_adj_1341.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1342 (.I0(n59437), .I1(\data_in_frame[19] [6]), 
            .I2(n55007), .I3(\data_in_frame[22] [2]), .O(n15_adj_5670));
    defparam i6_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1343 (.I0(n59285), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[22] [3]), .I3(n59647), .O(n10_adj_5671));
    defparam i4_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n28140), 
            .D(n5169[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1344 (.I0(n15_adj_5670), .I1(n54920), .I2(n14_adj_5669), 
            .I3(\data_in_frame[20][0] ), .O(n61218));
    defparam i8_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n28140), 
            .D(n5169[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n28140), 
            .D(n5169[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n28140), 
            .D(n5169[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n28140), 
            .D(n5169[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n28140), 
            .D(n5169[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1345 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(n59449), .I3(n54753), .O(n59383));
    defparam i1_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n28140), 
            .D(n5169[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n28140), 
            .D(n5169[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n28140), 
            .D(n5169[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n28140), 
            .D(n5169[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n28140), 
            .D(n5169[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2640 ), 
            .I2(GND_net), .I3(GND_net), .O(n58814));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n28140), 
            .D(n5169[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n28140), 
            .D(n5169[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n28140), 
            .D(n5169[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n28140), 
            .D(n5169[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n28140), 
            .D(n5169[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n28140), 
            .D(n5169[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n28140), 
            .D(n5169[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n28140), 
            .D(n5169[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n28140), 
            .D(n5169[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n28140), 
            .D(n5169[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n28140), 
            .D(n5169[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2636 ), 
            .C(clk16MHz), .D(n71150), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i3_4_lut_adj_1346 (.I0(\data_out_frame[17] [6]), .I1(n59660), 
            .I2(n59383), .I3(n26523), .O(n61719));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2637 ), 
            .C(clk16MHz), .D(n27436), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2638 ), 
            .C(clk16MHz), .D(n2533), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2534), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2640 ), 
            .C(clk16MHz), .D(n20798), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2641 ), 
            .C(clk16MHz), .D(n58084), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2642 ), 
            .C(clk16MHz), .D(n2545), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2643 ), 
            .C(clk16MHz), .D(n28024), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1][1] ), .C(clk16MHz), 
           .D(n30043));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5417), .S(n58989));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1347 (.I0(n61218), .I1(n54920), .I2(n10_adj_5671), 
            .I3(n60988), .O(n23_c));
    defparam i6_4_lut_adj_1347.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1348 (.I0(n59821), .I1(n54957), .I2(n59517), 
            .I3(\data_in_frame[18] [5]), .O(n14_adj_5672));
    defparam i6_4_lut_adj_1348.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1349 (.I0(\data_in_frame[22] [7]), .I1(n59735), 
            .I2(\data_in_frame[20][5] ), .I3(n55118), .O(n13_adj_5673));
    defparam i5_4_lut_adj_1349.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1350 (.I0(\data_in_frame[23] [6]), .I1(n59717), 
            .I2(n59488), .I3(\data_in_frame[21] [4]), .O(n60916));
    defparam i3_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1351 (.I0(n53451), .I1(Kp_23__N_1680), .I2(n10_adj_5662), 
            .I3(n61861), .O(n18_adj_5674));
    defparam i1_4_lut_adj_1351.LUT_INIT = 16'h1441;
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5416), .S(n58988));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i47881_3_lut (.I0(n60916), .I1(n13_adj_5673), .I2(n14_adj_5672), 
            .I3(GND_net), .O(n64044));
    defparam i47881_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i12_4_lut_adj_1352 (.I0(n23_c), .I1(n61145), .I2(\data_in_frame[23] [5]), 
            .I3(n59755), .O(n29_adj_5675));
    defparam i12_4_lut_adj_1352.LUT_INIT = 16'h0220;
    SB_LUT4 i2_2_lut_adj_1353 (.I0(\data_in_frame[22] [1]), .I1(n59437), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5676));
    defparam i2_2_lut_adj_1353.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1354 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[20][0] ), .I3(GND_net), .O(n7_adj_5677));
    defparam i1_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i47885_4_lut (.I0(n59423), .I1(n61385), .I2(n59553), .I3(\data_in_frame[23] [4]), 
            .O(n64048));
    defparam i47885_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i5_4_lut_adj_1355 (.I0(n27228), .I1(n7_adj_5677), .I2(\data_in_frame[19] [5]), 
            .I3(n8_adj_5676), .O(n61289));
    defparam i5_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1356 (.I0(\data_in_frame[22] [4]), .I1(n61318), 
            .I2(n10_adj_5667), .I3(\data_in_frame[20][3] ), .O(n22_adj_5678));
    defparam i5_4_lut_adj_1356.LUT_INIT = 16'h8448;
    SB_LUT4 i43841_2_lut_3_lut (.I0(n3942), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n59967));
    defparam i43841_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i47883_4_lut (.I0(\data_in_frame[23] [1]), .I1(n61138), .I2(n54957), 
            .I3(n59821), .O(n64046));
    defparam i47883_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 select_810_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15_4_lut_adj_1357 (.I0(n29_adj_5675), .I1(n64044), .I2(n61159), 
            .I3(n18_adj_5674), .O(n32_adj_5679));
    defparam i15_4_lut_adj_1357.LUT_INIT = 16'h0200;
    SB_LUT4 select_810_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i10_4_lut_adj_1358 (.I0(n61289), .I1(n64048), .I2(\data_in_frame[23] [7]), 
            .I3(n59476), .O(n27_adj_5680));
    defparam i10_4_lut_adj_1358.LUT_INIT = 16'h0110;
    SB_LUT4 i16_4_lut_adj_1359 (.I0(n27_adj_5680), .I1(n32_adj_5679), .I2(n64046), 
            .I3(n22_adj_5678), .O(Kp_23__N_741));
    defparam i16_4_lut_adj_1359.LUT_INIT = 16'h0800;
    SB_LUT4 i53761_4_lut (.I0(\FRAME_MATCHER.i_31__N_2642 ), .I1(Kp_23__N_741), 
            .I2(LED_N_3537), .I3(Kp_23__N_1877), .O(n28140));
    defparam i53761_4_lut.LUT_INIT = 16'hc4a0;
    SB_LUT4 i2_3_lut_adj_1360 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [6]), .I3(GND_net), .O(n59473));
    defparam i2_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(n53959), .I1(n55014), .I2(\data_out_frame[20] [3]), 
            .I3(\data_out_frame[22] [5]), .O(n55038));
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1362 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1362.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5415), .S(n58867));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5414), .S(n58868));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_5681));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1363 (.I0(n26113), .I1(n59404), .I2(n54669), 
            .I3(\data_out_frame[16] [3]), .O(n59416));
    defparam i2_3_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5413), .S(n58987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5412), .S(n58986));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5411), .S(n58985));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5410), .S(n58984));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5409), .S(n58869));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16_4_lut_adj_1364 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_5682));
    defparam i16_4_lut_adj_1364.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1365 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut_adj_1365.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1366 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_1366.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1367 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut_adj_1367.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut_adj_1368 (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut_adj_1368.LUT_INIT = 16'heeee;
    SB_LUT4 select_810_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5408), .S(n58840));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i24_4_lut_adj_1369 (.I0(n41), .I1(n43), .I2(n42_adj_5682), 
            .I3(n44_adj_5681), .O(n50));
    defparam i24_4_lut_adj_1369.LUT_INIT = 16'hfffe;
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5407), .S(n58839));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1370 (.I0(n45), .I1(n50), .I2(n39), .I3(n40), 
            .O(n25998));
    defparam i25_4_lut_adj_1370.LUT_INIT = 16'hfffe;
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5406), .S(n58983));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i29745_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25998), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i29745_4_lut.LUT_INIT = 16'h3230;
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5404), .S(n58982));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_218_i3_4_lut (.I0(n55038), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5683), .I3(n59547), .O(n3_adj_5684));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i503_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2643 ), .I2(GND_net), 
            .I3(GND_net), .O(n2553));   // verilog/coms.v(148[4] 304[11])
    defparam i503_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5402), .S(n58981));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5434));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\data_out_frame[23] [0]), .I1(n61040), 
            .I2(GND_net), .I3(GND_net), .O(n59547));
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1372 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[7] [5]), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1372.LUT_INIT = 16'ha088;
    SB_LUT4 select_810_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1373 (.I0(n26237), .I1(n59371), .I2(n59254), 
            .I3(\data_out_frame[16] [3]), .O(n54889));
    defparam i3_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1374 (.I0(\data_out_frame[13] [5]), .I1(n25546), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n59449));
    defparam i2_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54814 (.I0(byte_transmit_counter_c[3]), 
            .I1(n68989), .I2(n66942), .I3(byte_transmit_counter_c[4]), 
            .O(n70879));
    defparam byte_transmit_counter_3__bdd_4_lut_54814.LUT_INIT = 16'he4aa;
    SB_LUT4 n70879_bdd_4_lut (.I0(n70879), .I1(n70792), .I2(n7_adj_5685), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n70879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54689 (.I0(\byte_transmit_counter[1] ), 
            .I1(n4_adj_5686), .I2(n5_adj_5687), .I3(\byte_transmit_counter[2] ), 
            .O(n70873));
    defparam byte_transmit_counter_1__bdd_4_lut_54689.LUT_INIT = 16'he4aa;
    SB_LUT4 n70873_bdd_4_lut (.I0(n70873), .I1(n67007), .I2(n67006), .I3(\byte_transmit_counter[2] ), 
            .O(n70876));
    defparam n70873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54744 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n70867));
    defparam byte_transmit_counter_0__bdd_4_lut_54744.LUT_INIT = 16'he4aa;
    SB_LUT4 n70867_bdd_4_lut (.I0(n70867), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n64401));
    defparam n70867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5688), .S(n58870));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1375 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n42166), .O(n28770));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1375.LUT_INIT = 16'h4000;
    SB_LUT4 select_810_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5429));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1376 (.I0(\data_out_frame[18] [1]), .I1(n59693), 
            .I2(n59431), .I3(n54945), .O(n10_adj_5689));
    defparam i4_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5690), .S(n58871));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1377 (.I0(n59449), .I1(n10_adj_5689), .I2(\data_out_frame[15] [7]), 
            .I3(GND_net), .O(n59660));
    defparam i5_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1378 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n59083), .O(n59086));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1378.LUT_INIT = 16'hffbf;
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5691), .S(n29311));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5692), .S(n58872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5693), .S(n58873));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5694), .S(n58874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5695), .S(n58875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5696), .S(n58876));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_338_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5697));   // verilog/coms.v(157[7:23])
    defparam equal_338_i7_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1379 (.I0(n3942), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57), .I3(reset), .O(n42166));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1379.LUT_INIT = 16'h0020;
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5698), .S(n58877));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5699), .S(n58878));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1380 (.I0(n3942), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57), .I3(n8_adj_10), .O(n28725));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(n55014), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n55120));
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h6666;
    SB_LUT4 i14074_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28480));   // verilog/coms.v(109[34:55])
    defparam i14074_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5701), .S(n58879));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1382 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59527));
    defparam i1_2_lut_adj_1382.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5702), .S(n58838));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48275_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64449));
    defparam i48275_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5703), .S(n58880));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48276_4_lut (.I0(n64449), .I1(n28480), .I2(\byte_transmit_counter[2] ), 
            .I3(byte_transmit_counter[0]), .O(n64450));
    defparam i48276_4_lut.LUT_INIT = 16'haca0;
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5704), .S(n58837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5705), .S(n58881));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48274_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64448));
    defparam i48274_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5706), .S(n58882));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1117_3 (.CI(n51492), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n51493));
    SB_LUT4 add_1117_2_lut (.I0(n58814), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3545), .I3(GND_net), .O(n58815)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1117_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1383 (.I0(n3942), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57), .I3(n8_adj_11), .O(n28717));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1383.LUT_INIT = 16'hffdf;
    SB_CARRY add_1117_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3545), 
            .CO(n51492));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1384 (.I0(n3942), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57), .I3(n8_adj_12), .O(n28733));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1384.LUT_INIT = 16'hffdf;
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5709), .S(n58980));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5710), .S(n58979));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(n59578), .O(n28_adj_5626));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5711), .S(n58883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5712), .S(n58978));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5713), .S(n58977));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5714), .S(n58884));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5715), .S(n58885));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1386 (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5716));
    defparam i2_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i51031_2_lut (.I0(n70756), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n67088));
    defparam i51031_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1387 (.I0(n53903), .I1(n54889), .I2(n59547), 
            .I3(\data_out_frame[22] [6]), .O(n14_adj_5717));
    defparam i6_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5718), .S(n58831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5719), .S(n58830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5720), .S(n58886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5721), .S(n58887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5722), .S(n58888));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1388 (.I0(n59550), .I1(n14_adj_5717), .I2(n10_adj_5716), 
            .I3(n59527), .O(n59744));
    defparam i7_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5723), .S(n58889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5724), .S(n58890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5725), .S(n58891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5726), .S(n58892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5727), .S(n58893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5728), .S(n58894));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5729), .S(n29283));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5730), .S(n58816));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5731), .S(n58817));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5732), .S(n58818));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5733), .S(n58819));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5734), .S(n58820));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5735), .S(n58821));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), 
            .C(clk16MHz), .E(n3358), .D(n1_adj_5736), .S(n58822));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5737), .S(n58798));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27][6] ), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5738), .S(n58799));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5739), .S(n58800));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5740), .S(n58796));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5741), .S(n58801));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5684), .S(n58802));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5668), .S(n58803));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5647), .S(n58804));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5644), .S(n58805));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26][6] ), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5641), .S(n58806));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5637), .S(n58807));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5632), .S(n58797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n3358), .D(n5_adj_5613), 
            .S(n29263));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5603), .S(n58895));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n3358), .D(n27340), 
            .S(n29261));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5596), .S(n58824));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n31162), .D(n2_adj_5595), .S(n29256));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n31163), .D(n2_adj_5590), .S(n29255));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n31164), .D(n2_adj_5589), .S(n29254));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5584), .S(n58896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n31166), .D(n2_adj_5579), .S(n29251));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5557), .S(n58897));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5556), .S(n58898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5554), .S(n58828));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5553), .S(n58808));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3674[0]), .C(clk16MHz), 
            .E(n3358), .D(n1_adj_5547), .S(n29241));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52904_3_lut (.I0(n70732), .I1(n70984), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n69079));
    defparam i52904_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5545), .S(n58809));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5539), .S(n58976));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1389 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n59077), .O(n59079));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'hfffb;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5537), .S(n58975));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n3358), .D(n1_adj_5742), .S(n58815));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n3358), .D(n3_adj_5534), .S(n58810));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n3358), .D(n3), .S(n58795));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5495), .S(n58974));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_810_Select_219_i3_2_lut (.I0(n59744), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5741));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_219_i3_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n3358), .D(n2_adj_5477), .S(n58973));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1390 (.I0(n54669), .I1(n69908), .I2(GND_net), 
            .I3(GND_net), .O(n59371));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1391 (.I0(\data_out_frame[21] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(\data_out_frame[23] [1]), .I3(GND_net), .O(n59440));
    defparam i2_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1392 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59693));
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1393 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n42166), .O(n28778));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1393.LUT_INIT = 16'h0400;
    SB_LUT4 i4_4_lut_adj_1394 (.I0(n7_adj_5743), .I1(n26970), .I2(n69908), 
            .I3(n59693), .O(n59318));
    defparam i4_4_lut_adj_1394.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(n25517), .I1(\data_out_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5744));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_33_lut  (.I0(n67000), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n52702), .O(n28407)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_32_lut  (.I0(n66982), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n52701), .O(n28409)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_32  (.CI(n52701), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n52702));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_31_lut  (.I0(n66947), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n52700), .O(n28411)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_31  (.CI(n52700), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n52701));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_30_lut  (.I0(n66946), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n52699), .O(n28413)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut_adj_1396 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [5]), .I3(n6_adj_5744), .O(n59845));
    defparam i4_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_30  (.CI(n52699), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n52700));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_29_lut  (.I0(n66945), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n52698), .O(n28415)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_29  (.CI(n52698), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n52699));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_28_lut  (.I0(n66944), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n52697), .O(n28417)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_28  (.CI(n52697), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n52698));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_27_lut  (.I0(n66943), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n52696), .O(n28419)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_27  (.CI(n52696), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n52697));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_26_lut  (.I0(n66940), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n52695), .O(n28421)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_26  (.CI(n52695), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n52696));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_25_lut  (.I0(n66938), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n52694), .O(n28423)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_25  (.CI(n52694), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n52695));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_24_lut  (.I0(n66937), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n52693), .O(n28425)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_24  (.CI(n52693), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n52694));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_23_lut  (.I0(n66932), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n52692), .O(n28427)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_23  (.CI(n52692), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n52693));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_22_lut  (.I0(n66925), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n52691), .O(n28429)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_22  (.CI(n52691), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n52692));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_21_lut  (.I0(n66924), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n52690), .O(n28431)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_21  (.CI(n52690), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n52691));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_20_lut  (.I0(n66922), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n52689), .O(n28433)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_20  (.CI(n52689), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n52690));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_19_lut  (.I0(n66921), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n52688), .O(n28435)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut_adj_1397 (.I0(n59833), .I1(n59723), .I2(n59185), 
            .I3(n59845), .O(n10_adj_5745));
    defparam i4_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_19  (.CI(n52688), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n52689));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_18_lut  (.I0(n66919), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n52687), .O(n28437)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_18  (.CI(n52687), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n52688));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_17_lut  (.I0(n66918), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n52686), .O(n28439)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_17  (.CI(n52686), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n52687));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_16_lut  (.I0(n66917), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n52685), .O(n28441)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_16  (.CI(n52685), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n52686));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_15_lut  (.I0(n66913), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n52684), .O(n28443)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_15  (.CI(n52684), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n52685));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_14_lut  (.I0(n66912), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n52683), .O(n28445)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_14  (.CI(n52683), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n52684));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_13_lut  (.I0(n66909), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n52682), .O(n28447)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n26094));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1399 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(n59371), .I3(n6_adj_5746), .O(n61754));
    defparam i4_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_13  (.CI(n52682), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n52683));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_12_lut  (.I0(n66908), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n52681), .O(n28449)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i7_4_lut_adj_1400 (.I0(n59690), .I1(\data_out_frame[18] [5]), 
            .I2(n59440), .I3(\data_out_frame[16] [4]), .O(n18_adj_5747));
    defparam i7_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_12  (.CI(n52681), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n52682));
    SB_LUT4 i5_2_lut_adj_1401 (.I0(n54222), .I1(n61754), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_5748));
    defparam i5_2_lut_adj_1401.LUT_INIT = 16'h9999;
    SB_LUT4 i9_4_lut_adj_1402 (.I0(\data_out_frame[20] [7]), .I1(n18_adj_5747), 
            .I2(n25517), .I3(n59416), .O(n20_adj_5749));
    defparam i9_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_11_lut  (.I0(n66907), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n52680), .O(n28451)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_11  (.CI(n52680), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n52681));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54656 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n70855));
    defparam byte_transmit_counter_0__bdd_4_lut_54656.LUT_INIT = 16'he4aa;
    SB_LUT4 i10_4_lut_adj_1403 (.I0(n55026), .I1(n20_adj_5749), .I2(n16_adj_5748), 
            .I3(n61040), .O(n53903));
    defparam i10_4_lut_adj_1403.LUT_INIT = 16'h9669;
    SB_LUT4 n70855_bdd_4_lut (.I0(n70855), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n70858));
    defparam n70855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54651 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n70849));
    defparam byte_transmit_counter_0__bdd_4_lut_54651.LUT_INIT = 16'he4aa;
    SB_LUT4 n70849_bdd_4_lut (.I0(n70849), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n70852));
    defparam n70849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_10_lut  (.I0(n66906), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n52679), .O(n28453)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_10  (.CI(n52679), .I0(n28716), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n52680));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_9_lut  (.I0(n66905), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n52678), .O(n28455)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_9  (.CI(n52678), .I0(n28716), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n52679));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_8_lut  (.I0(n66904), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n52677), .O(n28457)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_8  (.CI(n52677), .I0(n28716), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n52678));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_7_lut  (.I0(n66903), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n52676), .O(n28459)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_7  (.CI(n52676), .I0(n28716), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n52677));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_6_lut  (.I0(n66902), .I1(n28716), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n52675), .O(n28461)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_6  (.CI(n52675), .I0(n28716), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n52676));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_5_lut  (.I0(n66901), .I1(n28716), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n52674), .O(n28463)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_5  (.CI(n52674), .I0(n28716), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n52675));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_4_lut  (.I0(n66900), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n52673), .O(n28465)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_4  (.CI(n52673), .I0(n28716), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n52674));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_3_lut  (.I0(n66899), .I1(n28716), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n52672), .O(n28467)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_3  (.CI(n52672), .I0(n28716), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n52673));
    SB_LUT4 \FRAME_MATCHER.i_2052_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2052_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2052_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n52672));
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n6_adj_5750));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1405 (.I0(n54991), .I1(n53903), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5751));
    defparam i2_2_lut_adj_1405.LUT_INIT = 16'h6666;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(n59121), .I2(n59245), 
            .I3(\data_in_frame[1] [7]), .O(n24));   // verilog/coms.v(169[9:87])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0990;
    SB_LUT4 select_810_Select_220_i3_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5751), .I3(\data_out_frame[25] [2]), 
            .O(n3_adj_5740));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_220_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i4_4_lut_adj_1406 (.I0(n59416), .I1(n59225), .I2(n54962), 
            .I3(n59663), .O(n10_adj_5752));
    defparam i4_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1407 (.I0(n59254), .I1(n10_adj_5752), .I2(n54916), 
            .I3(GND_net), .O(n55026));
    defparam i5_3_lut_adj_1407.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[20] [2]), .I1(n61719), 
            .I2(n55014), .I3(\data_out_frame[20] [3]), .O(n54966));
    defparam i1_2_lut_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26237));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h6666;
    SB_LUT4 select_812_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5742));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2640 ), 
            .I2(\FRAME_MATCHER.i_31__N_2643 ), .I3(GND_net), .O(n59060));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(n26523), .I1(n59360), .I2(GND_net), 
            .I3(GND_net), .O(n54161));
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1412 (.I0(\data_out_frame[22] [4]), .I1(n54966), 
            .I2(\data_out_frame[24] [0]), .I3(\data_out_frame[25] [7]), 
            .O(n59309));
    defparam i1_2_lut_3_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 select_812_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(\byte_transmit_counter[1] ), 
            .I3(GND_net), .O(n1_adj_5736));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1413 (.I0(\FRAME_MATCHER.i [5]), .I1(n57), .I2(GND_net), 
            .I3(GND_net), .O(n42164));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_adj_1413.LUT_INIT = 16'h4444;
    SB_LUT4 select_812_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n1_adj_5735));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_adj_1414 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n59100));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 select_812_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n1_adj_5734));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_812_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n1_adj_5733));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_812_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5732));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1415 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [0]), .O(n26509));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1416 (.I0(\data_out_frame[11] [1]), .I1(n59261), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n26123));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1416.LUT_INIT = 16'h9696;
    SB_LUT4 select_812_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5731));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_812_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2640 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5730));   // verilog/coms.v(148[4] 304[11])
    defparam select_812_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_810_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1417 (.I0(n26123), .I1(n61557), .I2(\data_out_frame[15] [3]), 
            .I3(\data_out_frame[17] [5]), .O(n59360));
    defparam i3_4_lut_adj_1417.LUT_INIT = 16'h9669;
    SB_LUT4 i15881_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n30288));
    defparam i15881_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15884_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n30291));
    defparam i15884_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1418 (.I0(n54982), .I1(n59360), .I2(GND_net), 
            .I3(GND_net), .O(n59361));
    defparam i1_2_lut_adj_1418.LUT_INIT = 16'h6666;
    SB_LUT4 i15887_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n30294));
    defparam i15887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1419 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[17] [3]), 
            .I2(n59784), .I3(\data_out_frame[19] [4]), .O(n30_adj_5753));
    defparam i11_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i15890_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n30297));
    defparam i15890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1420 (.I0(\data_out_frame[19] [3]), .I1(n30_adj_5753), 
            .I2(\data_out_frame[19] [5]), .I3(n59361), .O(n34));
    defparam i15_4_lut_adj_1420.LUT_INIT = 16'h9669;
    SB_LUT4 i15893_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n30300));
    defparam i15893_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15896_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n30303));
    defparam i15896_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15900_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n30307));
    defparam i15900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15903_3_lut_4_lut (.I0(n8_adj_11), .I1(n59077), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n30310));
    defparam i15903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1421 (.I0(n59811), .I1(n59100), .I2(n59635), 
            .I3(n54161), .O(n32_adj_5754));
    defparam i13_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1422 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[17] [4]), .I3(\data_out_frame[17] [1]), 
            .O(n33_adj_5755));
    defparam i14_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1423 (.I0(n59404), .I1(n26137), .I2(\data_out_frame[17] [7]), 
            .I3(\data_out_frame[18] [0]), .O(n31_adj_5756));
    defparam i12_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1424 (.I0(\FRAME_MATCHER.i_31__N_2637 ), .I1(\FRAME_MATCHER.i_31__N_2641 ), 
            .I2(n59060), .I3(LED_c), .O(n27759));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1424.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1425 (.I0(\FRAME_MATCHER.i_31__N_2637 ), .I1(\FRAME_MATCHER.i_31__N_2641 ), 
            .I2(\FRAME_MATCHER.i_31__N_2643 ), .I3(GND_net), .O(n3942));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1425.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_336_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_11));   // verilog/coms.v(157[7:23])
    defparam equal_336_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i18_4_lut_adj_1426 (.I0(n31_adj_5756), .I1(n33_adj_5755), .I2(n32_adj_5754), 
            .I3(n34), .O(n59833));
    defparam i18_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [5]), .I3(n59625), .O(n6_adj_5757));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 equal_343_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_12));   // verilog/coms.v(157[7:23])
    defparam equal_343_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_349_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5758));   // verilog/coms.v(158[12:15])
    defparam equal_349_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_341_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5759));   // verilog/coms.v(158[12:15])
    defparam equal_341_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1427 (.I0(n1519), .I1(n1516), .I2(n59347), 
            .I3(\data_out_frame[12] [4]), .O(n27181));
    defparam i2_3_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(n26113), .I1(n59404), .I2(n10_adj_5760), 
            .I3(\data_out_frame[18] [7]), .O(n54734));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59157));
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h6666;
    SB_LUT4 i29643_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43937));
    defparam i29643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1429 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(\data_out_frame[14] [5]), .I3(n59235), .O(n59196));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1430 (.I0(n69906), .I1(n59663), .I2(n59690), 
            .I3(n59150), .O(n22_adj_5761));
    defparam i9_4_lut_adj_1430.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1431 (.I0(n54994), .I1(n22_adj_5761), .I2(n16_adj_5762), 
            .I3(n59811), .O(n24_adj_5763));
    defparam i11_4_lut_adj_1431.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54646 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n70843));
    defparam byte_transmit_counter_0__bdd_4_lut_54646.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(n26509), .I3(n26087), .O(n1312));
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[7] [4]), .O(n59593));
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1434 (.I0(n26693), .I1(n24_adj_5763), .I2(n20_adj_5764), 
            .I3(\data_out_frame[23] [2]), .O(n54991));
    defparam i12_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1435 (.I0(n26113), .I1(n59635), .I2(n27181), 
            .I3(\data_out_frame[17] [0]), .O(n59606));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(n26113), .I1(n59635), .I2(\data_out_frame[17] [2]), 
            .I3(\data_out_frame[17] [0]), .O(n26137));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1437 (.I0(n59522), .I1(n54991), .I2(n59455), 
            .I3(n59157), .O(n59583));
    defparam i2_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5631));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1438 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n59629));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1438.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_221_i3_2_lut (.I0(n59583), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5739));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_221_i3_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_810_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5630));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n59114));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1440 (.I0(n26490), .I1(\data_out_frame[10] [0]), 
            .I2(n54935), .I3(GND_net), .O(n59368));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1440.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1441 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[20] [1]), 
            .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5624));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1441.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26651));
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5623));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i3_4_lut_adj_1443 (.I0(\data_out_frame[18] [4]), .I1(n59675), 
            .I2(n59641), .I3(n26504), .O(n54383));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5622));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_810_Select_8_i2_3_lut (.I0(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\data_out_frame[1][0] ), 
            .I3(GND_net), .O(n2_adj_5620));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(n26490), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[12] [1]), .O(n59793));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1445 (.I0(n54908), .I1(n54383), .I2(n26651), 
            .I3(n6_adj_5765), .O(n25517));
    defparam i4_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5619));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1446 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(n25517), .I3(\data_out_frame[21] [0]), .O(n59455));
    defparam i3_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(n26490), .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[8] [5]), 
            .I3(GND_net), .O(n10_adj_5766));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_222_i3_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5767), .I3(n59458), 
            .O(n3_adj_5738));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i48334_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64508));
    defparam i48334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1447 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26693));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1447.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1448 (.I0(n59225), .I1(n59585), .I2(n26137), 
            .I3(\data_out_frame[21] [4]), .O(n59827));
    defparam i3_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i48335_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64509));
    defparam i48335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1449 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[14] [7]), .I3(n59188), .O(n10_adj_5768));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5617));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i5_3_lut_adj_1450 (.I0(n59598), .I1(n10_adj_5768), .I2(\data_out_frame[10] [5]), 
            .I3(GND_net), .O(n59839));   // verilog/coms.v(76[16:42])
    defparam i5_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5615));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(GND_net), .I3(GND_net), .O(n59479));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(\FRAME_MATCHER.state_31__N_2741 [3]), .I3(GND_net), .O(n2_adj_5614));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1452 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .I2(\data_out_frame[0][2] ), .I3(GND_net), .O(n2_adj_5612));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1452.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3_4_lut_adj_1453 (.I0(\data_out_frame[17] [1]), .I1(n59212), 
            .I2(n59708), .I3(n59479), .O(n59165));
    defparam i3_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(n59225), .I1(n59606), .I2(GND_net), 
            .I3(GND_net), .O(n59781));
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1455 (.I0(\data_out_frame[21] [3]), .I1(n59781), 
            .I2(n59165), .I3(n54734), .O(n54750));
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [7]), 
            .O(n58798));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i3_4_lut_adj_1456 (.I0(\data_out_frame[14] [3]), .I1(n59616), 
            .I2(n59793), .I3(n59629), .O(n59404));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59150));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1458 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26504));
    defparam i1_2_lut_adj_1458.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1459 (.I0(n59619), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[9] [1]), .I3(n59767), .O(n10_adj_5769));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1460 (.I0(n54698), .I1(n54962), .I2(n10_adj_5745), 
            .I3(n59781), .O(n61040));
    defparam i5_3_lut_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1461 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27][6] ), 
            .O(n58799));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1461.LUT_INIT = 16'h5100;
    SB_LUT4 i2_3_lut_adj_1462 (.I0(n26490), .I1(n59270), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n27113));
    defparam i2_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5601));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1463 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [5]), 
            .O(n58800));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1463.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1464 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [4]), 
            .O(n58796));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1464.LUT_INIT = 16'h5100;
    SB_LUT4 i2_4_lut_adj_1465 (.I0(n27113), .I1(n53893), .I2(\data_out_frame[13] [5]), 
            .I3(n25546), .O(n54003));
    defparam i2_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1466 (.I0(\data_out_frame[17] [0]), .I1(n27181), 
            .I2(n59833), .I3(GND_net), .O(n59663));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1467 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [3]), 
            .O(n58801));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1467.LUT_INIT = 16'h5100;
    SB_LUT4 i3_2_lut_adj_1468 (.I0(n59808), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5770));
    defparam i3_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1469 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [2]), 
            .O(n58802));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1469.LUT_INIT = 16'h5100;
    SB_LUT4 i5_4_lut_adj_1470 (.I0(\data_out_frame[13] [1]), .I1(n59776), 
            .I2(n27029), .I3(\data_out_frame[11] [0]), .O(n13_adj_5771));
    defparam i5_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1471 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [1]), 
            .O(n58803));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1471.LUT_INIT = 16'h5100;
    SB_LUT4 select_810_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5600));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1472 (.I0(\data_out_frame[5] [4]), .I1(n10_adj_5772), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [2]), .O(n59222));   // verilog/coms.v(74[16:62])
    defparam i5_3_lut_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1473 (.I0(n13_adj_5771), .I1(n11_adj_5770), .I2(n32_adj_5773), 
            .I3(n61823), .O(n61557));
    defparam i7_4_lut_adj_1473.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1474 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[27] [0]), 
            .O(n58804));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1474.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1475 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [7]), 
            .O(n58805));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1475.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_adj_1476 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n59776));
    defparam i1_2_lut_adj_1476.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1477 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59162));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1477.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1478 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26][6] ), 
            .O(n58806));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1478.LUT_INIT = 16'h5100;
    SB_LUT4 select_810_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5599));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5774));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1480 (.I0(n59776), .I1(n59669), .I2(\data_out_frame[10] [7]), 
            .I3(n6_adj_5775), .O(n61686));   // verilog/coms.v(88[17:63])
    defparam i4_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1481 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [5]), 
            .O(n58807));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1481.LUT_INIT = 16'h5100;
    SB_LUT4 select_810_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5598));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1482 (.I0(n59327), .I1(n61686), .I2(n59598), 
            .I3(n6_adj_5774), .O(n59808));
    defparam i4_4_lut_adj_1482.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1483 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [4]), 
            .O(n58797));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1483.LUT_INIT = 16'h5100;
    SB_LUT4 select_810_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5597));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59401));
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1485 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [0]), 
            .O(n58808));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1485.LUT_INIT = 16'h5100;
    SB_LUT4 i5_4_lut_adj_1486 (.I0(n1130), .I1(n26660), .I2(\data_out_frame[9] [0]), 
            .I3(\data_out_frame[13] [2]), .O(n12_adj_5776));   // verilog/coms.v(77[16:43])
    defparam i5_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1487 (.I0(n26094), .I1(n12_adj_5776), .I2(\data_out_frame[6] [6]), 
            .I3(\data_out_frame[10] [6]), .O(n59261));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59350));
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h6666;
    SB_LUT4 i13999_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3942), 
            .I3(\FRAME_MATCHER.i_31__N_2636 ), .O(n28405));   // verilog/coms.v(158[12:15])
    defparam i13999_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i5_3_lut_4_lut_adj_1489 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(n10_adj_5777), .I3(n32_adj_5773), .O(n54753));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i48320_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64494));
    defparam i48320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48319_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64493));
    defparam i48319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1490 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [1]), 
            .O(n58809));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1490.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1491 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[19] [1]), 
            .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5582));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1491.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1492 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [2]), 
            .O(n58810));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1492.LUT_INIT = 16'h5100;
    SB_LUT4 i9_4_lut_adj_1493 (.I0(\data_out_frame[7] [0]), .I1(n59267), 
            .I2(n26660), .I3(\data_out_frame[4] [5]), .O(n24_adj_5778));
    defparam i9_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1494 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2638 ), .I3(\data_out_frame[26] [3]), 
            .O(n58795));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1494.LUT_INIT = 16'h5100;
    SB_LUT4 i11_4_lut_adj_1495 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(n59154), .I3(n1130), .O(n26_adj_5779));
    defparam i11_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1496 (.I0(\data_out_frame[6] [6]), .I1(n59222), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n59154));
    defparam i1_2_lut_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5581));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i10_4_lut_adj_1497 (.I0(\data_out_frame[7] [1]), .I1(n59327), 
            .I2(n59593), .I3(n59202), .O(n25_adj_5780));
    defparam i10_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5580));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_150_i2_4_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5578));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_150_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5577));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5576));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1498 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[4] [3]), .O(n32_adj_5773));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1499 (.I0(n59181), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[9] [6]), .I3(n26516), .O(n14_adj_5781));
    defparam i6_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5575));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16304_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30711));   // verilog/coms.v(130[12] 305[6])
    defparam i16304_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5574));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16325_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30732));   // verilog/coms.v(130[12] 305[6])
    defparam i16325_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1500 (.I0(\data_out_frame[7] [5]), .I1(n27_adj_5782), 
            .I2(n25_adj_5780), .I3(n26_adj_5779), .O(n9));
    defparam i1_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5573));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15620_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n30027));   // verilog/coms.v(130[12] 305[6])
    defparam i15620_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1501 (.I0(n9), .I1(n14_adj_5781), .I2(n59114), 
            .I3(\data_out_frame[9] [1]), .O(n54935));
    defparam i7_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5572));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16334_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30741));   // verilog/coms.v(130[12] 305[6])
    defparam i16334_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5783));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5571));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16333_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30740));   // verilog/coms.v(130[12] 305[6])
    defparam i16333_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1503 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(n1191), .I3(n6_adj_5783), .O(n59188));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1504 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[17] [6]), 
            .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5570));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1504.LUT_INIT = 16'ha088;
    SB_LUT4 i6_4_lut_adj_1505 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(n54935), .I3(\data_out_frame[4] [1]), .O(n14_adj_5784));
    defparam i6_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i16332_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30739));   // verilog/coms.v(130[12] 305[6])
    defparam i16332_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5569));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1506 (.I0(n59350), .I1(n14_adj_5784), .I2(n10_adj_5766), 
            .I3(\data_out_frame[6] [3]), .O(n61823));
    defparam i7_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i16331_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30738));   // verilog/coms.v(130[12] 305[6])
    defparam i16331_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5568));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5567));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16330_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30737));   // verilog/coms.v(130[12] 305[6])
    defparam i16330_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5566));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16329_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30736));   // verilog/coms.v(130[12] 305[6])
    defparam i16329_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1507 (.I0(n59666), .I1(n61823), .I2(n59188), 
            .I3(\data_out_frame[12] [6]), .O(n14_adj_5785));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1507.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5565));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16328_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30735));   // verilog/coms.v(130[12] 305[6])
    defparam i16328_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5564));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16327_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30734));   // verilog/coms.v(130[12] 305[6])
    defparam i16327_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5563));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1508 (.I0(n59669), .I1(n59368), .I2(\data_out_frame[8] [3]), 
            .I3(\data_out_frame[12] [7]), .O(n13_adj_5786));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i16324_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30731));   // verilog/coms.v(130[12] 305[6])
    defparam i16324_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5562));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1509 (.I0(n13_adj_5786), .I1(\data_out_frame[13] [0]), 
            .I2(n14_adj_5785), .I3(GND_net), .O(n53905));
    defparam i1_3_lut_adj_1509.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1510 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n59666));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1510.LUT_INIT = 16'h9696;
    SB_LUT4 i16323_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30730));   // verilog/coms.v(130[12] 305[6])
    defparam i16323_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5561));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1511 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[6] [2]), .O(n59598));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5560));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16322_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30729));   // verilog/coms.v(130[12] 305[6])
    defparam i16322_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_810_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5559));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1512 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59267));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1512.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5558));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27086));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i16321_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30728));   // verilog/coms.v(130[12] 305[6])
    defparam i16321_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1514 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[8] [7]), .I3(n59218), .O(n59619));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1515 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(n59222), .I3(GND_net), .O(n26768));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1515.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5555));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59181));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1517 (.I0(\data_out_frame[9] [2]), .I1(n10_adj_5787), 
            .I2(n26509), .I3(n27113), .O(n59675));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1518 (.I0(\data_out_frame[9] [2]), .I1(n10_adj_5787), 
            .I2(n26509), .I3(n53893), .O(n59431));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1519 (.I0(n59222), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n59153));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1519.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1520 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n27029));
    defparam i2_2_lut_3_lut_adj_1520.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n59767));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i12_3_lut_4_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(n59344), .I3(n24_adj_5778), .O(n27_adj_5782));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1522 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n59254), .I3(GND_net), .O(n59641));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1522.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1523 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n59675), .I3(GND_net), .O(n6_adj_5746));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16320_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30727));   // verilog/coms.v(130[12] 305[6])
    defparam i16320_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16319_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30726));   // verilog/coms.v(130[12] 305[6])
    defparam i16319_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1524 (.I0(n59154), .I1(n26768), .I2(n1130), .I3(n59767), 
            .O(n10_adj_5787));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i16318_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30725));   // verilog/coms.v(130[12] 305[6])
    defparam i16318_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i23650_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n23164), .I3(GND_net), .O(n30008));
    defparam i23650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1525 (.I0(\data_out_frame[15] [5]), .I1(n54753), 
            .I2(n26681), .I3(GND_net), .O(n54945));
    defparam i1_2_lut_3_lut_adj_1525.LUT_INIT = 16'h9696;
    SB_LUT4 i24127_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1]_c [0]), 
            .I2(n23230), .I3(GND_net), .O(n30009));
    defparam i24127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1526 (.I0(\data_out_frame[15] [5]), .I1(n54753), 
            .I2(n26123), .I3(\data_out_frame[15] [4]), .O(n54982));
    defparam i1_2_lut_3_lut_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1527 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n6_adj_5765));
    defparam i1_2_lut_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i16317_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30724));   // verilog/coms.v(130[12] 305[6])
    defparam i16317_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1528 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(n54698), .I3(\data_out_frame[18] [5]), .O(n54916));
    defparam i2_3_lut_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1529 (.I0(n59181), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[13] [4]), .I3(n59619), .O(n10_adj_5777));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16316_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30723));   // verilog/coms.v(130[12] 305[6])
    defparam i16316_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1530 (.I0(\data_out_frame[5] [0]), .I1(n1191), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[5] [5]), .O(n10_adj_5772));   // verilog/coms.v(74[16:62])
    defparam i4_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i16315_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30722));   // verilog/coms.v(130[12] 305[6])
    defparam i16315_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16314_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30721));   // verilog/coms.v(130[12] 305[6])
    defparam i16314_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1531 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n59324));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1531.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1532 (.I0(n54753), .I1(n59431), .I2(GND_net), 
            .I3(GND_net), .O(n26970));
    defparam i1_2_lut_adj_1532.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1533 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(n59153), .I3(GND_net), .O(n14_adj_5788));
    defparam i5_3_lut_adj_1533.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1534 (.I0(n59666), .I1(\data_out_frame[13] [3]), 
            .I2(n26768), .I3(n59324), .O(n15_adj_5789));
    defparam i6_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1535 (.I0(\data_out_frame[19] [3]), .I1(n59827), 
            .I2(\data_out_frame[21] [5]), .I3(GND_net), .O(n54694));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1535.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1536 (.I0(\data_out_frame[19] [3]), .I1(n59827), 
            .I2(\data_out_frame[23] [5]), .I3(n54750), .O(n61148));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1537 (.I0(\data_out_frame[23] [4]), .I1(n54750), 
            .I2(\data_out_frame[23] [6]), .I3(GND_net), .O(n59542));
    defparam i1_2_lut_3_lut_adj_1537.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1538 (.I0(\data_out_frame[23] [4]), .I1(n54750), 
            .I2(n59455), .I3(GND_net), .O(n6_adj_5767));
    defparam i2_2_lut_3_lut_adj_1538.LUT_INIT = 16'h9696;
    SB_LUT4 i16292_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n30699));
    defparam i16292_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8_4_lut_adj_1539 (.I0(n15_adj_5789), .I1(\data_out_frame[9] [1]), 
            .I2(n14_adj_5788), .I3(\data_out_frame[11] [2]), .O(n26681));
    defparam i8_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1540 (.I0(n59641), .I1(n1519), .I2(n59261), 
            .I3(\data_out_frame[11] [5]), .O(n44_adj_5790));   // verilog/coms.v(74[16:27])
    defparam i18_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i16338_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n30745));
    defparam i16338_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16_4_lut_adj_1541 (.I0(\data_out_frame[14] [4]), .I1(n59836), 
            .I2(n53905), .I3(n59347), .O(n42_adj_5791));   // verilog/coms.v(74[16:27])
    defparam i16_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i15391_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29798));
    defparam i15391_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_1542 (.I0(n26681), .I1(n26970), .I2(\data_out_frame[11] [4]), 
            .I3(n26113), .O(n43_adj_5792));   // verilog/coms.v(74[16:27])
    defparam i17_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1543 (.I0(n1835), .I1(\data_out_frame[15] [5]), 
            .I2(n59401), .I3(\data_out_frame[14] [7]), .O(n41_adj_5793));   // verilog/coms.v(74[16:27])
    defparam i15_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1544 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[8] [7]), .O(n26660));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i15388_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29795));
    defparam i15388_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16313_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30720));   // verilog/coms.v(130[12] 305[6])
    defparam i16313_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14_4_lut_adj_1545 (.I0(n59808), .I1(n59162), .I2(\data_out_frame[11] [7]), 
            .I3(\data_out_frame[15] [4]), .O(n40_adj_5794));   // verilog/coms.v(74[16:27])
    defparam i14_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i15385_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29792));
    defparam i15385_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15381_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29788));
    defparam i15381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16451_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n30858));
    defparam i16451_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19_4_lut_adj_1546 (.I0(n27086), .I1(\data_out_frame[14] [3]), 
            .I2(n61557), .I3(n54003), .O(n45_adj_5795));   // verilog/coms.v(74[16:27])
    defparam i19_4_lut_adj_1546.LUT_INIT = 16'h9669;
    SB_LUT4 i15378_3_lut_4_lut (.I0(n44625), .I1(n59083), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29785));
    defparam i15378_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i24_4_lut_adj_1547 (.I0(n41_adj_5793), .I1(n43_adj_5792), .I2(n42_adj_5791), 
            .I3(n44_adj_5790), .O(n50_adj_5796));   // verilog/coms.v(74[16:27])
    defparam i24_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n45_adj_5795), .I1(\data_out_frame[10] [5]), 
            .I2(n40_adj_5794), .I3(\data_out_frame[11] [6]), .O(n49));   // verilog/coms.v(74[16:27])
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1548 (.I0(n54222), .I1(n54383), .I2(n54900), 
            .I3(\data_out_frame[20] [0]), .O(n61790));
    defparam i2_3_lut_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 n70843_bdd_4_lut (.I0(n70843), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n70846));
    defparam n70843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_2_lut_3_lut (.I0(n54222), .I1(n54383), .I2(\data_out_frame[16] [1]), 
            .I3(GND_net), .O(n16_adj_5762));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1549 (.I0(\data_out_frame[20] [4]), .I1(n59185), 
            .I2(\data_out_frame[20] [5]), .I3(n59273), .O(n54222));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1550 (.I0(\data_out_frame[20] [4]), .I1(n59185), 
            .I2(\data_out_frame[22] [7]), .I3(GND_net), .O(n59690));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1550.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1551 (.I0(n49), .I1(n54945), .I2(n50_adj_5796), 
            .I3(\data_out_frame[16] [0]), .O(n59374));
    defparam i2_4_lut_adj_1551.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1552 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(n61255), .I3(n55014), .O(n54943));
    defparam i2_3_lut_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1553 (.I0(n26504), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[16] [7]), .I3(\data_out_frame[16] [1]), 
            .O(n59610));   // verilog/coms.v(88[17:28])
    defparam i2_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1554 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n59185));
    defparam i1_2_lut_3_lut_adj_1554.LUT_INIT = 16'h9696;
    SB_LUT4 i16312_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30719));   // verilog/coms.v(130[12] 305[6])
    defparam i16312_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1555 (.I0(\data_out_frame[15] [4]), .I1(n26123), 
            .I2(n26681), .I3(GND_net), .O(n26523));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1555.LUT_INIT = 16'h9696;
    SB_LUT4 i16311_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30718));   // verilog/coms.v(130[12] 305[6])
    defparam i16311_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut_adj_1556 (.I0(n59196), .I1(n59374), .I2(n54994), 
            .I3(GND_net), .O(n8_adj_5797));   // verilog/coms.v(88[17:28])
    defparam i3_3_lut_adj_1556.LUT_INIT = 16'h9696;
    SB_LUT4 i15636_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[1]), 
            .I3(\data_in_frame[1][1] ), .O(n30043));
    defparam i15636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15612_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[0]), 
            .I3(\data_in_frame[1]_c [0]), .O(n30019));
    defparam i15612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15709_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n30116));
    defparam i15709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1557 (.I0(n59610), .I1(n59150), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5798));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i15702_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n30109));
    defparam i15702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16310_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30717));   // verilog/coms.v(130[12] 305[6])
    defparam i16310_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15688_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n30095));
    defparam i15688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1558 (.I0(\data_out_frame[18] [6]), .I1(n7_adj_5798), 
            .I2(\data_out_frame[18] [7]), .I3(n8_adj_5797), .O(n59784));
    defparam i2_4_lut_adj_1558.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1559 (.I0(\data_out_frame[4] [0]), .I1(n59118), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[6] [1]), .O(n59327));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i15685_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n30092));
    defparam i15685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n59347));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h6666;
    SB_LUT4 i16309_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30716));   // verilog/coms.v(130[12] 305[6])
    defparam i16309_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15656_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n30063));
    defparam i15656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16308_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30715));   // verilog/coms.v(130[12] 305[6])
    defparam i16308_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15643_3_lut_4_lut (.I0(n8_adj_10), .I1(n59077), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n30050));
    defparam i15643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16307_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30714));   // verilog/coms.v(130[12] 305[6])
    defparam i16307_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 equal_339_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_10));   // verilog/coms.v(157[7:23])
    defparam equal_339_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut_3_lut_adj_1561 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_3_lut_adj_1561.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(\data_out_frame[12] [4]), .I1(n1516), 
            .I2(GND_net), .I3(GND_net), .O(n59632));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1563 (.I0(\data_out_frame[16] [7]), .I1(n59196), 
            .I2(GND_net), .I3(GND_net), .O(n59708));
    defparam i1_2_lut_adj_1563.LUT_INIT = 16'h6666;
    SB_LUT4 i15417_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29824));
    defparam i15417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1564 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [1]), .I3(GND_net), .O(n59669));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1564.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1565 (.I0(n59606), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[19] [1]), .I3(n59708), .O(n10_adj_5760));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 i16306_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30713));   // verilog/coms.v(130[12] 305[6])
    defparam i16306_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15414_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[6]), 
            .I3(\data_in_frame[16]_c [6]), .O(n29821));
    defparam i15414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15411_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[5]), 
            .I3(\data_in_frame[16]_c [5]), .O(n29818));
    defparam i15411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15408_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[4]), 
            .I3(\data_in_frame[16]_c [4]), .O(n29815));
    defparam i15408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15403_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[3]), 
            .I3(\data_in_frame[16]_c [3]), .O(n29810));
    defparam i15403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15400_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[2]), 
            .I3(\data_in_frame[16]_c [2]), .O(n29807));
    defparam i15400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23651_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6][4] ), 
            .I2(n23164), .I3(GND_net), .O(n30069));
    defparam i23651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23836_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6]_c [5]), 
            .I2(n23164), .I3(GND_net), .O(n30070));
    defparam i23836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23025_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(\data_in_frame[16]_c [1]), 
            .I3(rx_data[1]), .O(n29804));
    defparam i23025_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i23837_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6]_c [6]), 
            .I2(n23164), .I3(GND_net), .O(n30071));
    defparam i23837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1566 (.I0(\data_out_frame[19] [0]), .I1(n54734), 
            .I2(GND_net), .I3(GND_net), .O(n54962));
    defparam i1_2_lut_adj_1566.LUT_INIT = 16'h6666;
    SB_LUT4 i15394_3_lut_4_lut (.I0(n8), .I1(n59047), .I2(rx_data[0]), 
            .I3(\data_in_frame[16]_c [0]), .O(n29801));
    defparam i15394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71077_bdd_4_lut (.I0(n71077), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n64549));
    defparam n71077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1567 (.I0(n54908), .I1(n59784), .I2(n59610), 
            .I3(n59374), .O(n54698));
    defparam i3_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i16305_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30712));   // verilog/coms.v(130[12] 305[6])
    defparam i16305_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1568 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n59232));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1568.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1569 (.I0(\data_out_frame[8] [1]), .I1(n59629), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[10] [2]), .O(n12_adj_5799));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1569.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1570 (.I0(\data_out_frame[5] [7]), .I1(n12_adj_5799), 
            .I2(\data_out_frame[12] [3]), .I3(n59232), .O(n59235));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 i16326_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30733));   // verilog/coms.v(130[12] 305[6])
    defparam i16326_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1571 (.I0(n26490), .I1(\data_out_frame[10] [0]), 
            .I2(n54935), .I3(\data_out_frame[10] [5]), .O(n6_adj_5775));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_4_lut_adj_1571.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1572 (.I0(\data_out_frame[14] [4]), .I1(n59235), 
            .I2(GND_net), .I3(GND_net), .O(n59635));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1573 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(n59232), .I3(n6_adj_5757), .O(n26113));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1574 (.I0(\data_out_frame[7] [1]), .I1(n26509), 
            .I2(n10_adj_5769), .I3(n27029), .O(n25546));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1574.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5550));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1575 (.I0(n54698), .I1(\data_out_frame[19] [0]), 
            .I2(n54734), .I3(\data_out_frame[21] [2]), .O(n59522));
    defparam i1_2_lut_3_lut_4_lut_adj_1575.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1576 (.I0(n1312), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n59270));
    defparam i2_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 i48328_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64502));
    defparam i48328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48329_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64503));
    defparam i48329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48353_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64527));
    defparam i48353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48352_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64526));
    defparam i48352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(n61754), .I1(n59318), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n53959));
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1578 (.I0(n61754), .I1(n59318), .I2(n54222), 
            .I3(GND_net), .O(n59723));
    defparam i1_2_lut_3_lut_adj_1578.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1579 (.I0(\data_out_frame[12] [0]), .I1(n59793), 
            .I2(n59114), .I3(n59270), .O(n12_adj_5800));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64420), .I3(n64418), 
            .O(n7_adj_5801));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64417), .I3(n64415), 
            .O(n7_adj_5802));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i6_4_lut_adj_1580 (.I0(\data_out_frame[7] [6]), .I1(n12_adj_5800), 
            .I2(\data_out_frame[14] [2]), .I3(n59625), .O(n59254));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64426), .I3(n64424), 
            .O(n7_adj_5803));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n64450), .I3(n64448), 
            .O(n7));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i10_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), .I1(\byte_transmit_counter[1] ), 
            .I2(n64453), .I3(n64451), .O(n7_adj_5685));   // verilog/coms.v(109[34:55])
    defparam i10_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_4_lut_adj_1581 (.I0(\data_out_frame[15] [0]), .I1(n59598), 
            .I2(n10_adj_5768), .I3(\data_out_frame[10] [5]), .O(n59212));
    defparam i1_2_lut_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1582 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n59225));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1582.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1583 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(n53905), .I3(GND_net), .O(n59585));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_3_lut_adj_1583.LUT_INIT = 16'h9696;
    SB_LUT4 i15856_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n30263));
    defparam i15856_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15859_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n30266));
    defparam i15859_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15862_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n30269));
    defparam i15862_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15865_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n30272));
    defparam i15865_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15869_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n30276));
    defparam i15869_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15872_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n30279));
    defparam i15872_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1584 (.I0(\data_out_frame[14] [1]), .I1(n26490), 
            .I2(GND_net), .I3(GND_net), .O(n59836));
    defparam i1_2_lut_adj_1584.LUT_INIT = 16'h6666;
    SB_LUT4 i15875_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n30282));
    defparam i15875_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15878_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59077), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n30285));
    defparam i15878_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1585 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59344));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1586 (.I0(n26113), .I1(\data_out_frame[14] [4]), 
            .I2(n59235), .I3(n59254), .O(n54908));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\data_out_frame[7] [1]), .I1(n26509), 
            .I2(GND_net), .I3(GND_net), .O(n26954));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h6666;
    SB_LUT4 i7_3_lut_4_lut_adj_1588 (.I0(n54734), .I1(n54908), .I2(\data_out_frame[21] [1]), 
            .I3(\data_out_frame[23] [1]), .O(n20_adj_5764));
    defparam i7_3_lut_4_lut_adj_1588.LUT_INIT = 16'h6996;
    SB_LUT4 i30326_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n44625));
    defparam i30326_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_2_lut_3_lut_adj_1589 (.I0(\data_out_frame[22] [4]), .I1(n54966), 
            .I2(n59473), .I3(GND_net), .O(n6_adj_5683));
    defparam i2_2_lut_3_lut_adj_1589.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1590 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n55026), .I3(GND_net), .O(n59273));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1590.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1591 (.I0(n1519), .I1(n1516), .I2(\data_out_frame[7] [6]), 
            .I3(\data_out_frame[11] [7]), .O(n14_adj_5805));
    defparam i1_2_lut_3_lut_4_lut_adj_1591.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59218));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1593 (.I0(\data_out_frame[20] [2]), .I1(n61719), 
            .I2(\data_out_frame[22] [3]), .I3(n59560), .O(n54397));
    defparam i2_3_lut_4_lut_adj_1593.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1594 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26516));
    defparam i1_2_lut_adj_1594.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1595 (.I0(\data_out_frame[11] [5]), .I1(n26516), 
            .I2(n59218), .I3(\data_out_frame[4] [5]), .O(n12_adj_5806));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1596 (.I0(\data_out_frame[6] [7]), .I1(n12_adj_5806), 
            .I2(n1312), .I3(n26954), .O(n53893));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1596.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5541));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1597 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[8] [0]), .I3(n6_adj_5750), .O(n59202));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1597.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1598 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n59625));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1598.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1599 (.I0(reset), .I1(n3942), .I2(n161), 
            .I3(n10_adj_5758), .O(n59077));
    defparam i1_2_lut_3_lut_4_lut_adj_1599.LUT_INIT = 16'hffbf;
    SB_LUT4 select_810_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54641 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[20] [2]), .I2(\data_out_frame[21] [2]), 
            .I3(byte_transmit_counter_c[4]), .O(n70837));
    defparam byte_transmit_counter_0__bdd_4_lut_54641.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1600 (.I0(reset), .I1(n3942), .I2(n161), 
            .I3(n10_adj_5759), .O(n59083));
    defparam i1_2_lut_3_lut_4_lut_adj_1600.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_1601 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n59967), .O(n59093));
    defparam i1_2_lut_4_lut_adj_1601.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1602 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [3]), 
            .I2(\data_out_frame[18] [4]), .I3(GND_net), .O(n59811));
    defparam i1_2_lut_3_lut_adj_1602.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1603 (.I0(n3942), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n57), .I3(reset), .O(n59047));
    defparam i2_3_lut_4_lut_adj_1603.LUT_INIT = 16'hffdf;
    SB_LUT4 n70837_bdd_4_lut (.I0(n70837), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[4] [2]), .I3(byte_transmit_counter_c[4]), 
            .O(n70840));
    defparam n70837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1604 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5697), 
            .I2(n42164), .I3(n3942), .O(n28719));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1604.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1605 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_5697), 
            .I2(n59967), .I3(n10_adj_5759), .O(n28745));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1605.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1606 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n6_adj_5633));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1606.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1607 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(n24221), .I3(GND_net), .O(n18_adj_5648));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1608 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1][1] ), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n59354));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1608.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1609 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [5]), 
            .I2(n59625), .I3(GND_net), .O(n59790));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1609.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1610 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8] [1]), .I3(\data_out_frame[10] [4]), .O(n59398));
    defparam i3_4_lut_adj_1610.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1611 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1][1] ), 
            .I2(\data_in_frame[1]_c [0]), .I3(n59602), .O(n26302));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 i15928_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n30335));
    defparam i15928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15925_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n30332));
    defparam i15925_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15922_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n30329));
    defparam i15922_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1612 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59613));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1612.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1613 (.I0(\FRAME_MATCHER.i[4] ), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(\FRAME_MATCHER.i[3] ), 
            .O(n57));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1613.LUT_INIT = 16'h0008;
    SB_LUT4 i15919_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n30326));
    defparam i15919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54636 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter_c[4]), .O(n70831));
    defparam byte_transmit_counter_0__bdd_4_lut_54636.LUT_INIT = 16'he4aa;
    SB_LUT4 i15915_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n30322));
    defparam i15915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1614 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59787));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1614.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1615 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n59118));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1615.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15912_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n30319));
    defparam i15912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(n5), .O(n59174));   // verilog/coms.v(169[9:87])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15909_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n30316));
    defparam i15909_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15906_3_lut_4_lut (.I0(n8_adj_12), .I1(n59077), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n30313));
    defparam i15906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1616 (.I0(\data_in_frame[2] [7]), .I1(n26302), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n26617));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_3_lut_adj_1616.LUT_INIT = 16'h9696;
    SB_LUT4 n70831_bdd_4_lut (.I0(n70831), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[6] [2]), .I3(byte_transmit_counter_c[4]), 
            .O(n70834));
    defparam n70831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1617 (.I0(\data_in_frame[2] [7]), .I1(n26302), 
            .I2(\data_in_frame[2] [6]), .I3(n10_adj_5645), .O(n59644));   // verilog/coms.v(80[16:27])
    defparam i5_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1618 (.I0(\data_in_frame[1] [4]), .I1(n59539), 
            .I2(n59573), .I3(n59569), .O(n59761));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i21431_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n23230), .I3(GND_net), .O(n30122));
    defparam i21431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1619 (.I0(\data_out_frame[4] [0]), .I1(n59613), 
            .I2(n59202), .I3(\data_out_frame[10] [2]), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1620 (.I0(n59118), .I1(n59787), .I2(n59613), 
            .I3(n59398), .O(n1519));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1620.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1621 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(n59590), .O(n6_adj_5629));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1621.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59616));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'h6666;
    SB_LUT4 select_810_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1623 (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n7_adj_5743));
    defparam i2_2_lut_3_lut_adj_1623.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1624 (.I0(n3942), .I1(n42164), .I2(n43937), 
            .I3(\FRAME_MATCHER.i [0]), .O(n28723));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1624.LUT_INIT = 16'hff7f;
    SB_LUT4 i9_4_lut_adj_1625 (.I0(\data_out_frame[13] [7]), .I1(n59398), 
            .I2(n59790), .I3(n26094), .O(n22_adj_5807));
    defparam i9_4_lut_adj_1625.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(n26753), .I1(n59168), .I2(Kp_23__N_1007), 
            .I3(\data_in_frame[8][7] ), .O(n7_adj_5660));   // verilog/coms.v(78[16:43])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1626 (.I0(n26753), .I1(n59168), .I2(Kp_23__N_1007), 
            .I3(n53918), .O(n54912));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n70714), .I2(n64549), .I3(byte_transmit_counter_c[3]), 
            .O(n70825));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 select_810_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1627 (.I0(n26753), .I1(n59168), .I2(Kp_23__N_1007), 
            .I3(n59650), .O(n22_adj_5583));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1628 (.I0(n54030), .I1(\data_in_frame[13] [5]), 
            .I2(n26376), .I3(GND_net), .O(n6_adj_5610));
    defparam i1_2_lut_3_lut_adj_1628.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1629 (.I0(n54030), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[13] [6]), .I3(n59818), .O(n59729));
    defparam i2_3_lut_4_lut_adj_1629.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1630 (.I0(n59446), .I1(n59638), .I2(n7_adj_5660), 
            .I3(n26376), .O(n55066));
    defparam i1_2_lut_4_lut_adj_1630.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1631 (.I0(n59446), .I1(n59638), .I2(n7_adj_5660), 
            .I3(n26806), .O(n59711));
    defparam i1_2_lut_4_lut_adj_1631.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1632 (.I0(n59446), .I1(n59638), .I2(n7_adj_5660), 
            .I3(\data_in_frame[16]_c [0]), .O(n59818));
    defparam i1_2_lut_4_lut_adj_1632.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1633 (.I0(n53893), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[12] [0]), .I3(n14_adj_5805), .O(n23_adj_5808));
    defparam i10_4_lut_adj_1633.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(n26707), .I1(n54016), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n54030));
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1635 (.I0(n26707), .I1(n54016), .I2(\data_in_frame[11] [6]), 
            .I3(GND_net), .O(n6_adj_5548));
    defparam i1_2_lut_3_lut_adj_1635.LUT_INIT = 16'h9696;
    SB_LUT4 n70825_bdd_4_lut (.I0(n70825), .I1(n64401), .I2(n64400), .I3(byte_transmit_counter_c[3]), 
            .O(n70828));
    defparam n70825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1636 (.I0(control_mode[1]), .I1(n35592), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1636.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1637 (.I0(control_mode[1]), .I1(n35592), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15_adj_13));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1637.LUT_INIT = 16'hefef;
    SB_LUT4 i12_4_lut_adj_1638 (.I0(n23_adj_5808), .I1(\data_out_frame[10] [2]), 
            .I2(n22_adj_5807), .I3(n59836), .O(n54669));
    defparam i12_4_lut_adj_1638.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(n26113), .I1(n59404), .I2(GND_net), 
            .I3(GND_net), .O(n54994));
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1640 (.I0(n27142), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [4]), .I3(\data_in_frame[9] [3]), .O(n26395));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1640.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1641 (.I0(n27142), .I1(\data_in_frame[9] [2]), 
            .I2(n26189), .I3(n53899), .O(n14_adj_5609));   // verilog/coms.v(76[16:42])
    defparam i5_3_lut_4_lut_adj_1641.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1642 (.I0(n55014), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n59550));
    defparam i1_2_lut_3_lut_adj_1642.LUT_INIT = 16'h6969;
    SB_LUT4 i14395_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n43937), 
            .I2(n59093), .I3(reset), .O(n28801));   // verilog/coms.v(157[7:23])
    defparam i14395_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n71125));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71125_bdd_4_lut (.I0(n71125), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n71128));
    defparam n71125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1643 (.I0(n26848), .I1(n4_adj_5627), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n26455));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1643.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut (.I0(n26848), .I1(n4_adj_5627), .I2(n54912), 
            .I3(n26707), .O(n8_adj_5604));   // verilog/coms.v(77[16:43])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1644 (.I0(n54908), .I1(\data_out_frame[21] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59687));
    defparam i1_2_lut_adj_1644.LUT_INIT = 16'h6666;
    SB_LUT4 equal_337_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_5804));   // verilog/coms.v(157[7:23])
    defparam equal_337_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1645 (.I0(n54659), .I1(\data_in_frame[9] [7]), 
            .I2(n59699), .I3(GND_net), .O(n54986));
    defparam i1_2_lut_3_lut_adj_1645.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1646 (.I0(n54659), .I1(\data_in_frame[9] [7]), 
            .I2(n59251), .I3(GND_net), .O(n10_adj_5606));
    defparam i1_2_lut_3_lut_adj_1646.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54874 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n71119));
    defparam byte_transmit_counter_0__bdd_4_lut_54874.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1647 (.I0(Kp_23__N_1007), .I1(n59264), .I2(\data_in_frame[6]_c [5]), 
            .I3(\data_in_frame[11] [0]), .O(n59107));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1648 (.I0(n59318), .I1(n59449), .I2(n10_adj_5689), 
            .I3(\data_out_frame[15] [7]), .O(n55014));
    defparam i1_2_lut_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_2044_i7_2_lut_4_lut (.I0(Kp_23__N_1007), .I1(n59264), 
            .I2(\data_in_frame[6]_c [5]), .I3(\data_in_frame[8] [6]), .O(n7_adj_5655));   // verilog/coms.v(78[16:43])
    defparam equal_2044_i7_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1649 (.I0(Kp_23__N_1007), .I1(n59264), .I2(\data_in_frame[6]_c [5]), 
            .I3(\data_in_frame[9] [0]), .O(n59300));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15490_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29897));
    defparam i15490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15487_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29894));
    defparam i15487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_810_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1650 (.I0(n59416), .I1(\data_out_frame[20] [7]), 
            .I2(n59522), .I3(n59687), .O(n10_adj_5810));
    defparam i4_4_lut_adj_1650.LUT_INIT = 16'h9669;
    SB_LUT4 i15484_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29891));
    defparam i15484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15481_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29888));
    defparam i15481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15478_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29885));
    defparam i15478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15475_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29882));
    defparam i15475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71119_bdd_4_lut (.I0(n71119), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n71122));
    defparam n71119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54631 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n70819));
    defparam byte_transmit_counter_0__bdd_4_lut_54631.LUT_INIT = 16'he4aa;
    SB_LUT4 i15472_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29879));
    defparam i15472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[19] [0]), 
            .I2(n10_adj_5810), .I3(n54916), .O(n59363));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'h9669;
    SB_LUT4 n70819_bdd_4_lut (.I0(n70819), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n70822));
    defparam n70819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15469_3_lut_4_lut (.I0(n8_adj_5804), .I1(n59047), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29876));
    defparam i15469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14383_3_lut_4_lut (.I0(n10_adj_5759), .I1(n59967), .I2(reset), 
            .I3(n8_adj_11), .O(n59975));
    defparam i14383_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i14385_3_lut_4_lut (.I0(n10_adj_5759), .I1(n59967), .I2(reset), 
            .I3(n8_adj_5804), .O(n28791));
    defparam i14385_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i14391_3_lut_4_lut (.I0(n10_adj_5759), .I1(n59967), .I2(reset), 
            .I3(n8), .O(n59971));
    defparam i14391_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(n26447), .I3(GND_net), .O(n59741));
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1653 (.I0(\data_out_frame[25] [5]), .I1(n59363), 
            .I2(GND_net), .I3(GND_net), .O(n59458));
    defparam i1_2_lut_adj_1653.LUT_INIT = 16'h9999;
    SB_LUT4 i5_3_lut_4_lut_adj_1654 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(n10_adj_5482), .I3(\data_in_frame[15] [2]), .O(n59392));
    defparam i5_3_lut_4_lut_adj_1654.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(n54996), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[22] [0]), .I3(GND_net), .O(n27305));
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1656 (.I0(\data_in_frame[10] [5]), .I1(n26848), 
            .I2(n26365), .I3(GND_net), .O(n59653));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1656.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1657 (.I0(n26523), .I1(n59360), .I2(\data_out_frame[21] [6]), 
            .I3(GND_net), .O(n59749));
    defparam i1_2_lut_3_lut_adj_1657.LUT_INIT = 16'h9696;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1658 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(n59681), .I3(GND_net), .O(n54996));
    defparam i1_2_lut_3_lut_adj_1658.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1659 (.I0(\data_in_frame[6][1] ), .I1(\data_in_frame[6][3] ), 
            .I2(\data_in_frame[6][2] ), .I3(GND_net), .O(n59830));
    defparam i1_2_lut_3_lut_adj_1659.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1660 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6]_c [5]), 
            .I2(\data_in_frame[6]_c [6]), .I3(GND_net), .O(n59168));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1660.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1661 (.I0(n54982), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[17] [6]), .I3(\data_out_frame[19] [7]), 
            .O(n6_adj_5650));
    defparam i1_2_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1662 (.I0(n54982), .I1(n59360), .I2(n59383), 
            .I3(\data_out_frame[19] [7]), .O(n59104));
    defparam i2_3_lut_4_lut_adj_1662.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1663 (.I0(\data_in_frame[10] [5]), .I1(n26848), 
            .I2(\data_in_frame[10] [6]), .I3(GND_net), .O(n59657));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1663.LUT_INIT = 16'h9696;
    SB_LUT4 i16030_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n30437));
    defparam i16030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16027_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n30434));
    defparam i16027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_810_Select_223_i3_4_lut (.I0(n61148), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n59458), .I3(\data_out_frame[25] [6]), .O(n3_adj_5737));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_810_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1664 (.I0(\data_in_frame[2] [3]), .I1(n59410), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[2] [1]), .O(n59533));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 i16024_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n30431));
    defparam i16024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1665 (.I0(\data_out_frame[23] [7]), .I1(\data_out_frame[19] [3]), 
            .I2(n54411), .I3(GND_net), .O(n59824));
    defparam i1_2_lut_3_lut_adj_1665.LUT_INIT = 16'h9696;
    SB_LUT4 i16021_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n30428));
    defparam i16021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16018_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n30425));
    defparam i16018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16015_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n30422));
    defparam i16015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1666 (.I0(\data_in_frame[0] [3]), .I1(n59144), 
            .I2(\data_in_frame[2] [3]), .I3(n59410), .O(Kp_23__N_928));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1667 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(n26296), .O(n59602));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16012_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n30419));
    defparam i16012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16009_3_lut_4_lut (.I0(n8_adj_10), .I1(n59083), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n30416));
    defparam i16009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16055_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n30462));
    defparam i16055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16052_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n30459));
    defparam i16052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1668 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[1][1] ), .O(n59420));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i16049_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n30456));
    defparam i16049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1669 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n59191));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1669.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16046_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n30453));
    defparam i16046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1670 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(n59842), .I3(n59309), .O(n6_adj_5646));
    defparam i2_2_lut_4_lut_adj_1670.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16042_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n30449));
    defparam i16042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16039_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n30446));
    defparam i16039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n58460));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1671 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(n59842), .I3(GND_net), .O(n59705));
    defparam i1_2_lut_3_lut_adj_1671.LUT_INIT = 16'h9696;
    SB_LUT4 i16033_3_lut_4_lut (.I0(n28745), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n30440));
    defparam i16033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1672 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[0] [6]), 
            .I2(n26302), .I3(\data_in_frame[3] [0]), .O(n59281));
    defparam i1_2_lut_4_lut_adj_1672.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1673 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[25] [7]), 
            .I2(n53959), .I3(n59550), .O(n8_adj_5643));
    defparam i1_2_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1674 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(n26339), .O(n59251));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n6_adj_5639));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1676 (.I0(\data_in_frame[6][4] ), .I1(n59830), 
            .I2(\data_in_frame[6][7] ), .I3(\data_in_frame[4] [5]), .O(n6_adj_5638));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1677 (.I0(\data_in_frame[5] [1]), .I1(n59602), 
            .I2(\data_in_frame[3] [1]), .I3(n59354), .O(n6_adj_5635));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1677.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1678 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[2] [7]), 
            .I2(n26302), .I3(\data_in_frame[0] [5]), .O(n59365));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1678.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1679 (.I0(\data_in_frame[6][4] ), .I1(\data_in_frame[4] [2]), 
            .I2(n59357), .I3(Kp_23__N_901), .O(n59264));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1680 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2637 ), 
            .I2(n25927), .I3(\FRAME_MATCHER.i_31__N_2636 ), .O(n4_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1680.LUT_INIT = 16'hfff4;
    SB_LUT4 i5_3_lut_4_lut_adj_1681 (.I0(\data_in_frame[14] [3]), .I1(n55033), 
            .I2(\data_in_frame[18] [7]), .I3(n10_adj_5491), .O(n61489));
    defparam i5_3_lut_4_lut_adj_1681.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1682 (.I0(\data_in_frame[14] [3]), .I1(n55033), 
            .I2(\data_in_frame[16]_c [4]), .I3(n54954), .O(n61452));
    defparam i2_3_lut_4_lut_adj_1682.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54869 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n71113));
    defparam byte_transmit_counter_0__bdd_4_lut_54869.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54622 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n70813));
    defparam byte_transmit_counter_0__bdd_4_lut_54622.LUT_INIT = 16'he4aa;
    SB_LUT4 select_810_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_4_lut (.I0(n26523), .I1(n59360), .I2(n55073), .I3(n59104), 
            .O(n15_adj_5628));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16138_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n30545));
    defparam i16138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16134_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n30541));
    defparam i16134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16129_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30536));
    defparam i16129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16125_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n30532));
    defparam i16125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16122_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30529));
    defparam i16122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1683 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(n59144), .I3(n26786), .O(n26753));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1684 (.I0(n53944), .I1(n59569), .I2(n26809), 
            .I3(GND_net), .O(n59545));
    defparam i1_2_lut_3_lut_adj_1684.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1685 (.I0(n26523), .I1(n59360), .I2(n55073), 
            .I3(GND_net), .O(n59493));
    defparam i1_2_lut_3_lut_adj_1685.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1686 (.I0(\data_out_frame[17] [3]), .I1(n61557), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n8_adj_5618));
    defparam i1_2_lut_3_lut_adj_1686.LUT_INIT = 16'h6969;
    SB_LUT4 n71113_bdd_4_lut (.I0(n71113), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n71116));
    defparam n71113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1687 (.I0(\data_in_frame[7][1] ), .I1(\data_in_frame[4] [7]), 
            .I2(n59174), .I3(n26750), .O(n59276));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1687.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1688 (.I0(\data_in_frame[18] [3]), .I1(n60988), 
            .I2(\data_in_frame[20][4] ), .I3(\data_in_frame[20][3] ), .O(n59338));
    defparam i2_3_lut_4_lut_adj_1688.LUT_INIT = 16'h6996;
    SB_LUT4 i16118_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30525));
    defparam i16118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16115_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30522));
    defparam i16115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_810_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5507));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13] [4]), .I3(GND_net), .O(n59510));
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1690 (.I0(n26281), .I1(\data_in_frame[10] [7]), 
            .I2(n26365), .I3(\data_in_frame[11] [1]), .O(n59638));
    defparam i3_3_lut_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 i16112_3_lut_4_lut (.I0(n8_adj_12), .I1(n59083), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30519));
    defparam i16112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n69097), .I2(n66958), .I3(byte_transmit_counter_c[4]), 
            .O(n71107));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1691 (.I0(n54440), .I1(n59504), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16]_c [5]), .O(n59443));
    defparam i1_2_lut_4_lut_adj_1691.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1692 (.I0(n54440), .I1(n59504), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16]_c [6]), .O(n59110));
    defparam i1_2_lut_4_lut_adj_1692.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n70813_bdd_4_lut (.I0(n70813), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n70816));
    defparam n70813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1693 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(n59097), .I3(GND_net), .O(Kp_23__N_1209));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1693.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1694 (.I0(\FRAME_MATCHER.i_31__N_2642 ), .I1(Kp_23__N_1877), 
            .I2(\FRAME_MATCHER.i_31__N_2641 ), .I3(GND_net), .O(n6_adj_5602));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_adj_1694.LUT_INIT = 16'hfefe;
    SB_LUT4 i14854_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2637 ), 
            .I2(GND_net), .I3(GND_net), .O(n29261));   // verilog/coms.v(130[12] 305[6])
    defparam i14854_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_810_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n71107_bdd_4_lut (.I0(n71107), .I1(n14_adj_5461), .I2(n7_adj_5803), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n71107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1695 (.I0(\data_in_frame[8]_c [1]), .I1(n53944), 
            .I2(n59761), .I3(n26316), .O(n59762));
    defparam i2_3_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1696 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[5] [7]), .O(n6_adj_5594));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1697 (.I0(\data_in_frame[20][2] ), .I1(n26395), 
            .I2(n26376), .I3(\data_in_frame[13] [5]), .O(n6_adj_5592));
    defparam i1_2_lut_4_lut_adj_1697.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1698 (.I0(\data_in_frame[17][7] ), .I1(\data_in_frame[17][6] ), 
            .I2(n61866), .I3(GND_net), .O(n59647));
    defparam i1_2_lut_3_lut_adj_1698.LUT_INIT = 16'h6969;
    SB_LUT4 select_810_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1699 (.I0(\data_out_frame[23] [4]), .I1(n54750), 
            .I2(\data_out_frame[23] [6]), .I3(\data_out_frame[25] [7]), 
            .O(n4_adj_5552));
    defparam i1_2_lut_4_lut_adj_1699.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5729));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i43868_3_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i [0]), .I2(n43937), 
            .I3(n59093), .O(n59994));
    defparam i43868_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_adj_1700 (.I0(\data_in_frame[12] [4]), .I1(n26902), 
            .I2(n54440), .I3(GND_net), .O(n59377));
    defparam i1_2_lut_3_lut_adj_1700.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5728));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1701 (.I0(\data_in_frame[5] [6]), .I1(n26333), 
            .I2(\data_in_frame[8]_c [1]), .I3(\data_in_frame[8]_c [2]), 
            .O(n6_adj_5546));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1701.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5727));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14834_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n29241));   // verilog/coms.v(130[12] 305[6])
    defparam i14834_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54666 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64562), .I2(n64563), .I3(\byte_transmit_counter[2] ), 
            .O(n70807));
    defparam byte_transmit_counter_1__bdd_4_lut_54666.LUT_INIT = 16'he4aa;
    SB_LUT4 select_810_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5726));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5725));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1702 (.I0(n26376), .I1(\data_in_frame[11] [2]), 
            .I2(n26719), .I3(GND_net), .O(n6_adj_5544));
    defparam i1_2_lut_3_lut_adj_1702.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1703 (.I0(n26598), .I1(n54954), .I2(n59285), 
            .I3(GND_net), .O(n38));
    defparam i1_2_lut_3_lut_adj_1703.LUT_INIT = 16'h6969;
    SB_LUT4 select_810_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5724));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23_4_lut_4_lut (.I0(n55007), .I1(\data_in_frame[17]_c [0]), 
            .I2(n59726), .I3(GND_net), .O(n60_adj_5542));
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 select_810_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5723));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1704 (.I0(n26598), .I1(n54954), .I2(\data_in_frame[16]_c [3]), 
            .I3(GND_net), .O(n59517));
    defparam i1_2_lut_3_lut_adj_1704.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1705 (.I0(\data_out_frame[21] [5]), .I1(n54996), 
            .I2(n59141), .I3(\data_out_frame[21] [7]), .O(n59746));
    defparam i2_3_lut_4_lut_adj_1705.LUT_INIT = 16'h9669;
    SB_LUT4 select_810_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5722));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5721));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1706 (.I0(\data_in_frame[16]_c [5]), .I1(\data_in_frame[16]_c [6]), 
            .I2(\data_in_frame[16]_c [4]), .I3(GND_net), .O(n6_adj_5508));
    defparam i1_2_lut_3_lut_adj_1706.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5720));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[23] [3]), 
            .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5719));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'ha088;
    SB_LUT4 n70807_bdd_4_lut (.I0(n70807), .I1(n64554), .I2(n64553), .I3(\byte_transmit_counter[2] ), 
            .O(n70810));
    defparam n70807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_810_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5718));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5715));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1708 (.I0(n26395), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n6_adj_5485));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 select_810_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5714));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1709 (.I0(n26447), .I1(n59239), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[15] [1]), .O(n59678));
    defparam i1_2_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5713));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1710 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n55066), .I3(GND_net), .O(n54914));
    defparam i1_2_lut_3_lut_adj_1710.LUT_INIT = 16'h6969;
    SB_LUT4 select_810_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5712));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1711 (.I0(\data_in_frame[15] [5]), .I1(n26389), 
            .I2(n55066), .I3(n61866), .O(n26197));
    defparam i2_3_lut_4_lut_adj_1711.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5711));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(n55007), .I1(n54600), .I2(n26568), 
            .I3(GND_net), .O(n27228));
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1713 (.I0(n26568), .I1(n54732), .I2(\data_in_frame[19] [4]), 
            .I3(n54971), .O(n59488));
    defparam i1_2_lut_4_lut_adj_1713.LUT_INIT = 16'h6996;
    SB_LUT4 select_810_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5710));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1714 (.I0(n60966), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [3]), .I3(n59423), .O(n61159));
    defparam i2_3_lut_4_lut_adj_1714.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1715 (.I0(n60966), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[23] [2]), .I3(n59464), .O(n61145));
    defparam i2_3_lut_4_lut_adj_1715.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1084_i2_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n5169[1]));
    defparam mux_1084_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i3_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n5169[2]));
    defparam mux_1084_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i4_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n5169[3]));
    defparam mux_1084_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i5_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n5169[4]));
    defparam mux_1084_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i6_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n5169[5]));
    defparam mux_1084_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5709));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1084_i7_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n5169[6]));
    defparam mux_1084_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_4_lut_adj_1716 (.I0(\data_in_frame[15] [5]), .I1(n54914), 
            .I2(n61866), .I3(\data_in_frame[17][6] ), .O(n59437));
    defparam i1_2_lut_4_lut_adj_1716.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1084_i8_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n5169[7]));
    defparam mux_1084_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54859 (.I0(byte_transmit_counter_c[3]), 
            .I1(n70906), .I2(n67132), .I3(byte_transmit_counter_c[4]), 
            .O(n71101));
    defparam byte_transmit_counter_3__bdd_4_lut_54859.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1084_i9_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n5169[8]));
    defparam mux_1084_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i10_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n5169[9]));
    defparam mux_1084_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5706));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1084_i11_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n5169[10]));
    defparam mux_1084_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5705));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[22] [4]), 
            .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5704));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1084_i12_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n5169[11]));
    defparam mux_1084_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5703));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[22] [2]), 
            .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5702));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1084_i13_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n5169[12]));
    defparam mux_1084_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i14_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n5169[13]));
    defparam mux_1084_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 n71101_bdd_4_lut (.I0(n71101), .I1(n70786), .I2(n70876), .I3(byte_transmit_counter_c[4]), 
            .O(tx_data[4]));
    defparam n71101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1084_i15_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n5169[14]));
    defparam mux_1084_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54617 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n70795));
    defparam byte_transmit_counter_0__bdd_4_lut_54617.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1084_i16_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n5169[15]));
    defparam mux_1084_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i24124_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[1]_c [0]), 
            .I3(\data_in_frame[17]_c [0]), .O(n5169[16]));
    defparam i24124_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i18_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1][1] ), .I3(\data_in_frame[17] [1]), .O(n5169[17]));
    defparam mux_1084_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5701));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54854 (.I0(byte_transmit_counter_c[3]), 
            .I1(n69091), .I2(n66957), .I3(byte_transmit_counter_c[4]), 
            .O(n71095));
    defparam byte_transmit_counter_3__bdd_4_lut_54854.LUT_INIT = 16'he4aa;
    SB_LUT4 select_810_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2638 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5699));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_3_lut (.I0(LED_N_3537), .I1(\FRAME_MATCHER.i_31__N_2642 ), 
            .I2(reset), .I3(GND_net), .O(n23164));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mux_1084_i19_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n5169[18]));
    defparam mux_1084_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i20_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n5169[19]));
    defparam mux_1084_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5698));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_810_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5696));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1084_i21_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n5169[20]));
    defparam mux_1084_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i22_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n5169[21]));
    defparam mux_1084_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i23_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17][6] ), .O(n5169[22]));
    defparam mux_1084_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1084_i24_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17][7] ), .O(n5169[23]));
    defparam mux_1084_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_810_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5695));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23021_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[16]_c [0]), 
            .I3(deadband[0]), .O(n29998));
    defparam i23021_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15595_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n30002));
    defparam i15595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15599_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n30006));
    defparam i15599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15600_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n30007));
    defparam i15600_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70795_bdd_4_lut (.I0(n70795), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n70798));
    defparam n70795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54612 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64406), .I2(n64407), .I3(\byte_transmit_counter[2] ), 
            .O(n70789));
    defparam byte_transmit_counter_1__bdd_4_lut_54612.LUT_INIT = 16'he4aa;
    SB_LUT4 i15604_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n30011));
    defparam i15604_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70789_bdd_4_lut (.I0(n70789), .I1(n64524), .I2(n64523), .I3(\byte_transmit_counter[2] ), 
            .O(n70792));
    defparam n70789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15669_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8][7] ), 
            .I3(PWMLimit[23]), .O(n30076));
    defparam i15669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54598 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64511), .I2(n64512), .I3(\byte_transmit_counter[2] ), 
            .O(n70783));
    defparam byte_transmit_counter_1__bdd_4_lut_54598.LUT_INIT = 16'he4aa;
    SB_LUT4 i15670_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n30077));
    defparam i15670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70783_bdd_4_lut (.I0(n70783), .I1(n64506), .I2(n64505), .I3(\byte_transmit_counter[2] ), 
            .O(n70786));
    defparam n70783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_810_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5694));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15671_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8][5] ), 
            .I3(PWMLimit[21]), .O(n30078));
    defparam i15671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15672_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8][4] ), 
            .I3(PWMLimit[20]), .O(n30079));
    defparam i15672_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15673_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8][3] ), 
            .I3(PWMLimit[19]), .O(n30080));
    defparam i15673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23599_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8]_c [2]), 
            .I3(PWMLimit[18]), .O(n30081));
    defparam i23599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15675_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8]_c [1]), 
            .I3(PWMLimit[17]), .O(n30082));
    defparam i15675_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54603 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n70777));
    defparam byte_transmit_counter_0__bdd_4_lut_54603.LUT_INIT = 16'he4aa;
    SB_LUT4 i15676_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[8]_c [0]), 
            .I3(PWMLimit[16]), .O(n30083));
    defparam i15676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70777_bdd_4_lut (.I0(n70777), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n70780));
    defparam n70777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_810_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5693));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15677_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n30084));
    defparam i15677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54593 (.I0(\byte_transmit_counter[1] ), 
            .I1(n64559), .I2(n64560), .I3(\byte_transmit_counter[2] ), 
            .O(n70771));
    defparam byte_transmit_counter_1__bdd_4_lut_54593.LUT_INIT = 16'he4aa;
    SB_LUT4 i15678_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n30085));
    defparam i15678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70771_bdd_4_lut (.I0(n70771), .I1(n64569), .I2(n64568), .I3(\byte_transmit_counter[2] ), 
            .O(n70774));
    defparam n70771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15679_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n30086));
    defparam i15679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_810_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5692));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54588 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n70765));
    defparam byte_transmit_counter_0__bdd_4_lut_54588.LUT_INIT = 16'he4aa;
    SB_LUT4 n70765_bdd_4_lut (.I0(n70765), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n70768));
    defparam n70765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1719 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(n25998), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5419));
    defparam i1_3_lut_4_lut_adj_1719.LUT_INIT = 16'hfefc;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54579 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n70759));
    defparam byte_transmit_counter_0__bdd_4_lut_54579.LUT_INIT = 16'he4aa;
    SB_LUT4 n70759_bdd_4_lut (.I0(n70759), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n70762));
    defparam n70759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15680_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n30087));
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(\FRAME_MATCHER.i_31__N_2638 ), .I1(\data_out_frame[21] [1]), 
            .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5691));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54574 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70753));
    defparam byte_transmit_counter_0__bdd_4_lut_54574.LUT_INIT = 16'he4aa;
    SB_LUT4 n70753_bdd_4_lut (.I0(n70753), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70756));
    defparam n70753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_810_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5690));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54569 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n70747));
    defparam byte_transmit_counter_0__bdd_4_lut_54569.LUT_INIT = 16'he4aa;
    SB_LUT4 i15681_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n30088));
    defparam i15681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15682_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n30089));
    defparam i15682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15694_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n30101));
    defparam i15694_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15698_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n30105));
    defparam i15698_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70747_bdd_4_lut (.I0(n70747), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n70750));
    defparam n70747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_810_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2638 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2741 [3]), 
            .O(n2_adj_5688));   // verilog/coms.v(148[4] 304[11])
    defparam select_810_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54564 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n70741));
    defparam byte_transmit_counter_0__bdd_4_lut_54564.LUT_INIT = 16'he4aa;
    SB_LUT4 i15699_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n30106));
    defparam i15699_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71095_bdd_4_lut (.I0(n71095), .I1(n70810), .I2(n7_adj_5802), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n71095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15700_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n30107));
    defparam i15700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15701_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n30108));
    defparam i15701_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n70741_bdd_4_lut (.I0(n70741), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n70744));
    defparam n70741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15705_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n30112));
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15708_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n30115));
    defparam i15708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15712_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n30119));
    defparam i15712_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i50990_2_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67006));
    defparam i50990_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i23027_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n30120));
    defparam i23027_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51109_2_lut (.I0(\data_out_frame[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67007));
    defparam i51109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5687));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_adj_5686));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14101_2_lut (.I0(\byte_transmit_counter[1] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n28507));   // verilog/coms.v(109[34:55])
    defparam i14101_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15724_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n30131));
    defparam i15724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15725_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n30132));
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15726_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n30133));
    defparam i15726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15727_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n30134));
    defparam i15727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i29459_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n30135));
    defparam i29459_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15729_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n30136));
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54559 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n70729));
    defparam byte_transmit_counter_0__bdd_4_lut_54559.LUT_INIT = 16'he4aa;
    SB_LUT4 n70729_bdd_4_lut (.I0(n70729), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n70732));
    defparam n70729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15730_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n30137));
    defparam i15730_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15731_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n30138));
    defparam i15731_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54550 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n70723));
    defparam byte_transmit_counter_0__bdd_4_lut_54550.LUT_INIT = 16'he4aa;
    SB_LUT4 n70723_bdd_4_lut (.I0(n70723), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n70726));
    defparam n70723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54545 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n70717));
    defparam byte_transmit_counter_0__bdd_4_lut_54545.LUT_INIT = 16'he4aa;
    SB_LUT4 n70717_bdd_4_lut (.I0(n70717), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n70720));
    defparam n70717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54540 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n70711));
    defparam byte_transmit_counter_0__bdd_4_lut_54540.LUT_INIT = 16'he4aa;
    SB_LUT4 n70711_bdd_4_lut (.I0(n70711), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n70714));
    defparam n70711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15732_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n30139));
    defparam i15732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1721 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59127));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1721.LUT_INIT = 16'h6666;
    SB_LUT4 i23790_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n30140));
    defparam i23790_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15734_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n30141));
    defparam i15734_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1722 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n5));
    defparam i1_3_lut_adj_1722.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54849 (.I0(byte_transmit_counter_c[3]), 
            .I1(n69089), .I2(n67091), .I3(byte_transmit_counter_c[4]), 
            .O(n71089));
    defparam byte_transmit_counter_3__bdd_4_lut_54849.LUT_INIT = 16'he4aa;
    SB_LUT4 i15735_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n30142));
    defparam i15735_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15736_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n30143));
    defparam i15736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1723 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n26786));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1723.LUT_INIT = 16'h9696;
    SB_LUT4 i15737_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n30144));
    defparam i15737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_4_lut_adj_1724 (.I0(\data_in_frame[0] [4]), .I1(ID[6]), .I2(ID[4]), 
            .I3(\data_in_frame[0] [6]), .O(n6_adj_5811));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1724.LUT_INIT = 16'h7bde;
    SB_LUT4 n71089_bdd_4_lut (.I0(n71089), .I1(n14_adj_5453), .I2(n7_adj_5801), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n71089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[0]), .I3(ID[2]), .O(n5_adj_5812));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n5_adj_5812), .I1(\data_in_frame[0] [3]), 
            .I2(n6_adj_5811), .I3(ID[3]), .O(n6_adj_5813));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfbfe;
    SB_LUT4 i15738_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n30145));
    defparam i15738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15739_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n30146));
    defparam i15739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15740_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n30147));
    defparam i15740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_4_lut_adj_1727 (.I0(ID[1]), .I1(\data_in_frame[0] [5]), .I2(\data_in_frame[0] [1]), 
            .I3(ID[5]), .O(n7_adj_5814));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1727.LUT_INIT = 16'h7bde;
    SB_LUT4 i51108_2_lut (.I0(n70858), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66942));
    defparam i51108_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15741_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n30148));
    defparam i15741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1728 (.I0(n7_adj_5814), .I1(\data_in_frame[0] [7]), 
            .I2(n6_adj_5813), .I3(ID[7]), .O(n53451));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1728.LUT_INIT = 16'hfbfe;
    SB_LUT4 i15742_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n30149));
    defparam i15742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15743_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n30150));
    defparam i15743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1729 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n59144));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1730 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n59135));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1730.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1731 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59410));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1731.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1732 (.I0(\data_in_frame[0] [7]), .I1(n59410), 
            .I2(n59135), .I3(n59121), .O(Kp_23__N_877));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 i52814_3_lut (.I0(n70726), .I1(n70798), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n68989));
    defparam i52814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54844 (.I0(byte_transmit_counter_c[3]), 
            .I1(n70834), .I2(n67089), .I3(\byte_transmit_counter[1] ), 
            .O(n71083));
    defparam byte_transmit_counter_3__bdd_4_lut_54844.LUT_INIT = 16'he4aa;
    SB_LUT4 i15744_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n30151));
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1733 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n59121));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1733.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1734 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_877), 
            .I2(GND_net), .I3(GND_net), .O(n59245));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1734.LUT_INIT = 16'h6666;
    SB_LUT4 equal_2043_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // verilog/coms.v(169[9:87])
    defparam equal_2043_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1735 (.I0(n26231), .I1(Kp_23__N_877), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22));
    defparam i5_3_lut_adj_1735.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1736 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [6]), .O(n27_c));
    defparam i10_4_lut_adj_1736.LUT_INIT = 16'h8000;
    SB_LUT4 i15745_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n30152));
    defparam i15745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15746_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n30153));
    defparam i15746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15747_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [7]), 
            .I3(\Kp[7] ), .O(n30154));
    defparam i15747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15748_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [6]), 
            .I3(\Kp[6] ), .O(n30155));
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15749_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [5]), 
            .I3(\Kp[5] ), .O(n30156));
    defparam i15749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15750_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n30157));
    defparam i15750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15751_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [3]), 
            .I3(\Kp[3] ), .O(n30158));
    defparam i15751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15752_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [2]), 
            .I3(\Kp[2] ), .O(n30159));
    defparam i15752_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15753_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n30160));
    defparam i15753_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15754_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n30161));
    defparam i15754_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15755_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n30162));
    defparam i15755_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15756_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n30163));
    defparam i15756_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71083_bdd_4_lut (.I0(n71083), .I1(n67090), .I2(n70840), .I3(\byte_transmit_counter[1] ), 
            .O(n71086));
    defparam n71083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15757_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n30164));
    defparam i15757_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i47895_3_lut_4_lut (.I0(\data_in_frame[2] [3]), .I1(n59410), 
            .I2(\data_in_frame[2] [7]), .I3(n59135), .O(n64058));
    defparam i47895_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51146_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2636 ), 
            .I2(GND_net), .I3(GND_net), .O(n66924));   // verilog/coms.v(158[12:15])
    defparam i51146_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15758_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n30165));
    defparam i15758_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i22670_3_lut_4_lut (.I0(Kp_23__N_741), .I1(Kp_23__N_1877), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n30166));
    defparam i22670_3_lut_4_lut.LUT_INIT = 16'hf780;
    uart_tx tx (.\o_Rx_DV_N_3617[24] (\o_Rx_DV_N_3617[24] ), .r_SM_Main({r_SM_Main}), 
            .n27(n27), .n62584(n62584), .n28320(n28320), .clk16MHz(clk16MHz), 
            .n60079(n60079), .n1(n1), .tx_o(tx_o), .tx_data({tx_data}), 
            .GND_net(GND_net), .r_Clock_Count({r_Clock_Count}), .VCC_net(VCC_net), 
            .n30034(n30034), .tx_active(tx_active), .n71131(n71131), .n30847(n30847), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .\r_SM_Main_2__N_3674[0] (r_SM_Main_2__N_3674[0]), 
            .n62490(n62490), .\r_SM_Main_2__N_3665[1] (r_SM_Main_2__N_3665[1]), 
            .n60937(n60937), .n60609(n60609), .n6(n6), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .\o_Rx_DV_N_3617[12] (\o_Rx_DV_N_3617[12] ), 
            .n5254(n5254), .\o_Rx_DV_N_3617[8] (\o_Rx_DV_N_3617[8] ), .r_Rx_Data(r_Rx_Data), 
            .\o_Rx_DV_N_3617[24] (\o_Rx_DV_N_3617[24] ), .n29(n29), .n23(n23), 
            .\r_SM_Main[1] (\r_SM_Main[1]_adj_14 ), .n27(n27), .VCC_net(VCC_net), 
            .baudrate({baudrate}), .n28324(n28324), .clk16MHz(clk16MHz), 
            .n60053(n60053), .\r_SM_Main[2] (\r_SM_Main[2]_adj_15 ), .RX_N_2(RX_N_2), 
            .r_Clock_Count({r_Clock_Count_adj_25}), .n30256(n30256), .rx_data({rx_data}), 
            .n30255(n30255), .n30254(n30254), .n30253(n30253), .n30252(n30252), 
            .n25975(n25975), .\o_Rx_DV_N_3617[7] (\o_Rx_DV_N_3617[7] ), 
            .\o_Rx_DV_N_3617[6] (\o_Rx_DV_N_3617[6] ), .\o_Rx_DV_N_3617[5] (\o_Rx_DV_N_3617[5] ), 
            .\o_Rx_DV_N_3617[4] (\o_Rx_DV_N_3617[4] ), .\o_Rx_DV_N_3617[3] (\o_Rx_DV_N_3617[3] ), 
            .\o_Rx_DV_N_3617[2] (\o_Rx_DV_N_3617[2] ), .\o_Rx_DV_N_3617[1] (\o_Rx_DV_N_3617[1] ), 
            .\o_Rx_DV_N_3617[0] (\o_Rx_DV_N_3617[0] ), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_24 ), 
            .n62864(n62864), .n29921(n29921), .n59011(n59011), .n62764(n62764), 
            .n62780(n62780), .n62748(n62748), .n62828(n62828), .n62812(n62812), 
            .n30854(n30854), .n55126(n55126), .rx_data_ready(rx_data_ready), 
            .n30850(n30850), .n5257(n5257), .n60937(n60937), .n62490(n62490), 
            .n29791(n29791), .\r_SM_Main_2__N_3665[1] (r_SM_Main_2__N_3665[1]), 
            .n28127(n28127), .n62796(n62796), .n62846(n62846), .\r_SM_Main[0] (r_SM_Main[0]), 
            .n60609(n60609)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (\o_Rx_DV_N_3617[24] , r_SM_Main, n27, n62584, n28320, 
            clk16MHz, n60079, n1, tx_o, tx_data, GND_net, r_Clock_Count, 
            VCC_net, n30034, tx_active, n71131, n30847, \r_Bit_Index[0] , 
            \r_SM_Main_2__N_3674[0] , n62490, \r_SM_Main_2__N_3665[1] , 
            n60937, n60609, n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input \o_Rx_DV_N_3617[24] ;
    output [2:0]r_SM_Main;
    input n27;
    input n62584;
    output n28320;
    input clk16MHz;
    output n60079;
    output n1;
    output tx_o;
    input [7:0]tx_data;
    input GND_net;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n30034;
    output tx_active;
    input n71131;
    input n30847;
    output \r_Bit_Index[0] ;
    input \r_SM_Main_2__N_3674[0] ;
    input n62490;
    input \r_SM_Main_2__N_3665[1] ;
    output n60937;
    input n60609;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n3;
    wire [2:0]n460;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n3_adj_5400, n25486;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n22796;
    wire [8:0]n41;
    
    wire n52823, n52822, n52821, n52820, n52819, n52818, n52817, 
        n52816, n29506, n22795, n70738, n71074, o_Tx_Serial_N_3727, 
        n59997, n71071, n70735;
    
    SB_LUT4 i8916_4_lut (.I0(\o_Rx_DV_N_3617[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n62584), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i8916_4_lut.LUT_INIT = 16'hc9cc;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28320), 
            .D(n460[1]), .R(n60079));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28320), 
            .D(n460[2]), .R(n60079));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3_adj_5400));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n22796), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_2064_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n52823), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2064_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52822), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_9 (.CI(n52822), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n52823));
    SB_LUT4 r_Clock_Count_2064_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52821), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_8 (.CI(n52821), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52822));
    SB_LUT4 r_Clock_Count_2064_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52820), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_7 (.CI(n52820), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52821));
    SB_LUT4 r_Clock_Count_2064_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52819), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_6 (.CI(n52819), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52820));
    SB_LUT4 r_Clock_Count_2064_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52818), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_5 (.CI(n52818), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52819));
    SB_LUT4 r_Clock_Count_2064_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52817), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_4 (.CI(n52817), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52818));
    SB_LUT4 r_Clock_Count_2064_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52816), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_3 (.CI(n52816), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52817));
    SB_LUT4 r_Clock_Count_2064_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2064_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2064_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52816));
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n30034));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n71131));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_2064__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2064__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n29506));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30847));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25486), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i8667_4_lut (.I0(\r_SM_Main_2__N_3674[0] ), .I1(n62490), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n22795));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i8667_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i8668_3_lut (.I0(n22795), .I1(\r_SM_Main_2__N_3665[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n22796));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i8668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3070895_i1_3_lut (.I0(n70738), .I1(n71074), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3727));
    defparam i3070895_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3727), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_5400));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i2257_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2257_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i43871_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n59997));
    defparam i43871_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n60937));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2250_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2250_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54514_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_3665[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n28320));
    defparam i54514_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i54313_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3665[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n29506));
    defparam i54313_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n60609), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3674[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i54402_4_lut_4_lut (.I0(\r_SM_Main_2__N_3665[1] ), .I1(r_SM_Main[1]), 
            .I2(n59997), .I3(n60937), .O(n60079));
    defparam i54402_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3674[0] ), .O(n25486));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n71071));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71071_bdd_4_lut (.I0(n71071), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n71074));
    defparam n71071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_54829 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n70735));
    defparam r_Bit_Index_0__bdd_4_lut_54829.LUT_INIT = 16'he4aa;
    SB_LUT4 n70735_bdd_4_lut (.I0(n70735), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n70738));
    defparam n70735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, \o_Rx_DV_N_3617[12] , n5254, \o_Rx_DV_N_3617[8] , 
            r_Rx_Data, \o_Rx_DV_N_3617[24] , n29, n23, \r_SM_Main[1] , 
            n27, VCC_net, baudrate, n28324, clk16MHz, n60053, \r_SM_Main[2] , 
            RX_N_2, r_Clock_Count, n30256, rx_data, n30255, n30254, 
            n30253, n30252, n25975, \o_Rx_DV_N_3617[7] , \o_Rx_DV_N_3617[6] , 
            \o_Rx_DV_N_3617[5] , \o_Rx_DV_N_3617[4] , \o_Rx_DV_N_3617[3] , 
            \o_Rx_DV_N_3617[2] , \o_Rx_DV_N_3617[1] , \o_Rx_DV_N_3617[0] , 
            \r_Bit_Index[0] , n62864, n29921, n59011, n62764, n62780, 
            n62748, n62828, n62812, n30854, n55126, rx_data_ready, 
            n30850, n5257, n60937, n62490, n29791, \r_SM_Main_2__N_3665[1] , 
            n28127, n62796, n62846, \r_SM_Main[0] , n60609) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \o_Rx_DV_N_3617[12] ;
    input n5254;
    output \o_Rx_DV_N_3617[8] ;
    output r_Rx_Data;
    output \o_Rx_DV_N_3617[24] ;
    output n29;
    output n23;
    output \r_SM_Main[1] ;
    output n27;
    input VCC_net;
    input [31:0]baudrate;
    output n28324;
    input clk16MHz;
    output n60053;
    output \r_SM_Main[2] ;
    input RX_N_2;
    output [7:0]r_Clock_Count;
    input n30256;
    output [7:0]rx_data;
    input n30255;
    input n30254;
    input n30253;
    input n30252;
    output n25975;
    output \o_Rx_DV_N_3617[7] ;
    output \o_Rx_DV_N_3617[6] ;
    output \o_Rx_DV_N_3617[5] ;
    output \o_Rx_DV_N_3617[4] ;
    output \o_Rx_DV_N_3617[3] ;
    output \o_Rx_DV_N_3617[2] ;
    output \o_Rx_DV_N_3617[1] ;
    output \o_Rx_DV_N_3617[0] ;
    output \r_Bit_Index[0] ;
    output n62864;
    input n29921;
    input n59011;
    output n62764;
    output n62780;
    output n62748;
    output n62828;
    output n62812;
    input n30854;
    input n55126;
    output rx_data_ready;
    input n30850;
    input n5257;
    input n60937;
    output n62490;
    input n29791;
    output \r_SM_Main_2__N_3665[1] ;
    output n28127;
    output n62796;
    output n62846;
    input \r_SM_Main[0] ;
    output n60609;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2955;
    wire [23:0]n8825;
    wire [23:0]n294;
    
    wire n3063;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n67016, n58782, n67022, n64264, n60197, n67013, n2939, 
        n3047, n2941, n3049, n2940, n3048, n52438, n1977, n858, 
        n52439, n67019;
    wire [23:0]n8773;
    
    wire n2730, n52524, n3;
    wire [23:0]n8617;
    
    wire n538, n2944, n3052, n35, n2942, n3050, n39, n2945, 
        n3053, n33, n2943, n3051, n37, n52525, n2949, n3057, 
        n2950, n3058, n63984, n60171, n23_adj_5124, n25, n2947, 
        n3055, n2948, n3056, n27_adj_5125, n29_adj_5126, n2951, 
        n3059, n21, n2952, n3060, n2946, n3054, n2954, n3062, 
        n2953, n3061, n15, n17, n19, n31, n2956, n3064, n2957, 
        n3065, n11, n13, n67191, n68109, n68832, n68830, n67193, 
        n3066, n8, n69380, n69381, n16, n34, n67187, n14, n67182, 
        n69736, n69295, n10, n69382, n69383, n67203, n68097, n12, 
        n20, n69293, n69139, n69867, n69298, n69889, n69890, n69884, 
        n69300, n2828;
    wire [23:0]n8799;
    
    wire n2843, n2829, n2832, n37_adj_5127, n2830, n41, n2833, 
        n35_adj_5128, n2831, n39_adj_5129, n2835, n2836, n29_adj_5130, 
        n31_adj_5131, n2837, n2838, n2839, n23_adj_5132, n25_adj_5133, 
        n27_adj_5134, n2834;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n2840, n2842, n2841, n17_adj_5135, n19_adj_5136, n21_adj_5137, 
        n33_adj_5138, n2844, n2845, n13_adj_5139, n15_adj_5140, n67248, 
        n68151, n68852, n68850, n67250, n10_adj_5141, n69386, n69387, 
        n18, n36, n67243, n16_adj_5142, n67238, n69734, n69289, 
        n14_adj_5143, n22, n12_adj_5144, n67258, n69732, n69733, 
        n69592, n69149, n69865, n69558, n69893, n69894, n69888, 
        n2827, n2938, n3046, n3186;
    wire [23:0]n8851;
    
    wire n3151, n2713, n2714, n2719, n2717, n39_adj_5145, n2718, 
        n37_adj_5146, n2715, n43, n2716, n41_adj_5147, n2720, n2721, 
        n31_adj_5148, n33_adj_5149, n2722, n2724, n2723, n25_adj_5150, 
        n27_adj_5151, n29_adj_5152, n2725, n2726, n2729, n2728, 
        n15_adj_5153, n17_adj_5154, n2727, n19_adj_5155, n21_adj_5156, 
        n23_adj_5157, n35_adj_5158, n67310, n68241, n68864, n68862, 
        n64272, n60147, n67313, n12_adj_5159, n69392, n20_adj_5160, 
        n38, n69393, n67305, n18_adj_5161, n67302, n69390, n69281;
    wire [23:0]n8591;
    
    wire n1831, n2144, n52437, n16_adj_5162, n24, n14_adj_5163, 
        n67332, n69730, n69731, n69594, n69183, n69784, n69556, 
        n69859, n69860, n1832, n2013, n52436, n2596;
    wire [23:0]n8747;
    
    wire n2601, n2597, n45, n2599, n41_adj_5164, n2600, n39_adj_5165, 
        n2598, n43_adj_5166, n2604, n2606, n2605, n27_adj_5167, 
        n29_adj_5168, n31_adj_5169, n2602, n3_adj_5170, n2603, n33_adj_5171, 
        n35_adj_5172, r_Rx_Data_R, n2610, n2611, n2612, n17_adj_5173, 
        n19_adj_5174, n2607, n2608, n2609, n62394, n60155, n21_adj_5175, 
        n23_adj_5176, n2867, n52523, n1833, n1879, n52435, n25_adj_5177, 
        n37_adj_5178, n67352, n68275, n68878, n2754, n52522, n68876, 
        n67354, n14_adj_5179, n69396, n69397, n22_adj_5180, n40, 
        n67348, n20_adj_5181, n67345, n68941, n69277, n18_adj_5182, 
        n26, n2638, n52521, n16_adj_5183, n67367, n69728, n69729, 
        n1834, n1742, n52434, n69596, n2519, n52520, n69195, n69552, 
        n1835, n1602, n52433, n69551, n69554, n2397, n52519, n1836, 
        n1459, n52432, n2272, n52518, n2106, n31_adj_5184, n2107, 
        n29_adj_5185, n2105, n33_adj_5186, n2104, n35_adj_5187, n2102, 
        n39_adj_5188, n2103, n37_adj_5189, n2101, n41_adj_5190, n2236, 
        n29_adj_5191, n2235, n31_adj_5192, n2237, n27_adj_5193, n2233, 
        n35_adj_5194, n52517, n2238, n25_adj_5195, n52516, n1837, 
        n1460, n52431, n2232, n37_adj_5196, n2231, n39_adj_5197, 
        n2230, n41_adj_5198, n2234, n33_adj_5199, n2363, n27_adj_5200, 
        n2362, n29_adj_5201, n2364, n25_adj_5202, n52515, n2360, 
        n33_adj_5203, n2365, n23_adj_5204, n2359, n35_adj_5205, n1838, 
        n1011, n52430, n52514, n2358, n37_adj_5206, n2357, n39_adj_5207, 
        n2361, n31_adj_5208, n2356, n41_adj_5209, n1974, n31_adj_5210, 
        n1975, n29_adj_5211, n1973, n33_adj_5212, n1972, n35_adj_5213, 
        n1970, n39_adj_5214, n1971, n37_adj_5215, n1969, n41_adj_5216, 
        n2487, n25_adj_5217, n2486, n27_adj_5218, n2485, n29_adj_5219, 
        n2488, n23_adj_5220, n2484, n31_adj_5221, n2489, n21_adj_5222, 
        n2483, n33_adj_5223, n52513, n2482, n35_adj_5224, n2481, 
        n37_adj_5225, n2479, n41_adj_5226, n2478, n43_adj_5227, n2480, 
        n39_adj_5228, n1839, n856, n52429, n52512, n2477, n45_adj_5229, 
        n1697, n39_adj_5230, n1696, n41_adj_5231, n1556, n39_adj_5232, 
        n1555, n41_adj_5233, n1557, n37_adj_5234, n64187, n1840, 
        n698, n52428, n44073, n52511, n44071, n804, n21434, n21436, 
        n52510, n1411, n41_adj_5235, n1410, n43_adj_5236, n1412, 
        n39_adj_5237;
    wire [7:0]n1;
    
    wire n52815, n52509, n52814, n71130, n52508, n1841, n52427, 
        n51522, n26081, n60143, n51521, n62352, n64302, n51520, 
        n62432, n52813, n62384, n60180, n52507, n52812, n52811;
    wire [23:0]n8565;
    
    wire n1693, n52426, n52810, n1694, n52425, n62392, n60159, 
        n52809, n1695, n52424, n51519;
    wire [24:0]o_Rx_DV_N_3617;
    wire [23:0]n8721;
    
    wire n2476, n52506, n52423, n52505, n51518, n62430, n51517, 
        n62428, n52422, n51516, n52504, n51515, n62426, n51514, 
        n62424, n51513, n62350, n51512, n62422, n1698, n52421, 
        n51511, n52503, n52502, n1699, n52420, n51510, n51509, 
        n51508, n52501, n51507, n51506, n51505, n1700, n52419, 
        n51504, n51503, n1413, n1414, n67626, n52500, n1701, n52418, 
        n51502;
    wire [23:0]n8877;
    
    wire n52624, n3152, n3082, n52623, n3153, n3188, n52622, n52499, 
        n1702, n26055, n60151, n51501, n36_adj_5244, n51500, n51499, 
        n3154, n3084, n52621, n52498;
    wire [23:0]n8539;
    
    wire n1552, n52417, n61327, n3155, n2977, n52620, n1553, n52416, 
        n52497, n3156, n52619, n52496, n3157, n52618, n3158, n52617, 
        n1114, n40_adj_5245, n3159, n52616, n1115, n67641, n1554, 
        n52415, n52495, n52414, n3160, n52615, n3161, n52614, 
        n3162, n52613, n1558, n1559, n67614, n3163, n52612, n3164, 
        n52611, n52494, n34_adj_5246, n67603, n3165, n52610, n34_adj_5247, 
        n4, n62852, n62858, n63858, n62370, n62368, n63810, n26049, 
        n1265, n38_adj_5248, n62880, n62884, n1266, n67634, n62886, 
        n3166, n52609, n64062, n64064, n52413, n62882, n64236, 
        n62888, n64207, n63844, n64205, n63798, n64151, n59955, 
        n64298, n25994, n3167, n52608, n52493, n3168, n52607, 
        n3169, n52606, n26052, n62396, n3170, n52605, n2490, n52492, 
        n2491, n52491, n3171, n52604, n52412, n3172, n52603, n62402, 
        n52602, n60139, n28169, n29516, n14_adj_5249, n15_adj_5250, 
        n52601, n52600, n52599, n62752, n62758, n62768, n62774, 
        n52598, n62736, n62742, n62398, n62390, n60163, n52411, 
        n52597, n62816, n62822, n62800, n62806, n52410, n69702, 
        n26061, n52596, n1560, n52409;
    wire [23:0]n8695;
    
    wire n2353, n52490, n52595, n30, n52594, n67580, n2354, n52489, 
        n32, n8_adj_5251, n52593, n12_adj_5252, n68050, n14_adj_5253, 
        n69509, n26078, n10_adj_5254, n69511, n64246, n67158, n63964, 
        n62380, n48, n34_adj_5255, n2355, n52488, n52592, n11684, 
        n52591, n52487, n52590;
    wire [23:0]n8513;
    
    wire n1408, n52408, n52589, n63384, n960, n11848, n21444, 
        n44_adj_5256, n1409, n52407, n11855, n44_adj_5257, n48_adj_5258, 
        n44_adj_5259, n67315, n962, n48_adj_5260, n26011, n67321, 
        n42_adj_5261, n40_adj_5262, n62382, n48_adj_5263, n32_adj_5264, 
        n63820, n63776, n62908, n62928, n63804, n63846, n63802, 
        n52486, n62484, n63580, n3_adj_5265, n63584, n52588, n5, 
        n63588, n8_adj_5266, n61499, n62496, n52406, n52587, n62502, 
        n52586, n64185, n64286;
    wire [2:0]r_SM_Main_2__N_3575;
    
    wire n2, n12058, n52485, n67032, n52585, n63860, n63768, n63766, 
        n52405, n52484, n52584, n52483, n52583, n52582, n52404, 
        n52581, n52482, n52481, n52480, n52403, n52402, n52479, 
        n62400, n52478, n1415, n52401, n52580, n52579, n60189, 
        n52578;
    wire [23:0]n8487;
    
    wire n1261, n52400, n2366, n52477, n52577, n52576, n2367, 
        n52476, n1262, n52399, n62388, n60167, n52575, n1263, 
        n52398;
    wire [23:0]n8669;
    
    wire n2227, n52475, n52574, n52573, n52572, n1264, n52397, 
        n52571, n2228, n52474, n2229, n52473, n52396, n52570, 
        n52569, n52568, n52472, n52471, n52567, n52470, n52395, 
        n52566, n52565, n52469, n52468, n52564, n52563, n1267, 
        n52394, n52562, n52467, n52561, n60193, n52466, n52465;
    wire [23:0]n8461;
    
    wire n1111, n52393, n52560, n52464, n52559, n1112, n52392, 
        n52558, n52557, n52556, n1113, n52391, n2239, n52463, 
        n52390, n52555, n52554, n52389, n52553, n2240, n52462, 
        n62386, n1116, n52388;
    wire [23:0]n8643;
    
    wire n2098, n52461, n2099, n52460, n62378, n52552, n2100, 
        n52459, n52458, n52551, n52550, n52549, n52457, n52548, 
        n52547, n52456, n52546, n48_adj_5267, n26014, n52455, n52545, 
        n52544, n52454, n52543, n52453, n52542, n52452, n2108, 
        n52451, n2109, n52450, n2110, n1966, n52449, n52541, n52540, 
        n1967, n52448, n52539, n52538, n52537, n52536, n1968, 
        n52447, n52446, n52535, n52534, n52445, n52533, n52532, 
        n52444, n52531, n52443, n52530, n52442, n52529, n52441, 
        n52528, n52440, n52527, n18_adj_5268, n62288, n67418, n20_adj_5269, 
        n22_adj_5270, n67425, n62344, n6, n20_adj_5271, n52526, 
        n67450, n22_adj_5272, n24_adj_5273, n48_adj_5274, n18_adj_5275, 
        n1976, n67456, n62890, n48_adj_5276, n69614, n66996, n66993, 
        n69777, n26037, n62784, n62790, n48_adj_5277, n26_adj_5278, 
        n28, n67560, n30_adj_5279, n69747, n68936, n63978, n22_adj_5280, 
        n67474, n24_adj_5281, n67483, n26_adj_5282, n24_adj_5283, 
        n67507, n48_adj_5284, n63756, n26_adj_5285, n67514, n66991, 
        n66988, n66985, n62456, n62462, n28_adj_5286, n69650, n62834, 
        n62840, n28_adj_5287, n67531, n30_adj_5288, n37_adj_5289, 
        n43_adj_5290, n41_adj_5291, n39_adj_5292, n31_adj_5293, n33_adj_5294, 
        n35_adj_5295, n27_adj_5296, n29_adj_5297, n27_adj_5298, n67548, 
        n38_adj_5299, n60174, n26_adj_5300, n69193, n69194, n67537, 
        n69623, n68383, n69819, n69820, n48_adj_5301, n63854, n63852, 
        n63862, n43_adj_5302, n23_adj_5303, n67516, n67510, n22_adj_5304, 
        n30_adj_5305, n34_adj_5306, n69625, n69626, n69499, n69314, 
        n69412, n68395, n69649, n62438, n19_adj_5308, n21_adj_5309, 
        n21_adj_5310, n67486, n67476, n20_adj_5311, n28_adj_5312, 
        n32_adj_5313, n69720, n69721, n69606, n69231, n69722, n69535, 
        n69829, n69830, n69741, n27_adj_5314, n67570, n38_adj_5315, 
        n63962, n63800, n63960, n69199, n69200, n67564, n69619, 
        n68375, n69857, n69858, n69779, n19_adj_5316, n67459, n67454, 
        n69227, n69406, n69407, n68313, n26_adj_5317, n42_adj_5318, 
        n30_adj_5319, n69724, n69725, n69602, n68315, n68934, n69543, 
        n23_adj_5320, n25_adj_5321, n17_adj_5322, n67427, n67423, 
        n69223, n16_adj_5323, n69402, n69403, n68283, n68937, n69270, 
        n28_adj_5324, n63786, n69726, n69727, n69600, n68287, n69400, 
        n69547, n69746, n48_adj_5325, n37_adj_5326, n39_adj_5327, 
        n48_adj_5328, n43_adj_5329, n41_adj_5330, n961, n41_adj_5331, 
        n36_adj_5332, n40_adj_5333, n69617, n69618, n69515, n63850, 
        n63832, n63760, n63758, n63380, n63408, n69910, n46, n59901, 
        n63392, n805, n60200, n42_adj_5334, n69217, n959, n69218, 
        n59907, n43_adj_5335, n37_adj_5336, n63830, n63754, n60183, 
        n32_adj_5337, n69207, n69208, n68498, n69241, n68366, n69508, 
        n43_adj_5338, n64228, n69209, n69210, n68508, n69239, n68359, 
        n69510, n42_adj_5339, n43_adj_5340, n38_adj_5341, n42_adj_5342, 
        n69613, n42_adj_5343, n69221, n803, n69222, n59905, n62698, 
        n64222, n63958, n62726, n64155, n64292, n64282, n21446, 
        n41_adj_5344, n39_adj_5345, n29_adj_5346, n31_adj_5347, n23_adj_5348, 
        n25_adj_5349, n33_adj_5350, n35_adj_5351, n37_adj_5352, n7, 
        n45_adj_5353, n43_adj_5354, n11_adj_5355, n13_adj_5356, n15_adj_5357, 
        n27_adj_5358, n9, n17_adj_5359, n19_adj_5360, n21_adj_5361, 
        n67985, n68003, n16_adj_5362, n67930, n8_adj_5363, n24_adj_5364, 
        n3274, n68018, n64171, n68780, n68776, n69673, n69113, 
        n69752, n12_adj_5365, n48_adj_5366, n4_adj_5367, n62318, n69159, 
        n69160, n61397, n67977, n10_adj_5368, n30_adj_5369, n62642, 
        n67979, n69635, n62660, n68415, n69825, n69826, n6_adj_5370, 
        n64294, n69169, n60673, n62902, n62904, n69170, n67958, 
        n69310, n68413, n69769, n67960, n69710, n68421, n62330, 
        n3253, n69712, n62338, n62968, n66965, n66966, n46_adj_5371, 
        n33_adj_5372, n31_adj_5373, n46_adj_5374, n37_adj_5375, n35_adj_5376, 
        n45_adj_5377, n25_adj_5378, n27_adj_5379, n21_adj_5380, n23_adj_5381, 
        n69211, n69212, n9_adj_5382, n68516, n11_adj_5383, n19_adj_5384, 
        n38_adj_5385, n68357, n69237, n13_adj_5386, n15_adj_5387, 
        n17_adj_5388, n29_adj_5389, n67148, n68079, n68816, n68814, 
        n67150, n6_adj_5390, n69372, n31_adj_5391, n32_adj_5392, n69373, 
        n68055, n69627, n30_adj_5393, n33_adj_5394, n69374, n35_adj_5395, 
        n69375, n68067, n69306, n24_adj_5396, n69131, n29_adj_5397, 
        n67586, n40_adj_5398, n28_adj_5399, n69201, n69202, n67582, 
        n69607, n69821, n69492, n69891, n68373, n69892, n69882, 
        n69815, n69816, n69701;
    
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8825[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51603_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3617[12] ), 
            .I2(n5254), .I3(\o_Rx_DV_N_3617[8] ), .O(n67016));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51603_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i51700_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3617[12] ), .I2(n58782), 
            .I3(r_SM_Main[0]), .O(n67022));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51700_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i48100_1_lut (.I0(n64264), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60197));
    defparam i48100_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51600_4_lut (.I0(n67016), .I1(\o_Rx_DV_N_3617[24] ), .I2(n29), 
            .I3(n23), .O(n67013));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51600_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8825[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8825[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8825[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2860_3 (.CI(n52438), .I0(n1977), .I1(n858), .CO(n52439));
    SB_LUT4 i51608_4_lut (.I0(n67022), .I1(\o_Rx_DV_N_3617[24] ), .I2(n29), 
            .I3(n23), .O(n67019));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51608_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 add_2866_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n52524), 
            .O(n8773[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n67019), .I1(n67013), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 add_2860_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8617[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8825[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8825[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2860_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52438));
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8825[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8825[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2866_3 (.CI(n52524), .I0(n2730), .I1(n858), .CO(n52525));
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8825[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8825[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47823_1_lut (.I0(n63984), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60171));
    defparam i47823_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8825[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8825[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8825[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8825[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8825[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8825[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8825[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8825[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8825[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51017_4_lut (.I0(n31), .I1(n19), .I2(n17), .I3(n15), .O(n67191));
    defparam i51017_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51935_4_lut (.I0(n13), .I1(n11), .I2(n3065), .I3(baudrate[2]), 
            .O(n68109));
    defparam i51935_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52657_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n68109), 
            .O(n68832));
    defparam i52657_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52655_4_lut (.I0(n25), .I1(n23_adj_5124), .I2(n21), .I3(n68832), 
            .O(n68830));
    defparam i52655_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51019_4_lut (.I0(n31), .I1(n29_adj_5126), .I2(n27_adj_5125), 
            .I3(n68830), .O(n67193));
    defparam i51019_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53205_3_lut (.I0(n8), .I1(baudrate[13]), .I2(n31), .I3(GND_net), 
            .O(n69380));   // verilog/uart_rx.v(119[33:55])
    defparam i53205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53206_3_lut (.I0(n69380), .I1(baudrate[14]), .I2(n33), .I3(GND_net), 
            .O(n69381));   // verilog/uart_rx.v(119[33:55])
    defparam i53206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16), .I1(baudrate[17]), 
            .I2(n39), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51013_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67191), 
            .O(n67187));
    defparam i51013_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53561_4_lut (.I0(n34), .I1(n14), .I2(n39), .I3(n67182), 
            .O(n69736));   // verilog/uart_rx.v(119[33:55])
    defparam i53561_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53120_3_lut (.I0(n69381), .I1(baudrate[15]), .I2(n35), .I3(GND_net), 
            .O(n69295));   // verilog/uart_rx.v(119[33:55])
    defparam i53120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53207_3_lut (.I0(n10), .I1(baudrate[10]), .I2(n25), .I3(GND_net), 
            .O(n69382));   // verilog/uart_rx.v(119[33:55])
    defparam i53207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53208_3_lut (.I0(n69382), .I1(baudrate[11]), .I2(n27_adj_5125), 
            .I3(GND_net), .O(n69383));   // verilog/uart_rx.v(119[33:55])
    defparam i53208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51923_4_lut (.I0(n27_adj_5125), .I1(n25), .I2(n23_adj_5124), 
            .I3(n67203), .O(n68097));
    defparam i51923_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12), .I1(baudrate[9]), 
            .I2(n23_adj_5124), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53118_3_lut (.I0(n69383), .I1(baudrate[12]), .I2(n29_adj_5126), 
            .I3(GND_net), .O(n69293));   // verilog/uart_rx.v(119[33:55])
    defparam i53118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52964_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67193), 
            .O(n69139));
    defparam i52964_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53692_4_lut (.I0(n69295), .I1(n69736), .I2(n39), .I3(n67187), 
            .O(n69867));   // verilog/uart_rx.v(119[33:55])
    defparam i53692_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53123_4_lut (.I0(n69293), .I1(n20), .I2(n29_adj_5126), .I3(n68097), 
            .O(n69298));   // verilog/uart_rx.v(119[33:55])
    defparam i53123_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53714_4_lut (.I0(n69298), .I1(n69867), .I2(n39), .I3(n69139), 
            .O(n69889));   // verilog/uart_rx.v(119[33:55])
    defparam i53714_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53715_3_lut (.I0(n69889), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n69890));   // verilog/uart_rx.v(119[33:55])
    defparam i53715_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53709_3_lut (.I0(n69890), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n69884));   // verilog/uart_rx.v(119[33:55])
    defparam i53709_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53125_3_lut (.I0(n69884), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n69300));   // verilog/uart_rx.v(119[33:55])
    defparam i53125_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8799[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8799[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8799[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8799[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8799[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8799[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8799[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8799[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8799[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8799[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8799[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8799[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8799[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28324), 
            .D(n479[1]), .R(n60053));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8799[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8799[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8799[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28324), 
            .D(n479[2]), .R(n60053));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8799[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8799[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51074_4_lut (.I0(n33_adj_5138), .I1(n21_adj_5137), .I2(n19_adj_5136), 
            .I3(n17_adj_5135), .O(n67248));
    defparam i51074_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51977_4_lut (.I0(n15_adj_5140), .I1(n13_adj_5139), .I2(n2956), 
            .I3(baudrate[2]), .O(n68151));
    defparam i51977_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52677_4_lut (.I0(n21_adj_5137), .I1(n19_adj_5136), .I2(n17_adj_5135), 
            .I3(n68151), .O(n68852));
    defparam i52677_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52675_4_lut (.I0(n27_adj_5134), .I1(n25_adj_5133), .I2(n23_adj_5132), 
            .I3(n68852), .O(n68850));
    defparam i52675_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51076_4_lut (.I0(n33_adj_5138), .I1(n31_adj_5131), .I2(n29_adj_5130), 
            .I3(n68850), .O(n67250));
    defparam i51076_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53211_3_lut (.I0(n10_adj_5141), .I1(baudrate[13]), .I2(n33_adj_5138), 
            .I3(GND_net), .O(n69386));   // verilog/uart_rx.v(119[33:55])
    defparam i53211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53212_3_lut (.I0(n69386), .I1(baudrate[14]), .I2(n35_adj_5128), 
            .I3(GND_net), .O(n69387));   // verilog/uart_rx.v(119[33:55])
    defparam i53212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18), .I1(baudrate[17]), 
            .I2(n41), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51069_4_lut (.I0(n39_adj_5129), .I1(n37_adj_5127), .I2(n35_adj_5128), 
            .I3(n67248), .O(n67243));
    defparam i51069_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53559_4_lut (.I0(n36), .I1(n16_adj_5142), .I2(n41), .I3(n67238), 
            .O(n69734));   // verilog/uart_rx.v(119[33:55])
    defparam i53559_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53114_3_lut (.I0(n69387), .I1(baudrate[15]), .I2(n37_adj_5127), 
            .I3(GND_net), .O(n69289));   // verilog/uart_rx.v(119[33:55])
    defparam i53114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5143), .I1(baudrate[9]), 
            .I2(n25_adj_5133), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53557_4_lut (.I0(n22), .I1(n12_adj_5144), .I2(n25_adj_5133), 
            .I3(n67258), .O(n69732));   // verilog/uart_rx.v(119[33:55])
    defparam i53557_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53558_3_lut (.I0(n69732), .I1(baudrate[10]), .I2(n27_adj_5134), 
            .I3(GND_net), .O(n69733));   // verilog/uart_rx.v(119[33:55])
    defparam i53558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53417_3_lut (.I0(n69733), .I1(baudrate[11]), .I2(n29_adj_5130), 
            .I3(GND_net), .O(n69592));   // verilog/uart_rx.v(119[33:55])
    defparam i53417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52974_4_lut (.I0(n39_adj_5129), .I1(n37_adj_5127), .I2(n35_adj_5128), 
            .I3(n67250), .O(n69149));
    defparam i52974_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53690_4_lut (.I0(n69289), .I1(n69734), .I2(n41), .I3(n67243), 
            .O(n69865));   // verilog/uart_rx.v(119[33:55])
    defparam i53690_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53383_3_lut (.I0(n69592), .I1(baudrate[12]), .I2(n31_adj_5131), 
            .I3(GND_net), .O(n69558));   // verilog/uart_rx.v(119[33:55])
    defparam i53383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53718_4_lut (.I0(n69558), .I1(n69865), .I2(n41), .I3(n69149), 
            .O(n69893));   // verilog/uart_rx.v(119[33:55])
    defparam i53718_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53719_3_lut (.I0(n69893), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n69894));   // verilog/uart_rx.v(119[33:55])
    defparam i53719_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53713_3_lut (.I0(n69894), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n69888));   // verilog/uart_rx.v(119[33:55])
    defparam i53713_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8799[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8825[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8851[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8773[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8773[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8773[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8773[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8773[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8773[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8773[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8773[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8773[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8773[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8773[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8773[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8773[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8773[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8773[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8773[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8773[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8773[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51136_4_lut (.I0(n35_adj_5158), .I1(n23_adj_5157), .I2(n21_adj_5156), 
            .I3(n19_adj_5155), .O(n67310));
    defparam i51136_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52067_4_lut (.I0(n17_adj_5154), .I1(n15_adj_5153), .I2(n2844), 
            .I3(baudrate[2]), .O(n68241));
    defparam i52067_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52689_4_lut (.I0(n23_adj_5157), .I1(n21_adj_5156), .I2(n19_adj_5155), 
            .I3(n68241), .O(n68864));
    defparam i52689_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52687_4_lut (.I0(n29_adj_5152), .I1(n27_adj_5151), .I2(n25_adj_5150), 
            .I3(n68864), .O(n68862));
    defparam i52687_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48108_1_lut (.I0(n64272), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60147));
    defparam i48108_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51139_4_lut (.I0(n35_adj_5158), .I1(n33_adj_5149), .I2(n31_adj_5148), 
            .I3(n68862), .O(n67313));
    defparam i51139_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53217_3_lut (.I0(n12_adj_5159), .I1(baudrate[13]), .I2(n35_adj_5158), 
            .I3(GND_net), .O(n69392));   // verilog/uart_rx.v(119[33:55])
    defparam i53217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5160), .I1(baudrate[17]), 
            .I2(n43), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53218_3_lut (.I0(n69392), .I1(baudrate[14]), .I2(n37_adj_5146), 
            .I3(GND_net), .O(n69393));   // verilog/uart_rx.v(119[33:55])
    defparam i53218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51131_4_lut (.I0(n41_adj_5147), .I1(n39_adj_5145), .I2(n37_adj_5146), 
            .I3(n67310), .O(n67305));
    defparam i51131_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53215_4_lut (.I0(n38), .I1(n18_adj_5161), .I2(n43), .I3(n67302), 
            .O(n69390));   // verilog/uart_rx.v(119[33:55])
    defparam i53215_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53106_3_lut (.I0(n69393), .I1(baudrate[15]), .I2(n39_adj_5145), 
            .I3(GND_net), .O(n69281));   // verilog/uart_rx.v(119[33:55])
    defparam i53106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2859_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n52437), 
            .O(n8591[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5162), .I1(baudrate[9]), 
            .I2(n27_adj_5151), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53555_4_lut (.I0(n24), .I1(n14_adj_5163), .I2(n27_adj_5151), 
            .I3(n67332), .O(n69730));   // verilog/uart_rx.v(119[33:55])
    defparam i53555_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53556_3_lut (.I0(n69730), .I1(baudrate[10]), .I2(n29_adj_5152), 
            .I3(GND_net), .O(n69731));   // verilog/uart_rx.v(119[33:55])
    defparam i53556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53419_3_lut (.I0(n69731), .I1(baudrate[11]), .I2(n31_adj_5148), 
            .I3(GND_net), .O(n69594));   // verilog/uart_rx.v(119[33:55])
    defparam i53419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53008_4_lut (.I0(n41_adj_5147), .I1(n39_adj_5145), .I2(n37_adj_5146), 
            .I3(n67313), .O(n69183));
    defparam i53008_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53609_4_lut (.I0(n69281), .I1(n69390), .I2(n43), .I3(n67305), 
            .O(n69784));   // verilog/uart_rx.v(119[33:55])
    defparam i53609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53381_3_lut (.I0(n69594), .I1(baudrate[12]), .I2(n33_adj_5149), 
            .I3(GND_net), .O(n69556));   // verilog/uart_rx.v(119[33:55])
    defparam i53381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53684_4_lut (.I0(n69556), .I1(n69784), .I2(n43), .I3(n69183), 
            .O(n69859));   // verilog/uart_rx.v(119[33:55])
    defparam i53684_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53685_3_lut (.I0(n69859), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n69860));   // verilog/uart_rx.v(119[33:55])
    defparam i53685_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2859_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n52436), 
            .O(n8591[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8747[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8747[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8747[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8747[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8747[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8747[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8747[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8747[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8747[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8747[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3_adj_5170), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8747[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8747[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8747[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8747[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8747[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8747[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8747[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2866_2_lut (.I0(n60155), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62394)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2866_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52524));
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2859_12 (.CI(n52436), .I0(n1832), .I1(n2013), .CO(n52437));
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2865_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n52523), 
            .O(n8747[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2859_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n52435), 
            .O(n8591[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51178_4_lut (.I0(n37_adj_5178), .I1(n25_adj_5177), .I2(n23_adj_5176), 
            .I3(n21_adj_5175), .O(n67352));
    defparam i51178_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52101_4_lut (.I0(n19_adj_5174), .I1(n17_adj_5173), .I2(n2729), 
            .I3(baudrate[2]), .O(n68275));
    defparam i52101_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52703_4_lut (.I0(n25_adj_5177), .I1(n23_adj_5176), .I2(n21_adj_5175), 
            .I3(n68275), .O(n68878));
    defparam i52703_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_2865_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n52522), 
            .O(n8747[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52701_4_lut (.I0(n31_adj_5169), .I1(n29_adj_5168), .I2(n27_adj_5167), 
            .I3(n68878), .O(n68876));
    defparam i52701_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51180_4_lut (.I0(n37_adj_5178), .I1(n35_adj_5172), .I2(n33_adj_5171), 
            .I3(n68876), .O(n67354));
    defparam i51180_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53221_3_lut (.I0(n14_adj_5179), .I1(baudrate[13]), .I2(n37_adj_5178), 
            .I3(GND_net), .O(n69396));   // verilog/uart_rx.v(119[33:55])
    defparam i53221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53222_3_lut (.I0(n69396), .I1(baudrate[14]), .I2(n39_adj_5165), 
            .I3(GND_net), .O(n69397));   // verilog/uart_rx.v(119[33:55])
    defparam i53222_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2859_11 (.CI(n52435), .I0(n1833), .I1(n1879), .CO(n52436));
    SB_CARRY add_2865_18 (.CI(n52522), .I0(n2597), .I1(n2754), .CO(n52523));
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5180), .I1(baudrate[17]), 
            .I2(n45), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51174_4_lut (.I0(n43_adj_5166), .I1(n41_adj_5164), .I2(n39_adj_5165), 
            .I3(n67352), .O(n67348));
    defparam i51174_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52766_4_lut (.I0(n40), .I1(n20_adj_5181), .I2(n45), .I3(n67345), 
            .O(n68941));   // verilog/uart_rx.v(119[33:55])
    defparam i52766_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53102_3_lut (.I0(n69397), .I1(baudrate[15]), .I2(n41_adj_5164), 
            .I3(GND_net), .O(n69277));   // verilog/uart_rx.v(119[33:55])
    defparam i53102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5182), .I1(baudrate[9]), 
            .I2(n29_adj_5168), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2865_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n52521), 
            .O(n8747[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53553_4_lut (.I0(n26), .I1(n16_adj_5183), .I2(n29_adj_5168), 
            .I3(n67367), .O(n69728));   // verilog/uart_rx.v(119[33:55])
    defparam i53553_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2865_17 (.CI(n52521), .I0(n2598), .I1(n2638), .CO(n52522));
    SB_LUT4 i53554_3_lut (.I0(n69728), .I1(baudrate[10]), .I2(n31_adj_5169), 
            .I3(GND_net), .O(n69729));   // verilog/uart_rx.v(119[33:55])
    defparam i53554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2859_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n52434), 
            .O(n8591[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53421_3_lut (.I0(n69729), .I1(baudrate[11]), .I2(n33_adj_5171), 
            .I3(GND_net), .O(n69596));   // verilog/uart_rx.v(119[33:55])
    defparam i53421_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2859_10 (.CI(n52434), .I0(n1834), .I1(n1742), .CO(n52435));
    SB_LUT4 add_2865_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n52520), 
            .O(n8747[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53020_4_lut (.I0(n43_adj_5166), .I1(n41_adj_5164), .I2(n39_adj_5165), 
            .I3(n67354), .O(n69195));
    defparam i53020_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53377_4_lut (.I0(n69277), .I1(n68941), .I2(n45), .I3(n67348), 
            .O(n69552));   // verilog/uart_rx.v(119[33:55])
    defparam i53377_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2859_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n52433), 
            .O(n8591[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2859_9 (.CI(n52433), .I0(n1835), .I1(n1602), .CO(n52434));
    SB_LUT4 i53376_3_lut (.I0(n69596), .I1(baudrate[12]), .I2(n35_adj_5172), 
            .I3(GND_net), .O(n69551));   // verilog/uart_rx.v(119[33:55])
    defparam i53376_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2865_16 (.CI(n52520), .I0(n2599), .I1(n2519), .CO(n52521));
    SB_LUT4 i53379_4_lut (.I0(n69551), .I1(n69552), .I2(n45), .I3(n69195), 
            .O(n69554));   // verilog/uart_rx.v(119[33:55])
    defparam i53379_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2865_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n52519), 
            .O(n8747[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2859_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n52432), 
            .O(n8591[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2865_15 (.CI(n52519), .I0(n2600), .I1(n2397), .CO(n52520));
    SB_CARRY add_2859_8 (.CI(n52432), .I0(n1836), .I1(n1459), .CO(n52433));
    SB_LUT4 add_2865_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n52518), 
            .O(n8747[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2865_14 (.CI(n52518), .I0(n2601), .I1(n2272), .CO(n52519));
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2865_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n52517), 
            .O(n8747[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2865_13 (.CI(n52517), .I0(n2602), .I1(n2144), .CO(n52518));
    SB_LUT4 add_2865_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n52516), 
            .O(n8747[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2859_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n52431), 
            .O(n8591[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2865_12 (.CI(n52516), .I0(n2603), .I1(n2013), .CO(n52517));
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2865_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n52515), 
            .O(n8747[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2859_7 (.CI(n52431), .I0(n1837), .I1(n1460), .CO(n52432));
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2865_11 (.CI(n52515), .I0(n2604), .I1(n1879), .CO(n52516));
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2859_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n52430), 
            .O(n8591[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2865_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n52514), 
            .O(n8747[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2865_10 (.CI(n52514), .I0(n2605), .I1(n1742), .CO(n52515));
    SB_CARRY add_2859_6 (.CI(n52430), .I0(n1838), .I1(n1011), .CO(n52431));
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2865_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n52513), 
            .O(n8747[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2859_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n52429), 
            .O(n8591[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2865_9 (.CI(n52513), .I0(n2606), .I1(n1602), .CO(n52514));
    SB_LUT4 add_2865_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n52512), 
            .O(n8747[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2859_5 (.CI(n52429), .I0(n1839), .I1(n856), .CO(n52430));
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2865_8 (.CI(n52512), .I0(n2607), .I1(n1459), .CO(n52513));
    SB_LUT4 i48022_2_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n64187));
    defparam i48022_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2859_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n52428), 
            .O(n8591[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29776_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44073));
    defparam i29776_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_2865_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n52511), 
            .O(n8747[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29774_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44071));
    defparam i29774_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7335_4_lut (.I0(n804), .I1(n44071), .I2(n21434), .I3(baudrate[2]), 
            .O(n21436));   // verilog/uart_rx.v(119[33:55])
    defparam i7335_4_lut.LUT_INIT = 16'ha2aa;
    SB_CARRY add_2865_7 (.CI(n52511), .I0(n2608), .I1(n1460), .CO(n52512));
    SB_LUT4 add_2865_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n52510), 
            .O(n8747[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Clock_Count_2062_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n52815), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2865_6 (.CI(n52510), .I0(n2609), .I1(n1011), .CO(n52511));
    SB_CARRY add_2859_4 (.CI(n52428), .I0(n1840), .I1(n698), .CO(n52429));
    SB_LUT4 add_2865_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n52509), 
            .O(n8747[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2062_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n52814), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_8 (.CI(n52814), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n52815));
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n30256));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n30255));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n30254));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n30253));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n30252));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n71130));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2865_5 (.CI(n52509), .I0(n2610), .I1(n856), .CO(n52510));
    SB_LUT4 add_2865_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n52508), 
            .O(n8747[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2859_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n52427), 
            .O(n8591[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2859_3 (.CI(n52427), .I0(n1841), .I1(n858), .CO(n52428));
    SB_CARRY add_2865_4 (.CI(n52508), .I0(n2611), .I1(n698), .CO(n52509));
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n51522), .O(\o_Rx_DV_N_3617[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i44011_1_lut (.I0(n26081), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60143));
    defparam i44011_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n62352), .I1(n25975), .I2(VCC_net), 
            .I3(n51521), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n51521), .I0(n25975), .I1(VCC_net), 
            .CO(n51522));
    SB_LUT4 sub_38_add_2_24_lut (.I0(n62432), .I1(n64302), .I2(VCC_net), 
            .I3(n51520), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 r_Clock_Count_2062_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n52813), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2859_2_lut (.I0(n60180), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62384)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2859_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2865_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n52507), 
            .O(n8747[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2859_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52427));
    SB_CARRY r_Clock_Count_2062_add_4_7 (.CI(n52813), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n52814));
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Clock_Count_2062_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n52812), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_6 (.CI(n52812), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n52813));
    SB_LUT4 r_Clock_Count_2062_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n52811), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_5 (.CI(n52811), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n52812));
    SB_LUT4 add_2858_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n52426), 
            .O(n8565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2062_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n52810), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2858_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n52425), 
            .O(n8565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_4 (.CI(n52810), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n52811));
    SB_CARRY add_2865_3 (.CI(n52507), .I0(n2612), .I1(n858), .CO(n52508));
    SB_LUT4 add_2865_2_lut (.I0(n60159), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62392)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2865_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 r_Clock_Count_2062_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n52809), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_3 (.CI(n52809), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n52810));
    SB_CARRY add_2865_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52507));
    SB_CARRY add_2858_10 (.CI(n52425), .I0(n1694), .I1(n1879), .CO(n52426));
    SB_CARRY sub_38_add_2_24 (.CI(n51520), .I0(n64302), .I1(VCC_net), 
            .CO(n51521));
    SB_LUT4 add_2858_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n52424), 
            .O(n8565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3617[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n51519), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2864_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n52506), 
            .O(n8721[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2062_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2062_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2062_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n52809));
    SB_CARRY add_2858_9 (.CI(n52424), .I0(n1695), .I1(n1742), .CO(n52425));
    SB_LUT4 add_2858_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n52423), 
            .O(n8565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n52505), 
            .O(n8721[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_23 (.CI(n51519), .I0(n294[21]), .I1(VCC_net), 
            .CO(n51520));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n62430), .I1(n294[20]), .I2(VCC_net), 
            .I3(n51518), .O(n62432)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_22 (.CI(n51518), .I0(n294[20]), .I1(VCC_net), 
            .CO(n51519));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n62428), .I1(n294[19]), .I2(VCC_net), 
            .I3(n51517), .O(n62430)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_21 (.CI(n51517), .I0(n294[19]), .I1(VCC_net), 
            .CO(n51518));
    SB_CARRY add_2858_8 (.CI(n52423), .I0(n1696), .I1(n1602), .CO(n52424));
    SB_LUT4 add_2858_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n52422), 
            .O(n8565[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n51516), .O(o_Rx_DV_N_3617[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_17 (.CI(n52505), .I0(n2477), .I1(n2638), .CO(n52506));
    SB_CARRY add_2858_7 (.CI(n52422), .I0(n1697), .I1(n1459), .CO(n52423));
    SB_LUT4 add_2864_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n52504), 
            .O(n8721[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n51516), .I0(n294[18]), .I1(VCC_net), 
            .CO(n51517));
    SB_CARRY add_2864_16 (.CI(n52504), .I0(n2478), .I1(n2519), .CO(n52505));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n62426), .I1(n294[17]), .I2(VCC_net), 
            .I3(n51515), .O(n62428)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_38_add_2_19 (.CI(n51515), .I0(n294[17]), .I1(VCC_net), 
            .CO(n51516));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n62424), .I1(n294[16]), .I2(VCC_net), 
            .I3(n51514), .O(n62426)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_18 (.CI(n51514), .I0(n294[16]), .I1(VCC_net), 
            .CO(n51515));
    SB_LUT4 sub_38_add_2_17_lut (.I0(n62350), .I1(n294[15]), .I2(VCC_net), 
            .I3(n51513), .O(n62352)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n51513), .I0(n294[15]), .I1(VCC_net), 
            .CO(n51514));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n62422), .I1(n294[14]), .I2(VCC_net), 
            .I3(n51512), .O(n62424)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n51512), .I0(n294[14]), .I1(VCC_net), 
            .CO(n51513));
    SB_LUT4 add_2858_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n52421), 
            .O(n8565[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3617[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n51511), .O(n62422)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2858_6 (.CI(n52421), .I0(n1698), .I1(n1460), .CO(n52422));
    SB_LUT4 add_2864_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n52503), 
            .O(n8721[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n51511), .I0(n294[13]), .I1(VCC_net), 
            .CO(n51512));
    SB_CARRY add_2864_15 (.CI(n52503), .I0(n2479), .I1(n2397), .CO(n52504));
    SB_LUT4 add_2864_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n52502), 
            .O(n8721[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2858_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n52420), 
            .O(n8565[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_14 (.CI(n52502), .I0(n2480), .I1(n2272), .CO(n52503));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n51510), .O(\o_Rx_DV_N_3617[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_14 (.CI(n51510), .I0(n294[12]), .I1(VCC_net), 
            .CO(n51511));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3617[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n51509), .O(n62350)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n51509), .I0(n294[11]), .I1(VCC_net), 
            .CO(n51510));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n51508), .O(o_Rx_DV_N_3617[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n52501), 
            .O(n8721[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n51508), .I0(n294[10]), .I1(VCC_net), 
            .CO(n51509));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n51507), .O(o_Rx_DV_N_3617[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n51507), .I0(n294[9]), .I1(VCC_net), 
            .CO(n51508));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n51506), .O(\o_Rx_DV_N_3617[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2858_5 (.CI(n52420), .I0(n1699), .I1(n1011), .CO(n52421));
    SB_CARRY sub_38_add_2_10 (.CI(n51506), .I0(n294[8]), .I1(VCC_net), 
            .CO(n51507));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n51505), .O(\o_Rx_DV_N_3617[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2858_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n52419), 
            .O(n8565[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_13 (.CI(n52501), .I0(n2481), .I1(n2144), .CO(n52502));
    SB_CARRY sub_38_add_2_9 (.CI(n51505), .I0(n294[7]), .I1(VCC_net), 
            .CO(n51506));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n51504), .O(\o_Rx_DV_N_3617[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n51504), .I0(n294[6]), .I1(VCC_net), 
            .CO(n51505));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n51503), .O(\o_Rx_DV_N_3617[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51452_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n67626));   // verilog/uart_rx.v(119[33:55])
    defparam i51452_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2858_4 (.CI(n52419), .I0(n1700), .I1(n856), .CO(n52420));
    SB_CARRY sub_38_add_2_7 (.CI(n51503), .I0(n294[5]), .I1(VCC_net), 
            .CO(n51504));
    SB_LUT4 add_2864_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n52500), 
            .O(n8721[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2858_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n52418), 
            .O(n8565[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n51502), .O(\o_Rx_DV_N_3617[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2870_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n52624), 
            .O(n8877[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n51502), .I0(n294[4]), .I1(VCC_net), 
            .CO(n51503));
    SB_CARRY add_2864_12 (.CI(n52500), .I0(n2482), .I1(n2013), .CO(n52501));
    SB_LUT4 add_2870_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n52623), 
            .O(n8877[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_24 (.CI(n52623), .I0(n3152), .I1(n3082), .CO(n52624));
    SB_LUT4 add_2870_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n52622), 
            .O(n8877[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n52499), 
            .O(n8721[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2858_3 (.CI(n52418), .I0(n1701), .I1(n698), .CO(n52419));
    SB_LUT4 add_2858_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8565[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2858_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_11 (.CI(n52499), .I0(n2483), .I1(n1879), .CO(n52500));
    SB_LUT4 i44019_1_lut (.I0(n26055), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60151));
    defparam i44019_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n51501), .O(\o_Rx_DV_N_3617[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n51501), .I0(n294[3]), .I1(VCC_net), 
            .CO(n51502));
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n51500), .O(\o_Rx_DV_N_3617[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n51500), .I0(n294[2]), .I1(VCC_net), 
            .CO(n51501));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n51499), .O(\o_Rx_DV_N_3617[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n51499), .I0(n294[1]), .I1(VCC_net), 
            .CO(n51500));
    SB_CARRY add_2870_23 (.CI(n52622), .I0(n3153), .I1(n3188), .CO(n52623));
    SB_LUT4 add_2870_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n52621), 
            .O(n8877[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2858_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n52418));
    SB_LUT4 add_2864_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n52498), 
            .O(n8721[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_22 (.CI(n52621), .I0(n3154), .I1(n3084), .CO(n52622));
    SB_LUT4 add_2857_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n52417), 
            .O(n8539[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n61327), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3617[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2870_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n52620), 
            .O(n8877[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_10 (.CI(n52498), .I0(n2484), .I1(n1742), .CO(n52499));
    SB_LUT4 add_2857_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n52416), 
            .O(n8539[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n61327), .I1(GND_net), 
            .CO(n51499));
    SB_LUT4 add_2864_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n52497), 
            .O(n8721[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_9 (.CI(n52497), .I0(n2485), .I1(n1602), .CO(n52498));
    SB_CARRY add_2870_21 (.CI(n52620), .I0(n3155), .I1(n2977), .CO(n52621));
    SB_LUT4 add_2870_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n52619), 
            .O(n8877[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n52496), 
            .O(n8721[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_20 (.CI(n52619), .I0(n3156), .I1(n2867), .CO(n52620));
    SB_LUT4 add_2870_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n52618), 
            .O(n8877[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_19 (.CI(n52618), .I0(n3157), .I1(n2754), .CO(n52619));
    SB_LUT4 add_2870_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n52617), 
            .O(n8877[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_2864_8 (.CI(n52496), .I0(n2486), .I1(n1459), .CO(n52497));
    SB_CARRY add_2870_18 (.CI(n52617), .I0(n3158), .I1(n2638), .CO(n52618));
    SB_LUT4 add_2870_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n52616), 
            .O(n8877[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2857_10 (.CI(n52416), .I0(n1553), .I1(n1742), .CO(n52417));
    SB_LUT4 i51467_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n67641));   // verilog/uart_rx.v(119[33:55])
    defparam i51467_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2870_17 (.CI(n52616), .I0(n3159), .I1(n2519), .CO(n52617));
    SB_LUT4 add_2857_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n52415), 
            .O(n8539[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n52495), 
            .O(n8721[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2857_9 (.CI(n52415), .I0(n1554), .I1(n1602), .CO(n52416));
    SB_LUT4 add_2857_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n52414), 
            .O(n8539[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2857_8 (.CI(n52414), .I0(n1555), .I1(n1459), .CO(n52415));
    SB_LUT4 add_2870_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n52615), 
            .O(n8877[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_7 (.CI(n52495), .I0(n2487), .I1(n1460), .CO(n52496));
    SB_CARRY add_2870_16 (.CI(n52615), .I0(n3160), .I1(n2397), .CO(n52616));
    SB_LUT4 add_2870_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n52614), 
            .O(n8877[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_15 (.CI(n52614), .I0(n3161), .I1(n2272), .CO(n52615));
    SB_LUT4 add_2870_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n52613), 
            .O(n8877[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_14 (.CI(n52613), .I0(n3162), .I1(n2144), .CO(n52614));
    SB_LUT4 i51440_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n67614));   // verilog/uart_rx.v(119[33:55])
    defparam i51440_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2870_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n52612), 
            .O(n8877[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_13 (.CI(n52612), .I0(n3163), .I1(n2013), .CO(n52613));
    SB_LUT4 add_2870_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n52611), 
            .O(n8877[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_12 (.CI(n52611), .I0(n3164), .I1(n1879), .CO(n52612));
    SB_LUT4 add_2864_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n52494), 
            .O(n8721[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51429_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n67603));   // verilog/uart_rx.v(119[33:55])
    defparam i51429_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2870_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n52610), 
            .O(n8877[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_11 (.CI(n52610), .I0(n3165), .I1(n1742), .CO(n52611));
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_4_lut (.I0(n4), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[1]), 
            .I3(\r_Bit_Index[0] ), .O(n62852));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_adj_989 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62852), .O(n62858));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_990 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62858), .O(n62864));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_991 (.I0(n63858), .I1(n62370), .I2(n62368), .I3(n63810), 
            .O(n26049));
    defparam i1_4_lut_adj_991.LUT_INIT = 16'hfffe;
    SB_LUT4 i44027_1_lut (.I0(n26049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60159));
    defparam i44027_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n62880));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_992 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n62884));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'heeee;
    SB_LUT4 i51460_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n67634));   // verilog/uart_rx.v(119[33:55])
    defparam i51460_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_adj_993 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n62886));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'heeee;
    SB_LUT4 add_2870_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n52609), 
            .O(n8877[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47899_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n64062));
    defparam i47899_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_994 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n64064));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 add_2857_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n52413), 
            .O(n8539[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_6 (.CI(n52494), .I0(n2488), .I1(n1011), .CO(n52495));
    SB_LUT4 i48071_4_lut (.I0(n62886), .I1(n62882), .I2(n62884), .I3(n62880), 
            .O(n64236));
    defparam i48071_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_995 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n62888));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'heeee;
    SB_LUT4 i48042_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n64207));
    defparam i48042_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i48107_4_lut (.I0(n64207), .I1(n63844), .I2(n64205), .I3(n63798), 
            .O(n64272));
    defparam i48107_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48133_4_lut (.I0(n64272), .I1(n64151), .I2(n59955), .I3(baudrate[4]), 
            .O(n64298));
    defparam i48133_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53961_4_lut (.I0(n64236), .I1(n64064), .I2(n64298), .I3(n64062), 
            .O(n64302));
    defparam i53961_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53965_3_lut (.I0(n25994), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25975));   // verilog/uart_rx.v(119[33:55])
    defparam i53965_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_4_lut (.I0(n69554), .I1(baudrate[18]), .I2(n2713), 
            .I3(n62394), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_CARRY add_2870_10 (.CI(n52609), .I0(n3166), .I1(n1602), .CO(n52610));
    SB_LUT4 add_2870_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n52608), 
            .O(n8877[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n52493), 
            .O(n8721[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_9 (.CI(n52608), .I0(n3167), .I1(n1459), .CO(n52609));
    SB_LUT4 add_2870_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n52607), 
            .O(n8877[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_8 (.CI(n52607), .I0(n3168), .I1(n1460), .CO(n52608));
    SB_LUT4 add_2870_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n52606), 
            .O(n8877[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_5 (.CI(n52493), .I0(n2489), .I1(n856), .CO(n52494));
    SB_CARRY add_2857_7 (.CI(n52413), .I0(n1556), .I1(n1460), .CO(n52414));
    SB_LUT4 i54490_2_lut_4_lut (.I0(n69554), .I1(baudrate[18]), .I2(n2713), 
            .I3(n26052), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i54490_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_996 (.I0(n69860), .I1(baudrate[19]), .I2(n2827), 
            .I3(n62396), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_996.LUT_INIT = 16'h7100;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29921));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2870_7 (.CI(n52606), .I0(n3169), .I1(n1011), .CO(n52607));
    SB_LUT4 add_2870_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n52605), 
            .O(n8877[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2864_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n52492), 
            .O(n8721[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_4 (.CI(n52492), .I0(n2490), .I1(n698), .CO(n52493));
    SB_LUT4 add_2864_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n52491), 
            .O(n8721[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_6 (.CI(n52605), .I0(n3170), .I1(n856), .CO(n52606));
    SB_LUT4 add_2870_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n52604), 
            .O(n8877[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_3 (.CI(n52491), .I0(n2491), .I1(n858), .CO(n52492));
    SB_CARRY add_2870_5 (.CI(n52604), .I0(n3171), .I1(n698), .CO(n52605));
    SB_LUT4 add_2857_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n52412), 
            .O(n8539[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2870_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n52603), 
            .O(n8877[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2870_4 (.CI(n52603), .I0(n3172), .I1(n858), .CO(n52604));
    SB_LUT4 add_2870_3_lut (.I0(n60139), .I1(GND_net), .I2(n538), .I3(n52602), 
            .O(n62402)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2870_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2870_3 (.CI(n52602), .I0(GND_net), .I1(n538), .CO(n52603));
    SB_LUT4 i54493_2_lut_4_lut (.I0(n69860), .I1(baudrate[19]), .I2(n2827), 
            .I3(n26055), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i54493_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_DFFESR r_Clock_Count_2062__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n28169), .D(n1[0]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n28169), .D(n1[1]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n28169), .D(n1[2]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n28169), .D(n1[3]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n28169), .D(n1[4]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n28169), .D(n1[5]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n28169), .D(n1[6]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2062__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n28169), .D(n1[7]), .R(n29516));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3617[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5249));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3617[12] ), .I2(n23), .I3(n5254), 
            .O(n15_adj_5250));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5250), .I1(\o_Rx_DV_N_3617[8] ), .I2(n14_adj_5249), 
            .I3(n59011), .O(n71130));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY add_2870_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n52602));
    SB_LUT4 add_2869_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n52601), 
            .O(n8851[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2869_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n52600), 
            .O(n8851[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_22 (.CI(n52600), .I0(n3047), .I1(n3188), .CO(n52601));
    SB_LUT4 add_2869_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n52599), 
            .O(n8851[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_997 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62752), .O(n62758));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_998 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62758), .O(n62764));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_CARRY add_2869_21 (.CI(n52599), .I0(n3048), .I1(n3084), .CO(n52600));
    SB_LUT4 i1_4_lut_adj_999 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62768), .O(n62774));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62774), .O(n62780));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2869_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n52598), 
            .O(n8851[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2857_6 (.CI(n52412), .I0(n1557), .I1(n1011), .CO(n52413));
    SB_CARRY add_2869_20 (.CI(n52598), .I0(n3049), .I1(n2977), .CO(n52599));
    SB_LUT4 i1_4_lut_adj_1001 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62736), .O(n62742));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1002 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62742), .O(n62748));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1003 (.I0(n69888), .I1(baudrate[20]), .I2(n2938), 
            .I3(n62398), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1003.LUT_INIT = 16'h7100;
    SB_LUT4 add_2864_2_lut (.I0(n60163), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62390)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2864_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2857_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n52411), 
            .O(n8539[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2869_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n52597), 
            .O(n8851[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_19 (.CI(n52597), .I0(n3050), .I1(n2867), .CO(n52598));
    SB_LUT4 i1_4_lut_adj_1004 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62816), .O(n62822));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_CARRY add_2857_5 (.CI(n52411), .I0(n1558), .I1(n856), .CO(n52412));
    SB_LUT4 i1_4_lut_adj_1005 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62822), .O(n62828));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62800), .O(n62806));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62806), .O(n62812));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2857_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n52410), 
            .O(n8539[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2864_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52491));
    SB_LUT4 i54502_2_lut_4_lut (.I0(n69702), .I1(baudrate[22]), .I2(n3151), 
            .I3(n26061), .O(n294[1]));
    defparam i54502_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i54496_2_lut_4_lut (.I0(n69888), .I1(baudrate[20]), .I2(n2938), 
            .I3(n64272), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i54496_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2857_4 (.CI(n52410), .I0(n1559), .I1(n698), .CO(n52411));
    SB_LUT4 add_2869_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n52596), 
            .O(n8851[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2857_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n52409), 
            .O(n8539[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n52490), 
            .O(n8695[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_18 (.CI(n52596), .I0(n3051), .I1(n2754), .CO(n52597));
    SB_LUT4 add_2869_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n52595), 
            .O(n8851[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_17 (.CI(n52595), .I0(n3052), .I1(n2638), .CO(n52596));
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2869_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n52594), 
            .O(n8851[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30854));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n55126));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2869_16 (.CI(n52594), .I0(n3053), .I1(n2519), .CO(n52595));
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30850));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i51406_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n67580));
    defparam i51406_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_2857_3 (.CI(n52409), .I0(n1560), .I1(n858), .CO(n52410));
    SB_LUT4 add_2863_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n52489), 
            .O(n8695[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2869_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n52593), 
            .O(n8851[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51876_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n68050));
    defparam i51876_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54142_2_lut_4_lut (.I0(n69509), .I1(baudrate[10]), .I2(n1693), 
            .I3(n26078), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i54142_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54336_2_lut_4_lut (.I0(n69511), .I1(baudrate[9]), .I2(n1552), 
            .I3(n64246), .O(n294[14]));
    defparam i54336_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50984_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n67158));
    defparam i50984_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n63964));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62380), .I3(n48), .O(n34_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_CARRY add_2863_16 (.CI(n52489), .I0(n2354), .I1(n2519), .CO(n52490));
    SB_CARRY add_2869_15 (.CI(n52593), .I0(n3054), .I1(n2397), .CO(n52594));
    SB_LUT4 add_2863_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n52488), 
            .O(n8695[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_15 (.CI(n52488), .I0(n2355), .I1(n2397), .CO(n52489));
    SB_LUT4 add_2869_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n52592), 
            .O(n8851[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2857_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8539[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2857_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5650_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n21434), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n11684));   // verilog/uart_rx.v(119[33:55])
    defparam i5650_2_lut_3_lut_4_lut.LUT_INIT = 16'h4445;
    SB_CARRY add_2869_14 (.CI(n52592), .I0(n3055), .I1(n2272), .CO(n52593));
    SB_CARRY add_2857_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52409));
    SB_LUT4 add_2869_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n52591), 
            .O(n8851[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n52487), 
            .O(n8695[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_13 (.CI(n52591), .I0(n3056), .I1(n2144), .CO(n52592));
    SB_LUT4 add_2869_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n52590), 
            .O(n8851[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_12 (.CI(n52590), .I0(n3057), .I1(n2013), .CO(n52591));
    SB_LUT4 add_2856_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n52408), 
            .O(n8513[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_14 (.CI(n52487), .I0(n2356), .I1(n2272), .CO(n52488));
    SB_LUT4 add_2869_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n52589), 
            .O(n8851[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1008 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n63384));
    defparam i1_2_lut_4_lut_adj_1008.LUT_INIT = 16'hfffe;
    SB_LUT4 i5823_2_lut_4_lut (.I0(n960), .I1(n11848), .I2(n21444), .I3(baudrate[3]), 
            .O(n44_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam i5823_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 add_2856_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n52407), 
            .O(n8513[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5821_2_lut_3_lut (.I0(baudrate[3]), .I1(n21444), .I2(n11848), 
            .I3(GND_net), .O(n11855));   // verilog/uart_rx.v(119[33:55])
    defparam i5821_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i5652_2_lut_4_lut (.I0(n804), .I1(n44071), .I2(n21434), .I3(baudrate[2]), 
            .O(n44_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam i5652_2_lut_4_lut.LUT_INIT = 16'ha2fb;
    SB_LUT4 i1_3_lut_4_lut (.I0(n25994), .I1(n48_adj_5258), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5259));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i51141_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5258), .I2(n25994), 
            .I3(GND_net), .O(n67315));   // verilog/uart_rx.v(119[33:55])
    defparam i51141_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5814_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11848));   // verilog/uart_rx.v(119[33:55])
    defparam i5814_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i51147_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5260), .I2(n26011), 
            .I3(GND_net), .O(n67321));   // verilog/uart_rx.v(119[33:55])
    defparam i51147_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i5645_2_lut_3_lut (.I0(n21434), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam i5645_2_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i5808_2_lut_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), 
            .I3(GND_net), .O(n40_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam i5808_2_lut_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62382), .I3(n48_adj_5263), .O(n32_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1009 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n63820));
    defparam i1_2_lut_4_lut_adj_1009.LUT_INIT = 16'hfffe;
    SB_CARRY add_2869_11 (.CI(n52589), .I0(n3058), .I1(n1879), .CO(n52590));
    SB_LUT4 i1_4_lut_adj_1010 (.I0(n63844), .I1(n63776), .I2(n62908), 
            .I3(baudrate[19]), .O(n62928));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n62928), .I1(n63804), .I2(n63846), 
            .I3(n63802), .O(n26052));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 i44023_1_lut (.I0(n26052), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n60155));
    defparam i44023_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2856_9 (.CI(n52407), .I0(n1409), .I1(n1602), .CO(n52408));
    SB_LUT4 add_2863_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n52486), 
            .O(n8695[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5257), .I2(n60937), 
            .I3(GND_net), .O(n62484));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62484), .O(n62490));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i1_4_lut_adj_1013 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3617[2] ), .I3(\o_Rx_DV_N_3617[1] ), .O(n63580));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_305_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3617[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5265));   // verilog/uart_rx.v(69[17:62])
    defparam equal_305_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(r_Clock_Count[3]), .I1(n3_adj_5265), 
            .I2(\o_Rx_DV_N_3617[4] ), .I3(n63580), .O(n63584));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hffde;
    SB_LUT4 add_2869_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n52588), 
            .O(n8851[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_305_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3617[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_305_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3617[6] ), 
            .I3(n63584), .O(n63588));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'hffde;
    SB_LUT4 equal_305_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3617[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5266));   // verilog/uart_rx.v(69[17:62])
    defparam equal_305_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(r_Clock_Count[6]), .I1(n8_adj_5266), 
            .I2(n63588), .I3(\o_Rx_DV_N_3617[7] ), .O(n58782));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n61499), .O(n62496));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'hfeff;
    SB_CARRY add_2869_10 (.CI(n52588), .I0(n3059), .I1(n1742), .CO(n52589));
    SB_LUT4 add_2856_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n52406), 
            .O(n8513[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2869_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n52587), 
            .O(n8851[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2856_8 (.CI(n52406), .I0(n1410), .I1(n1459), .CO(n52407));
    SB_CARRY add_2869_9 (.CI(n52587), .I0(n3060), .I1(n1602), .CO(n52588));
    SB_LUT4 i1_4_lut_adj_1018 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62496), .O(n62502));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2869_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n52586), 
            .O(n8851[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48020_2_lut (.I0(\o_Rx_DV_N_3617[12] ), .I1(n58782), .I2(GND_net), 
            .I3(GND_net), .O(n64185));
    defparam i48020_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48121_4_lut (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n64185), .O(n64286));
    defparam i48121_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n62502), .I1(r_SM_Main_2__N_3575[1]), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n64286), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n12058));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n12058), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3_adj_5170));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY add_2863_13 (.CI(n52486), .I0(n2357), .I1(n2144), .CO(n52487));
    SB_CARRY add_2869_8 (.CI(n52586), .I0(n3061), .I1(n1459), .CO(n52587));
    SB_LUT4 add_2863_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n52485), 
            .O(n8695[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51752_2_lut_3_lut (.I0(n25994), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n67032));   // verilog/uart_rx.v(119[33:55])
    defparam i51752_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 add_2869_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n52585), 
            .O(n8851[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1019 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n63860));
    defparam i1_2_lut_4_lut_adj_1019.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1020 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n63858));
    defparam i1_2_lut_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1021 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n63768));
    defparam i1_2_lut_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1022 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n63766));
    defparam i1_2_lut_4_lut_adj_1022.LUT_INIT = 16'hfffe;
    SB_CARRY add_2863_12 (.CI(n52485), .I0(n2358), .I1(n2013), .CO(n52486));
    SB_LUT4 add_2856_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n52405), 
            .O(n8513[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n52484), 
            .O(n8695[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2856_7 (.CI(n52405), .I0(n1411), .I1(n1460), .CO(n52406));
    SB_CARRY add_2863_11 (.CI(n52484), .I0(n2359), .I1(n1879), .CO(n52485));
    SB_CARRY add_2869_7 (.CI(n52585), .I0(n3062), .I1(n1460), .CO(n52586));
    SB_LUT4 add_2869_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n52584), 
            .O(n8851[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n52483), 
            .O(n8695[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_6 (.CI(n52584), .I0(n3063), .I1(n1011), .CO(n52585));
    SB_LUT4 add_2869_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n52583), 
            .O(n8851[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29791));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2869_5 (.CI(n52583), .I0(n3064), .I1(n856), .CO(n52584));
    SB_CARRY add_2863_10 (.CI(n52483), .I0(n2360), .I1(n1742), .CO(n52484));
    SB_LUT4 add_2869_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n52582), 
            .O(n8851[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_4 (.CI(n52582), .I0(n3065), .I1(n698), .CO(n52583));
    SB_LUT4 add_2856_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n52404), 
            .O(n8513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2869_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n52581), 
            .O(n8851[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n52482), 
            .O(n8695[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2869_3 (.CI(n52581), .I0(n3066), .I1(n858), .CO(n52582));
    SB_CARRY add_2863_9 (.CI(n52482), .I0(n2361), .I1(n1602), .CO(n52483));
    SB_LUT4 add_2863_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n52481), 
            .O(n8695[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_8 (.CI(n52481), .I0(n2362), .I1(n1459), .CO(n52482));
    SB_LUT4 add_2863_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n52480), 
            .O(n8695[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2856_6 (.CI(n52404), .I0(n1412), .I1(n1011), .CO(n52405));
    SB_LUT4 add_2856_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n52403), 
            .O(n8513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_7 (.CI(n52480), .I0(n2363), .I1(n1460), .CO(n52481));
    SB_CARRY add_2856_5 (.CI(n52403), .I0(n1413), .I1(n856), .CO(n52404));
    SB_LUT4 add_2856_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n52402), 
            .O(n8513[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2863_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n52479), 
            .O(n8695[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2856_4 (.CI(n52402), .I0(n1414), .I1(n698), .CO(n52403));
    SB_LUT4 add_2869_2_lut (.I0(n60143), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62400)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2869_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2863_6 (.CI(n52479), .I0(n2364), .I1(n1011), .CO(n52480));
    SB_CARRY add_2869_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52581));
    SB_LUT4 add_2863_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n52478), 
            .O(n8695[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2856_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n52401), 
            .O(n8513[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n52580), 
            .O(n8825[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2856_3 (.CI(n52401), .I0(n1415), .I1(n858), .CO(n52402));
    SB_LUT4 add_2868_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n52579), 
            .O(n8825[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2856_2_lut (.I0(n60189), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62382)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2856_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2868_21 (.CI(n52579), .I0(n2939), .I1(n3084), .CO(n52580));
    SB_CARRY add_2863_5 (.CI(n52478), .I0(n2365), .I1(n856), .CO(n52479));
    SB_LUT4 add_2868_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n52578), 
            .O(n8825[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_20 (.CI(n52578), .I0(n2940), .I1(n2977), .CO(n52579));
    SB_CARRY add_2856_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52401));
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2855_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n52400), 
            .O(n8487[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2863_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n52477), 
            .O(n8695[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n52577), 
            .O(n8825[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_4 (.CI(n52477), .I0(n2366), .I1(n698), .CO(n52478));
    SB_CARRY add_2868_19 (.CI(n52577), .I0(n2941), .I1(n2867), .CO(n52578));
    SB_LUT4 add_2868_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n52576), 
            .O(n8825[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_18 (.CI(n52576), .I0(n2942), .I1(n2754), .CO(n52577));
    SB_LUT4 add_2863_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n52476), 
            .O(n8695[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2855_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n52399), 
            .O(n8487[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_3 (.CI(n52476), .I0(n2367), .I1(n858), .CO(n52477));
    SB_LUT4 add_2863_2_lut (.I0(n60167), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62388)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2863_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2868_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n52575), 
            .O(n8825[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_17 (.CI(n52575), .I0(n2943), .I1(n2638), .CO(n52576));
    SB_CARRY add_2855_8 (.CI(n52399), .I0(n1262), .I1(n1459), .CO(n52400));
    SB_LUT4 add_2855_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n52398), 
            .O(n8487[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2863_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52476));
    SB_LUT4 add_2862_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n52475), 
            .O(n8669[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n52574), 
            .O(n8825[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_16 (.CI(n52574), .I0(n2944), .I1(n2519), .CO(n52575));
    SB_CARRY add_2855_7 (.CI(n52398), .I0(n1263), .I1(n1460), .CO(n52399));
    SB_LUT4 add_2868_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n52573), 
            .O(n8825[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_15 (.CI(n52573), .I0(n2945), .I1(n2397), .CO(n52574));
    SB_LUT4 add_2868_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n52572), 
            .O(n8825[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_14 (.CI(n52572), .I0(n2946), .I1(n2272), .CO(n52573));
    SB_LUT4 add_2855_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n52397), 
            .O(n8487[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n52571), 
            .O(n8825[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2862_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n52474), 
            .O(n8669[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2855_6 (.CI(n52397), .I0(n1264), .I1(n1011), .CO(n52398));
    SB_CARRY add_2868_13 (.CI(n52571), .I0(n2947), .I1(n2144), .CO(n52572));
    SB_CARRY add_2862_15 (.CI(n52474), .I0(n2228), .I1(n2397), .CO(n52475));
    SB_LUT4 add_2862_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n52473), 
            .O(n8669[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2855_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n52396), 
            .O(n8487[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n52570), 
            .O(n8825[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_12 (.CI(n52570), .I0(n2948), .I1(n2013), .CO(n52571));
    SB_LUT4 add_2868_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n52569), 
            .O(n8825[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_14 (.CI(n52473), .I0(n2229), .I1(n2272), .CO(n52474));
    SB_CARRY add_2868_11 (.CI(n52569), .I0(n2949), .I1(n1879), .CO(n52570));
    SB_LUT4 add_2868_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n52568), 
            .O(n8825[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_10 (.CI(n52568), .I0(n2950), .I1(n1742), .CO(n52569));
    SB_LUT4 add_2862_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n52472), 
            .O(n8669[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2855_5 (.CI(n52396), .I0(n1265), .I1(n856), .CO(n52397));
    SB_CARRY add_2862_13 (.CI(n52472), .I0(n2230), .I1(n2144), .CO(n52473));
    SB_LUT4 add_2862_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n52471), 
            .O(n8669[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n52567), 
            .O(n8825[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2862_12 (.CI(n52471), .I0(n2231), .I1(n2013), .CO(n52472));
    SB_CARRY add_2868_9 (.CI(n52567), .I0(n2951), .I1(n1602), .CO(n52568));
    SB_LUT4 add_2862_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n52470), 
            .O(n8669[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2855_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n52395), 
            .O(n8487[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n52566), 
            .O(n8825[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_8 (.CI(n52566), .I0(n2952), .I1(n1459), .CO(n52567));
    SB_CARRY add_2862_11 (.CI(n52470), .I0(n2232), .I1(n1879), .CO(n52471));
    SB_LUT4 add_2868_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n52565), 
            .O(n8825[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2862_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n52469), 
            .O(n8669[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2862_10 (.CI(n52469), .I0(n2233), .I1(n1742), .CO(n52470));
    SB_LUT4 add_2862_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n52468), 
            .O(n8669[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_7 (.CI(n52565), .I0(n2953), .I1(n1460), .CO(n52566));
    SB_LUT4 add_2868_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n52564), 
            .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_9 (.CI(n52468), .I0(n2234), .I1(n1602), .CO(n52469));
    SB_CARRY add_2855_4 (.CI(n52395), .I0(n1266), .I1(n698), .CO(n52396));
    SB_CARRY add_2868_6 (.CI(n52564), .I0(n2954), .I1(n1011), .CO(n52565));
    SB_LUT4 add_2868_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n52563), 
            .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_5 (.CI(n52563), .I0(n2955), .I1(n856), .CO(n52564));
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2855_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n52394), 
            .O(n8487[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n52562), 
            .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2855_3 (.CI(n52394), .I0(n1267), .I1(n858), .CO(n52395));
    SB_LUT4 add_2862_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n52467), 
            .O(n8669[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_8 (.CI(n52467), .I0(n2235), .I1(n1459), .CO(n52468));
    SB_CARRY add_2868_4 (.CI(n52562), .I0(n2956), .I1(n698), .CO(n52563));
    SB_LUT4 add_2868_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n52561), 
            .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2855_2_lut (.I0(n60193), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62380)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2855_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2862_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n52466), 
            .O(n8669[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2855_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52394));
    SB_CARRY add_2862_7 (.CI(n52466), .I0(n2236), .I1(n1460), .CO(n52467));
    SB_CARRY add_2868_3 (.CI(n52561), .I0(n2957), .I1(n858), .CO(n52562));
    SB_LUT4 add_2862_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n52465), 
            .O(n8669[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2868_2_lut (.I0(n60147), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62398)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2868_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2862_6 (.CI(n52465), .I0(n2237), .I1(n1011), .CO(n52466));
    SB_LUT4 add_2854_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n52393), 
            .O(n8461[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2868_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52561));
    SB_LUT4 add_2867_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n52560), 
            .O(n8799[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2862_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n52464), 
            .O(n8669[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2867_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n52559), 
            .O(n8799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_20 (.CI(n52559), .I0(n2828), .I1(n2977), .CO(n52560));
    SB_LUT4 add_2854_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n52392), 
            .O(n8461[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_5 (.CI(n52464), .I0(n2238), .I1(n856), .CO(n52465));
    SB_LUT4 add_2867_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n52558), 
            .O(n8799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_19 (.CI(n52558), .I0(n2829), .I1(n2867), .CO(n52559));
    SB_LUT4 add_2867_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n52557), 
            .O(n8799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_18 (.CI(n52557), .I0(n2830), .I1(n2754), .CO(n52558));
    SB_CARRY add_2854_7 (.CI(n52392), .I0(n1112), .I1(n1460), .CO(n52393));
    SB_LUT4 add_2867_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n52556), 
            .O(n8799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2854_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n52391), 
            .O(n8461[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2862_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n52463), 
            .O(n8669[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2854_6 (.CI(n52391), .I0(n1113), .I1(n1011), .CO(n52392));
    SB_CARRY add_2867_17 (.CI(n52556), .I0(n2831), .I1(n2638), .CO(n52557));
    SB_LUT4 add_2854_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n52390), 
            .O(n8461[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2867_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n52555), 
            .O(n8799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2854_5 (.CI(n52390), .I0(n1114), .I1(n856), .CO(n52391));
    SB_CARRY add_2867_16 (.CI(n52555), .I0(n2832), .I1(n2519), .CO(n52556));
    SB_LUT4 add_2867_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n52554), 
            .O(n8799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_4 (.CI(n52463), .I0(n2239), .I1(n698), .CO(n52464));
    SB_LUT4 add_2854_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n52389), 
            .O(n8461[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_15 (.CI(n52554), .I0(n2833), .I1(n2397), .CO(n52555));
    SB_CARRY add_2854_4 (.CI(n52389), .I0(n1115), .I1(n698), .CO(n52390));
    SB_LUT4 add_2867_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n52553), 
            .O(n8799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2862_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n52462), 
            .O(n8669[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2862_3 (.CI(n52462), .I0(n2240), .I1(n858), .CO(n52463));
    SB_LUT4 add_2862_2_lut (.I0(n60171), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62386)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2862_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2862_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52462));
    SB_LUT4 add_2854_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n52388), 
            .O(n8461[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2854_3 (.CI(n52388), .I0(n1116), .I1(n858), .CO(n52389));
    SB_LUT4 add_2861_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n52461), 
            .O(n8643[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2861_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n52460), 
            .O(n8643[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2854_2_lut (.I0(n60197), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62378)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2854_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2867_14 (.CI(n52553), .I0(n2834), .I1(n2272), .CO(n52554));
    SB_LUT4 add_2867_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n52552), 
            .O(n8799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2854_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52388));
    SB_CARRY add_2861_13 (.CI(n52460), .I0(n2099), .I1(n2272), .CO(n52461));
    SB_CARRY add_2867_13 (.CI(n52552), .I0(n2835), .I1(n2144), .CO(n52553));
    SB_LUT4 add_2861_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n52459), 
            .O(n8643[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_12 (.CI(n52459), .I0(n2100), .I1(n2144), .CO(n52460));
    SB_LUT4 add_2861_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n52458), 
            .O(n8643[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2867_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n52551), 
            .O(n8799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_12 (.CI(n52551), .I0(n2836), .I1(n2013), .CO(n52552));
    SB_LUT4 add_2867_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n52550), 
            .O(n8799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_11 (.CI(n52550), .I0(n2837), .I1(n1879), .CO(n52551));
    SB_CARRY add_2861_11 (.CI(n52458), .I0(n2101), .I1(n2013), .CO(n52459));
    SB_LUT4 add_2867_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n52549), 
            .O(n8799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2861_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n52457), 
            .O(n8643[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_10 (.CI(n52549), .I0(n2838), .I1(n1742), .CO(n52550));
    SB_LUT4 add_2867_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n52548), 
            .O(n8799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_9 (.CI(n52548), .I0(n2839), .I1(n1602), .CO(n52549));
    SB_LUT4 add_2867_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n52547), 
            .O(n8799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_10 (.CI(n52457), .I0(n2102), .I1(n1879), .CO(n52458));
    SB_LUT4 add_2861_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n52456), 
            .O(n8643[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_8 (.CI(n52547), .I0(n2840), .I1(n1459), .CO(n52548));
    SB_LUT4 add_2867_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n52546), 
            .O(n8799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_9 (.CI(n52456), .I0(n2103), .I1(n1742), .CO(n52457));
    SB_CARRY add_2867_7 (.CI(n52546), .I0(n2841), .I1(n1460), .CO(n52547));
    SB_LUT4 i51821_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48_adj_5267), 
            .I3(n26014), .O(n1115));
    defparam i51821_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 add_2861_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n52455), 
            .O(n8643[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2867_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n52545), 
            .O(n8799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_6 (.CI(n52545), .I0(n2842), .I1(n1011), .CO(n52546));
    SB_LUT4 add_2867_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n52544), 
            .O(n8799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_8 (.CI(n52455), .I0(n2104), .I1(n1602), .CO(n52456));
    SB_LUT4 add_2861_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n52454), 
            .O(n8643[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_7 (.CI(n52454), .I0(n2105), .I1(n1459), .CO(n52455));
    SB_CARRY add_2867_5 (.CI(n52544), .I0(n2843), .I1(n856), .CO(n52545));
    SB_LUT4 add_2867_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n52543), 
            .O(n8799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2861_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n52453), 
            .O(n8643[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_6 (.CI(n52453), .I0(n2106), .I1(n1460), .CO(n52454));
    SB_CARRY add_2867_4 (.CI(n52543), .I0(n2844), .I1(n698), .CO(n52544));
    SB_LUT4 add_2867_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n52542), 
            .O(n8799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2867_3 (.CI(n52542), .I0(n2845), .I1(n858), .CO(n52543));
    SB_LUT4 add_2867_2_lut (.I0(n60151), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n62396)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2867_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2861_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n52452), 
            .O(n8643[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_5 (.CI(n52452), .I0(n2107), .I1(n1011), .CO(n52453));
    SB_LUT4 add_2861_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n52451), 
            .O(n8643[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_4 (.CI(n52451), .I0(n2108), .I1(n856), .CO(n52452));
    SB_CARRY add_2867_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n52542));
    SB_LUT4 add_2861_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n52450), 
            .O(n8643[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_3 (.CI(n52450), .I0(n2109), .I1(n698), .CO(n52451));
    SB_LUT4 add_2861_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8643[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2861_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2861_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n52450));
    SB_LUT4 add_2860_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n52449), 
            .O(n8617[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n52541), 
            .O(n8773[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n52540), 
            .O(n8773[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_19 (.CI(n52540), .I0(n2714), .I1(n2867), .CO(n52541));
    SB_LUT4 add_2860_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n52448), 
            .O(n8617[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n52539), 
            .O(n8773[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_18 (.CI(n52539), .I0(n2715), .I1(n2754), .CO(n52540));
    SB_CARRY add_2860_13 (.CI(n52448), .I0(n1967), .I1(n2144), .CO(n52449));
    SB_LUT4 add_2866_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n52538), 
            .O(n8773[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_17 (.CI(n52538), .I0(n2716), .I1(n2638), .CO(n52539));
    SB_LUT4 add_2866_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n52537), 
            .O(n8773[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_16 (.CI(n52537), .I0(n2717), .I1(n2519), .CO(n52538));
    SB_LUT4 add_2866_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n52536), 
            .O(n8773[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2860_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n52447), 
            .O(n8617[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_12 (.CI(n52447), .I0(n1968), .I1(n2013), .CO(n52448));
    SB_LUT4 add_2860_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n52446), 
            .O(n8617[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_15 (.CI(n52536), .I0(n2718), .I1(n2397), .CO(n52537));
    SB_LUT4 add_2866_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n52535), 
            .O(n8773[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_11 (.CI(n52446), .I0(n1969), .I1(n1879), .CO(n52447));
    SB_CARRY add_2866_14 (.CI(n52535), .I0(n2719), .I1(n2272), .CO(n52536));
    SB_LUT4 add_2866_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n52534), 
            .O(n8773[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_13 (.CI(n52534), .I0(n2720), .I1(n2144), .CO(n52535));
    SB_LUT4 add_2860_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n52445), 
            .O(n8617[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n52533), 
            .O(n8773[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_12 (.CI(n52533), .I0(n2721), .I1(n2013), .CO(n52534));
    SB_LUT4 add_2866_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n52532), 
            .O(n8773[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_11 (.CI(n52532), .I0(n2722), .I1(n1879), .CO(n52533));
    SB_CARRY add_2860_10 (.CI(n52445), .I0(n1970), .I1(n1742), .CO(n52446));
    SB_LUT4 add_2860_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n52444), 
            .O(n8617[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_9 (.CI(n52444), .I0(n1971), .I1(n1602), .CO(n52445));
    SB_LUT4 add_2866_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n52531), 
            .O(n8773[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_10 (.CI(n52531), .I0(n2723), .I1(n1742), .CO(n52532));
    SB_LUT4 add_2860_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n52443), 
            .O(n8617[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_8 (.CI(n52443), .I0(n1972), .I1(n1459), .CO(n52444));
    SB_LUT4 add_2866_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n52530), 
            .O(n8773[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_9 (.CI(n52530), .I0(n2724), .I1(n1602), .CO(n52531));
    SB_LUT4 add_2860_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n52442), 
            .O(n8617[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n52529), 
            .O(n8773[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_7 (.CI(n52442), .I0(n1973), .I1(n1460), .CO(n52443));
    SB_CARRY add_2866_8 (.CI(n52529), .I0(n2725), .I1(n1459), .CO(n52530));
    SB_LUT4 add_2860_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n52441), 
            .O(n8617[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2866_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n52528), 
            .O(n8773[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2860_6 (.CI(n52441), .I0(n1974), .I1(n1011), .CO(n52442));
    SB_LUT4 add_2860_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n52440), 
            .O(n8617[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2866_7 (.CI(n52528), .I0(n2726), .I1(n1460), .CO(n52529));
    SB_LUT4 add_2866_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n52527), 
            .O(n8773[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1023 (.I0(n23), .I1(\o_Rx_DV_N_3617[12] ), .I2(n5257), 
            .I3(GND_net), .O(n62288));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_1023.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1024 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n27), .I2(n29), 
            .I3(n62288), .O(\r_SM_Main_2__N_3665[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1024.LUT_INIT = 16'hfffe;
    SB_LUT4 i51244_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n67418));
    defparam i51244_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2235_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2235_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i48096_1_lut_2_lut (.I0(baudrate[9]), .I1(n64246), .I2(GND_net), 
            .I3(GND_net), .O(n60189));
    defparam i48096_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54235_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n64246), .I2(n48), 
            .I3(baudrate[8]), .O(n294[16]));
    defparam i54235_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54264_2_lut_3_lut (.I0(baudrate[9]), .I1(n64246), .I2(n48_adj_5263), 
            .I3(GND_net), .O(n294[15]));
    defparam i54264_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i48099_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n64246), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n64264));
    defparam i48099_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48098_1_lut_2_lut_3_lut (.I0(baudrate[9]), .I1(n64246), .I2(baudrate[8]), 
            .I3(GND_net), .O(n60193));
    defparam i48098_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i51251_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n67425));
    defparam i51251_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n23), .I1(\o_Rx_DV_N_3617[12] ), .I2(n5254), 
            .I3(\o_Rx_DV_N_3617[8] ), .O(n62344));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n27), .I2(n29), 
            .I3(n62344), .O(r_SM_Main_2__N_3575[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_CARRY add_2866_6 (.CI(n52527), .I0(n2727), .I1(n1011), .CO(n52528));
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n61499));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2228_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2228_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2866_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n52526), 
            .O(n8773[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51276_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n67450));
    defparam i51276_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2860_5 (.CI(n52440), .I0(n1975), .I1(n856), .CO(n52441));
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62388), .I3(n48_adj_5274), .O(n18_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 add_2860_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n52439), 
            .O(n8617[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51282_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n67456));
    defparam i51282_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1027 (.I0(n62890), .I1(n64264), .I2(baudrate[0]), 
            .I3(n48_adj_5276), .O(n962));
    defparam i1_3_lut_4_lut_adj_1027.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_4_lut_adj_1028 (.I0(n69614), .I1(baudrate[6]), .I2(n1111), 
            .I3(n62378), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1028.LUT_INIT = 16'h7100;
    SB_CARRY add_2866_5 (.CI(n52526), .I0(n2728), .I1(n856), .CO(n52527));
    SB_LUT4 i53971_2_lut_4_lut (.I0(n69614), .I1(baudrate[6]), .I2(n1111), 
            .I3(n64264), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i53971_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51792_4_lut (.I0(\o_Rx_DV_N_3617[8] ), .I1(\o_Rx_DV_N_3617[12] ), 
            .I2(n5254), .I3(n59011), .O(n66996));
    defparam i51792_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i51788_4_lut (.I0(n66996), .I1(\o_Rx_DV_N_3617[24] ), .I2(n29), 
            .I3(n23), .O(n66993));
    defparam i51788_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n66993), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n28127));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 add_2866_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n52525), 
            .O(n8773[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2866_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54145_2_lut_4_lut (.I0(n69777), .I1(baudrate[13]), .I2(n2098), 
            .I3(n26037), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i54145_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2860_4 (.CI(n52439), .I0(n1976), .I1(n698), .CO(n52440));
    SB_LUT4 i1_4_lut_adj_1029 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62784), .O(n62790));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62790), .O(n62796));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62384), .I3(n48_adj_5277), .O(n26_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53748_2_lut_3_lut_4_lut (.I0(r_SM_Main_2__N_3575[1]), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n28324));
    defparam i53748_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i51386_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n67560));
    defparam i51386_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2860_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n52438), 
            .O(n8617[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2860_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54487_2_lut_4_lut (.I0(n69747), .I1(baudrate[17]), .I2(n2596), 
            .I3(n26049), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i54487_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1031 (.I0(n69747), .I1(baudrate[17]), .I2(n2596), 
            .I3(n62392), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1031.LUT_INIT = 16'h7100;
    SB_CARRY add_2866_4 (.CI(n52525), .I0(n2729), .I1(n698), .CO(n52526));
    SB_LUT4 i1_2_lut_4_lut_adj_1032 (.I0(n68936), .I1(baudrate[16]), .I2(n2476), 
            .I3(n62390), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1032.LUT_INIT = 16'h7100;
    SB_LUT4 i54484_2_lut_4_lut (.I0(n68936), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63978), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i54484_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51300_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n67474));
    defparam i51300_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51309_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n67483));
    defparam i51309_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54423_2_lut_3_lut_4_lut (.I0(n62882), .I1(n63984), .I2(n48_adj_5277), 
            .I3(baudrate[12]), .O(n294[12]));
    defparam i54423_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51333_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n67507));
    defparam i51333_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1033 (.I0(n62882), .I1(n63984), .I2(n8617[11]), 
            .I3(n48_adj_5284), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1033.LUT_INIT = 16'h0010;
    SB_LUT4 i48081_2_lut_3_lut_4_lut (.I0(n62882), .I1(n63984), .I2(n63756), 
            .I3(baudrate[12]), .O(n64246));
    defparam i48081_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51340_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n67514));
    defparam i51340_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51817_2_lut (.I0(n58782), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n66991));
    defparam i51817_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51814_4_lut (.I0(n66991), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3617[12] ), 
            .O(n66988));
    defparam i51814_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51279_4_lut (.I0(n66988), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3617[24] ), 
            .O(n66985));
    defparam i51279_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i54238_4_lut (.I0(\r_SM_Main[2] ), .I1(n66985), .I2(r_SM_Main_2__N_3575[1]), 
            .I3(\r_SM_Main[1] ), .O(n29516));
    defparam i54238_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n58782), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n62456));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3617[12] ), 
            .I3(n62456), .O(n62462));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h0100;
    SB_LUT4 i53751_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3617[24] ), 
            .I2(n27), .I3(n62462), .O(n28169));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i53751_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5286));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1036 (.I0(n69650), .I1(baudrate[14]), .I2(n2227), 
            .I3(n62386), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1036.LUT_INIT = 16'h7100;
    SB_LUT4 i54473_2_lut_4_lut (.I0(n69650), .I1(baudrate[14]), .I2(n2227), 
            .I3(n63984), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i54473_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(n4), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(r_Bit_Index[2]), .O(n62834));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(\o_Rx_DV_N_3617[12] ), .I1(n5254), .I2(\o_Rx_DV_N_3617[8] ), 
            .I3(n62834), .O(n62840));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5287));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51357_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n67531));
    defparam i51357_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n29), .I2(n23), 
            .I3(n62840), .O(n62846));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5288));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8721[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8617[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8643[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8669[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8695[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8721[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8695[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8721[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8591[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8617[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8643[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8669[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8695[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8721[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5289));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8695[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8721[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5290));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8591[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8617[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8643[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8669[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8695[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8721[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5291));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8591[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8617[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8643[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8669[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8695[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8721[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5292));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8591[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8617[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8643[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8669[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8695[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8591[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8617[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8643[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8669[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8695[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8721[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8591[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8617[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8643[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8669[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8695[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8721[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8721[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5293));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5294));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5295));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8591[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8617[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8643[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8669[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8695[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8591[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8617[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8643[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8669[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8695[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8721[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8721[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5296));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5297));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n62908));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n63804));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5298));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51374_4_lut (.I0(n33_adj_5186), .I1(n31_adj_5184), .I2(n29_adj_5185), 
            .I3(n27_adj_5298), .O(n67548));
    defparam i51374_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5288), .I1(baudrate[10]), 
            .I2(n41_adj_5190), .I3(GND_net), .O(n38_adj_5299));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29817_rep_4_2_lut (.I0(n8617[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n60174));   // verilog/uart_rx.v(119[33:55])
    defparam i29817_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n60174), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5300));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53018_3_lut (.I0(n26_adj_5300), .I1(baudrate[6]), .I2(n33_adj_5186), 
            .I3(GND_net), .O(n69193));   // verilog/uart_rx.v(119[33:55])
    defparam i53018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53019_3_lut (.I0(n69193), .I1(baudrate[7]), .I2(n35_adj_5187), 
            .I3(GND_net), .O(n69194));   // verilog/uart_rx.v(119[33:55])
    defparam i53019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51363_4_lut (.I0(n39_adj_5188), .I1(n37_adj_5189), .I2(n35_adj_5187), 
            .I3(n67548), .O(n67537));
    defparam i51363_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53448_4_lut (.I0(n38_adj_5299), .I1(n28_adj_5287), .I2(n41_adj_5190), 
            .I3(n67531), .O(n69623));   // verilog/uart_rx.v(119[33:55])
    defparam i53448_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52209_3_lut (.I0(n69194), .I1(baudrate[8]), .I2(n37_adj_5189), 
            .I3(GND_net), .O(n68383));   // verilog/uart_rx.v(119[33:55])
    defparam i52209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53644_4_lut (.I0(n68383), .I1(n69623), .I2(n41_adj_5190), 
            .I3(n67537), .O(n69819));   // verilog/uart_rx.v(119[33:55])
    defparam i53644_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53645_3_lut (.I0(n69819), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n69820));   // verilog/uart_rx.v(119[33:55])
    defparam i53645_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53602_3_lut (.I0(n69820), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n69777));   // verilog/uart_rx.v(119[33:55])
    defparam i53602_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52215_3_lut (.I0(n69777), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5301));   // verilog/uart_rx.v(119[33:55])
    defparam i52215_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n63854));
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1043 (.I0(n63804), .I1(n63852), .I2(n62908), 
            .I3(GND_net), .O(n63862));
    defparam i1_3_lut_adj_1043.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(n63862), .I1(n63858), .I2(n63860), 
            .I3(n63854), .O(n26037));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1045 (.I0(n26037), .I1(n48_adj_5301), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1045.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8669[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8695[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5302));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5303));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51342_4_lut (.I0(n29_adj_5191), .I1(n27_adj_5193), .I2(n25_adj_5195), 
            .I3(n23_adj_5303), .O(n67516));
    defparam i51342_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51336_4_lut (.I0(n35_adj_5194), .I1(n33_adj_5199), .I2(n31_adj_5192), 
            .I3(n67516), .O(n67510));
    defparam i51336_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5304));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5286), .I1(baudrate[7]), 
            .I2(n33_adj_5199), .I3(GND_net), .O(n30_adj_5305));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5285), .I1(baudrate[9]), 
            .I2(n37_adj_5196), .I3(GND_net), .O(n34_adj_5306));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53450_4_lut (.I0(n34_adj_5306), .I1(n24_adj_5283), .I2(n37_adj_5196), 
            .I3(n67507), .O(n69625));   // verilog/uart_rx.v(119[33:55])
    defparam i53450_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53451_3_lut (.I0(n69625), .I1(baudrate[10]), .I2(n39_adj_5197), 
            .I3(GND_net), .O(n69626));   // verilog/uart_rx.v(119[33:55])
    defparam i53451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53324_3_lut (.I0(n69626), .I1(baudrate[11]), .I2(n41_adj_5198), 
            .I3(GND_net), .O(n69499));   // verilog/uart_rx.v(119[33:55])
    defparam i53324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53139_4_lut (.I0(n41_adj_5198), .I1(n39_adj_5197), .I2(n37_adj_5196), 
            .I3(n67510), .O(n69314));
    defparam i53139_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53237_4_lut (.I0(n30_adj_5305), .I1(n22_adj_5304), .I2(n33_adj_5199), 
            .I3(n67514), .O(n69412));   // verilog/uart_rx.v(119[33:55])
    defparam i53237_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52221_3_lut (.I0(n69499), .I1(baudrate[12]), .I2(n43_adj_5302), 
            .I3(GND_net), .O(n68395));   // verilog/uart_rx.v(119[33:55])
    defparam i52221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53474_4_lut (.I0(n68395), .I1(n69412), .I2(n43_adj_5302), 
            .I3(n69314), .O(n69649));   // verilog/uart_rx.v(119[33:55])
    defparam i53474_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53475_3_lut (.I0(n69649), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n69650));   // verilog/uart_rx.v(119[33:55])
    defparam i53475_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n23), .I1(\o_Rx_DV_N_3617[12] ), .I2(n5257), 
            .I3(\r_SM_Main[0] ), .O(n62438));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(\o_Rx_DV_N_3617[24] ), .I1(n27), .I2(n29), 
            .I3(n62438), .O(n60609));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8695[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8721[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8721[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5308));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5309));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8591[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8617[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8643[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8591[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8617[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8643[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8669[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8669[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5310));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51312_4_lut (.I0(n27_adj_5200), .I1(n25_adj_5202), .I2(n23_adj_5204), 
            .I3(n21_adj_5310), .O(n67486));
    defparam i51312_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51302_4_lut (.I0(n33_adj_5203), .I1(n31_adj_5208), .I2(n29_adj_5201), 
            .I3(n67486), .O(n67476));
    defparam i51302_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_5311));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5282), .I1(baudrate[7]), 
            .I2(n31_adj_5208), .I3(GND_net), .O(n28_adj_5312));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5281), .I1(baudrate[9]), 
            .I2(n35_adj_5205), .I3(GND_net), .O(n32_adj_5313));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53545_4_lut (.I0(n32_adj_5313), .I1(n22_adj_5280), .I2(n35_adj_5205), 
            .I3(n67474), .O(n69720));   // verilog/uart_rx.v(119[33:55])
    defparam i53545_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53546_3_lut (.I0(n69720), .I1(baudrate[10]), .I2(n37_adj_5206), 
            .I3(GND_net), .O(n69721));   // verilog/uart_rx.v(119[33:55])
    defparam i53546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53431_3_lut (.I0(n69721), .I1(baudrate[11]), .I2(n39_adj_5207), 
            .I3(GND_net), .O(n69606));   // verilog/uart_rx.v(119[33:55])
    defparam i53431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53056_4_lut (.I0(n39_adj_5207), .I1(n37_adj_5206), .I2(n35_adj_5205), 
            .I3(n67476), .O(n69231));
    defparam i53056_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53547_4_lut (.I0(n28_adj_5312), .I1(n20_adj_5311), .I2(n31_adj_5208), 
            .I3(n67483), .O(n69722));   // verilog/uart_rx.v(119[33:55])
    defparam i53547_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53360_3_lut (.I0(n69606), .I1(baudrate[12]), .I2(n41_adj_5209), 
            .I3(GND_net), .O(n69535));   // verilog/uart_rx.v(119[33:55])
    defparam i53360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53654_4_lut (.I0(n69535), .I1(n69722), .I2(n41_adj_5209), 
            .I3(n69231), .O(n69829));   // verilog/uart_rx.v(119[33:55])
    defparam i53654_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53655_3_lut (.I0(n69829), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n69830));   // verilog/uart_rx.v(119[33:55])
    defparam i53655_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53566_3_lut (.I0(n69830), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n69741));   // verilog/uart_rx.v(119[33:55])
    defparam i53566_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53364_3_lut (.I0(n69741), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam i53364_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(n62388), .I1(n48_adj_5274), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8721[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8591[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8617[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8643[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8669[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8695[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n62882));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5314));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51396_4_lut (.I0(n33_adj_5212), .I1(n31_adj_5210), .I2(n29_adj_5211), 
            .I3(n27_adj_5314), .O(n67570));
    defparam i51396_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5279), .I1(baudrate[9]), 
            .I2(n41_adj_5216), .I3(GND_net), .O(n38_adj_5315));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44007_1_lut_4_lut (.I0(n63962), .I1(n63964), .I2(n63800), 
            .I3(n63960), .O(n60139));
    defparam i44007_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54406_4_lut_4_lut (.I0(r_SM_Main_2__N_3575[1]), .I1(\r_SM_Main[1] ), 
            .I2(n6), .I3(n61499), .O(n60053));
    defparam i54406_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i53024_3_lut (.I0(n26_adj_5278), .I1(baudrate[5]), .I2(n33_adj_5212), 
            .I3(GND_net), .O(n69199));   // verilog/uart_rx.v(119[33:55])
    defparam i53024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53025_3_lut (.I0(n69199), .I1(baudrate[6]), .I2(n35_adj_5213), 
            .I3(GND_net), .O(n69200));   // verilog/uart_rx.v(119[33:55])
    defparam i53025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51390_4_lut (.I0(n39_adj_5214), .I1(n37_adj_5215), .I2(n35_adj_5213), 
            .I3(n67570), .O(n67564));
    defparam i51390_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53444_4_lut (.I0(n38_adj_5315), .I1(n28), .I2(n41_adj_5216), 
            .I3(n67560), .O(n69619));   // verilog/uart_rx.v(119[33:55])
    defparam i53444_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52201_3_lut (.I0(n69200), .I1(baudrate[7]), .I2(n37_adj_5215), 
            .I3(GND_net), .O(n68375));   // verilog/uart_rx.v(119[33:55])
    defparam i52201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53682_4_lut (.I0(n68375), .I1(n69619), .I2(n41_adj_5216), 
            .I3(n67564), .O(n69857));   // verilog/uart_rx.v(119[33:55])
    defparam i53682_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53683_3_lut (.I0(n69857), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n69858));   // verilog/uart_rx.v(119[33:55])
    defparam i53683_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53604_3_lut (.I0(n69858), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n69779));   // verilog/uart_rx.v(119[33:55])
    defparam i53604_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52207_3_lut (.I0(n69779), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam i52207_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8643[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8669[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5316));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51285_4_lut (.I0(n25_adj_5217), .I1(n23_adj_5220), .I2(n21_adj_5222), 
            .I3(n19_adj_5316), .O(n67459));
    defparam i51285_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51280_4_lut (.I0(n31_adj_5221), .I1(n29_adj_5219), .I2(n27_adj_5218), 
            .I3(n67459), .O(n67454));
    defparam i51280_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53052_4_lut (.I0(n37_adj_5225), .I1(n35_adj_5224), .I2(n33_adj_5223), 
            .I3(n67454), .O(n69227));
    defparam i53052_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53231_3_lut (.I0(n18_adj_5275), .I1(baudrate[13]), .I2(n41_adj_5226), 
            .I3(GND_net), .O(n69406));   // verilog/uart_rx.v(119[33:55])
    defparam i53231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53232_3_lut (.I0(n69406), .I1(baudrate[14]), .I2(n43_adj_5227), 
            .I3(GND_net), .O(n69407));   // verilog/uart_rx.v(119[33:55])
    defparam i53232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52139_4_lut (.I0(n43_adj_5227), .I1(n41_adj_5226), .I2(n29_adj_5219), 
            .I3(n67456), .O(n68313));
    defparam i52139_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5273), .I1(baudrate[7]), 
            .I2(n29_adj_5219), .I3(GND_net), .O(n26_adj_5317));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53091_3_lut (.I0(n69407), .I1(baudrate[15]), .I2(n45_adj_5229), 
            .I3(GND_net), .O(n42_adj_5318));   // verilog/uart_rx.v(119[33:55])
    defparam i53091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48070_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n63984), .I3(baudrate[12]), .O(n60180));
    defparam i48070_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54441_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n63984), .I3(n48_adj_5284), .O(n294[11]));
    defparam i54441_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5272), .I1(baudrate[9]), 
            .I2(n33_adj_5223), .I3(GND_net), .O(n30_adj_5319));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47817_1_lut_2_lut (.I0(baudrate[17]), .I1(n26049), .I2(GND_net), 
            .I3(GND_net), .O(n60163));
    defparam i47817_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i53549_4_lut (.I0(n30_adj_5319), .I1(n20_adj_5271), .I2(n33_adj_5223), 
            .I3(n67450), .O(n69724));   // verilog/uart_rx.v(119[33:55])
    defparam i53549_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53550_3_lut (.I0(n69724), .I1(baudrate[10]), .I2(n35_adj_5224), 
            .I3(GND_net), .O(n69725));   // verilog/uart_rx.v(119[33:55])
    defparam i53550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53427_3_lut (.I0(n69725), .I1(baudrate[11]), .I2(n37_adj_5225), 
            .I3(GND_net), .O(n69602));   // verilog/uart_rx.v(119[33:55])
    defparam i53427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52141_4_lut (.I0(n43_adj_5227), .I1(n41_adj_5226), .I2(n39_adj_5228), 
            .I3(n69227), .O(n68315));
    defparam i52141_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52759_4_lut (.I0(n42_adj_5318), .I1(n26_adj_5317), .I2(n45_adj_5229), 
            .I3(n68313), .O(n68934));   // verilog/uart_rx.v(119[33:55])
    defparam i52759_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53368_3_lut (.I0(n69602), .I1(baudrate[12]), .I2(n39_adj_5228), 
            .I3(GND_net), .O(n69543));   // verilog/uart_rx.v(119[33:55])
    defparam i53368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52761_4_lut (.I0(n69543), .I1(n68934), .I2(n45_adj_5229), 
            .I3(n68315), .O(n68936));   // verilog/uart_rx.v(119[33:55])
    defparam i52761_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48040_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n64205));
    defparam i48040_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8695[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8721[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5320));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5321));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5322));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51253_4_lut (.I0(n23_adj_5320), .I1(n21_adj_5309), .I2(n19_adj_5308), 
            .I3(n17_adj_5322), .O(n67427));
    defparam i51253_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51249_4_lut (.I0(n29_adj_5297), .I1(n27_adj_5296), .I2(n25_adj_5321), 
            .I3(n67427), .O(n67423));
    defparam i51249_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53048_4_lut (.I0(n35_adj_5295), .I1(n33_adj_5294), .I2(n31_adj_5293), 
            .I3(n67423), .O(n69223));
    defparam i53048_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5323));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53227_3_lut (.I0(n16_adj_5323), .I1(baudrate[13]), .I2(n39_adj_5292), 
            .I3(GND_net), .O(n69402));   // verilog/uart_rx.v(119[33:55])
    defparam i53227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53228_3_lut (.I0(n69402), .I1(baudrate[14]), .I2(n41_adj_5291), 
            .I3(GND_net), .O(n69403));   // verilog/uart_rx.v(119[33:55])
    defparam i53228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52109_4_lut (.I0(n41_adj_5291), .I1(n39_adj_5292), .I2(n27_adj_5296), 
            .I3(n67425), .O(n68283));
    defparam i52109_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52762_3_lut (.I0(n22_adj_5270), .I1(baudrate[7]), .I2(n27_adj_5296), 
            .I3(GND_net), .O(n68937));   // verilog/uart_rx.v(119[33:55])
    defparam i52762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53095_3_lut (.I0(n69403), .I1(baudrate[15]), .I2(n43_adj_5290), 
            .I3(GND_net), .O(n69270));   // verilog/uart_rx.v(119[33:55])
    defparam i53095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5269), .I1(baudrate[9]), 
            .I2(n31_adj_5293), .I3(GND_net), .O(n28_adj_5324));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n63786));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53551_4_lut (.I0(n28_adj_5324), .I1(n18_adj_5268), .I2(n31_adj_5293), 
            .I3(n67418), .O(n69726));   // verilog/uart_rx.v(119[33:55])
    defparam i53551_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53552_3_lut (.I0(n69726), .I1(baudrate[10]), .I2(n33_adj_5294), 
            .I3(GND_net), .O(n69727));   // verilog/uart_rx.v(119[33:55])
    defparam i53552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53425_3_lut (.I0(n69727), .I1(baudrate[11]), .I2(n35_adj_5295), 
            .I3(GND_net), .O(n69600));   // verilog/uart_rx.v(119[33:55])
    defparam i53425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52113_4_lut (.I0(n41_adj_5291), .I1(n39_adj_5292), .I2(n37_adj_5289), 
            .I3(n69223), .O(n68287));
    defparam i52113_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53225_4_lut (.I0(n69270), .I1(n68937), .I2(n43_adj_5290), 
            .I3(n68283), .O(n69400));   // verilog/uart_rx.v(119[33:55])
    defparam i53225_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53372_3_lut (.I0(n69600), .I1(baudrate[12]), .I2(n37_adj_5289), 
            .I3(GND_net), .O(n69547));   // verilog/uart_rx.v(119[33:55])
    defparam i53372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53920_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n64264), .I3(n48_adj_5276), .O(n294[19]));
    defparam i53920_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i53571_4_lut (.I0(n69547), .I1(n69400), .I2(n43_adj_5290), 
            .I3(n68287), .O(n69746));   // verilog/uart_rx.v(119[33:55])
    defparam i53571_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53572_3_lut (.I0(n69746), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n69747));   // verilog/uart_rx.v(119[33:55])
    defparam i53572_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8565[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1050 (.I0(n64246), .I1(n48_adj_5325), .I2(n8539[14]), 
            .I3(GND_net), .O(n1702));
    defparam i1_3_lut_adj_1050.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8565[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8461[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8487[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8513[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8539[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8565[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8565[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5326));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5327));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1051 (.I0(n26078), .I1(n48_adj_5328), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1051.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8565[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5329));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8487[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8513[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8539[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8565[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5330));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(n62382), .I1(n48_adj_5263), .I2(GND_net), 
            .I3(GND_net), .O(n1560));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8539[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5262), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8461[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5331));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5332));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5248), .I1(baudrate[4]), 
            .I2(n41_adj_5331), .I3(GND_net), .O(n40_adj_5333));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53442_4_lut (.I0(n40_adj_5333), .I1(n36_adj_5332), .I2(n41_adj_5331), 
            .I3(n67634), .O(n69617));   // verilog/uart_rx.v(119[33:55])
    defparam i53442_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53443_3_lut (.I0(n69617), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n69618));   // verilog/uart_rx.v(119[33:55])
    defparam i53443_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53340_3_lut (.I0(n69618), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n69515));   // verilog/uart_rx.v(119[33:55])
    defparam i53340_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52177_3_lut (.I0(n69515), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i52177_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(n62380), .I1(n48), .I2(GND_net), .I3(GND_net), 
            .O(n1415));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8513[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1054 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62800));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1054.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1055 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62816));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1055.LUT_INIT = 16'hfffb;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8539[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8565[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63776));
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n63960));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63962));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n63850));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n63810));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n63852), .I1(n63810), .I2(n63850), 
            .I3(n63846), .O(n63832));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1062 (.I0(n63960), .I1(n63786), .I2(n63844), 
            .I3(n63776), .O(n26081));
    defparam i1_4_lut_adj_1062.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n63760));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n63758));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1065 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62736));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1065.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1066 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62768));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1066.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n63380));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n63844));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n63846));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63798));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n63802));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n63408));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1073 (.I0(n63408), .I1(n63858), .I2(n63802), 
            .I3(n63798), .O(n26055));
    defparam i1_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1074 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62752));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1074.LUT_INIT = 16'hffef;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n67032), .I1(baudrate[2]), 
            .I2(n69910), .I3(n48_adj_5258), .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46), .I1(baudrate[3]), .I2(n59901), 
            .I3(GND_net), .O(n48_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n63380), .I1(n63758), .I2(n63760), 
            .I3(n63756), .O(n63392));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1076 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n62784));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1076.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1077 (.I0(n63392), .I1(n26055), .I2(n63384), 
            .I3(n63860), .O(n26011));
    defparam i1_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1078 (.I0(n26011), .I1(n48_adj_5260), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1078.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i29785_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n60200));   // verilog/uart_rx.v(119[33:55])
    defparam i29785_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n60200), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5334));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53042_3_lut (.I0(n42_adj_5334), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n69217));   // verilog/uart_rx.v(119[33:55])
    defparam i53042_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53043_3_lut (.I0(n69217), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n69218));   // verilog/uart_rx.v(119[33:55])
    defparam i53043_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n69218), .I1(baudrate[5]), 
            .I2(n59907), .I3(GND_net), .O(n48_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(n63768), .I1(n26081), .I2(n63832), 
            .I3(n63766), .O(n26014));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1080 (.I0(n26014), .I1(n48_adj_5267), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1080.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8461[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8487[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8513[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8539[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8539[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8539[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5335));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8539[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5336));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(n63844), .I1(n63800), .I2(n63802), 
            .I3(baudrate[11]), .O(n63830));
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1082 (.I0(n63830), .I1(n63832), .I2(n63820), 
            .I3(n63754), .O(n26078));
    defparam i1_4_lut_adj_1082.LUT_INIT = 16'hfffe;
    SB_LUT4 i29808_rep_5_2_lut (.I0(n8539[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n60183));   // verilog/uart_rx.v(119[33:55])
    defparam i29808_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n60183), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5337));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53032_3_lut (.I0(n32_adj_5337), .I1(baudrate[6]), .I2(n39_adj_5230), 
            .I3(GND_net), .O(n69207));   // verilog/uart_rx.v(119[33:55])
    defparam i53032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53033_3_lut (.I0(n69207), .I1(baudrate[7]), .I2(n41_adj_5231), 
            .I3(GND_net), .O(n69208));   // verilog/uart_rx.v(119[33:55])
    defparam i53033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52324_4_lut (.I0(n41_adj_5231), .I1(n39_adj_5230), .I2(n37_adj_5336), 
            .I3(n67603), .O(n68498));
    defparam i52324_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53066_3_lut (.I0(n34_adj_5247), .I1(baudrate[5]), .I2(n37_adj_5336), 
            .I3(GND_net), .O(n69241));   // verilog/uart_rx.v(119[33:55])
    defparam i53066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52192_3_lut (.I0(n69208), .I1(baudrate[8]), .I2(n43_adj_5335), 
            .I3(GND_net), .O(n68366));   // verilog/uart_rx.v(119[33:55])
    defparam i52192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53333_4_lut (.I0(n68366), .I1(n69241), .I2(n43_adj_5335), 
            .I3(n68498), .O(n69508));   // verilog/uart_rx.v(119[33:55])
    defparam i53333_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53334_3_lut (.I0(n69508), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n69509));   // verilog/uart_rx.v(119[33:55])
    defparam i53334_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n69509), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5328));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8461[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8487[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8513[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8513[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8513[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5338));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1083 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n62368));
    defparam i1_3_lut_4_lut_adj_1083.LUT_INIT = 16'hfffe;
    SB_LUT4 i48063_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n64228));
    defparam i48063_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53034_3_lut (.I0(n32_adj_5264), .I1(baudrate[5]), .I2(n39_adj_5232), 
            .I3(GND_net), .O(n69209));   // verilog/uart_rx.v(119[33:55])
    defparam i53034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53035_3_lut (.I0(n69209), .I1(baudrate[6]), .I2(n41_adj_5233), 
            .I3(GND_net), .O(n69210));   // verilog/uart_rx.v(119[33:55])
    defparam i53035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52334_4_lut (.I0(n41_adj_5233), .I1(n39_adj_5232), .I2(n37_adj_5234), 
            .I3(n67614), .O(n68508));
    defparam i52334_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53064_3_lut (.I0(n34_adj_5246), .I1(baudrate[4]), .I2(n37_adj_5234), 
            .I3(GND_net), .O(n69239));   // verilog/uart_rx.v(119[33:55])
    defparam i53064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52185_3_lut (.I0(n69210), .I1(baudrate[7]), .I2(n43_adj_5338), 
            .I3(GND_net), .O(n68359));   // verilog/uart_rx.v(119[33:55])
    defparam i52185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53335_4_lut (.I0(n68359), .I1(n69239), .I2(n43_adj_5338), 
            .I3(n68508), .O(n69510));   // verilog/uart_rx.v(119[33:55])
    defparam i53335_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53336_3_lut (.I0(n69510), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n69511));   // verilog/uart_rx.v(119[33:55])
    defparam i53336_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n69511), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5325));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5816_2_lut (.I0(n21444), .I1(n11848), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_5339));   // verilog/uart_rx.v(119[33:55])
    defparam i5816_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5339), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5340));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5341));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5245), .I1(baudrate[4]), 
            .I2(n43_adj_5340), .I3(GND_net), .O(n42_adj_5342));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53438_4_lut (.I0(n42_adj_5342), .I1(n38_adj_5341), .I2(n43_adj_5340), 
            .I3(n67641), .O(n69613));   // verilog/uart_rx.v(119[33:55])
    defparam i53438_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53439_3_lut (.I0(n69613), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n69614));   // verilog/uart_rx.v(119[33:55])
    defparam i53439_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n62890));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5343));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53046_3_lut (.I0(n42_adj_5343), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n69221));   // verilog/uart_rx.v(119[33:55])
    defparam i53046_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53047_3_lut (.I0(n69221), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n69222));   // verilog/uart_rx.v(119[33:55])
    defparam i53047_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n69222), .I1(baudrate[4]), 
            .I2(n59905), .I3(GND_net), .O(n48_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_2_lut_3_lut_adj_1085 (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[2] ), .I3(GND_net), .O(n4));
    defparam i1_2_lut_3_lut_adj_1085.LUT_INIT = 16'hfdfd;
    SB_LUT4 i51822_4_lut (.I0(n25994), .I1(n67321), .I2(n48_adj_5258), 
            .I3(baudrate[0]), .O(n804));
    defparam i51822_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i7341_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21444));   // verilog/uart_rx.v(119[33:55])
    defparam i7341_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5261), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n62698));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'h0100;
    SB_LUT4 i48057_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n64222));
    defparam i48057_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(n59955), .I1(n62698), .I2(n63958), 
            .I3(baudrate[16]), .O(n62726));
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'h0004;
    SB_LUT4 i48127_4_lut (.I0(n64222), .I1(n64151), .I2(n64155), .I3(n64064), 
            .O(n64292));
    defparam i48127_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53735_4_lut (.I0(n64282), .I1(n67315), .I2(n64292), .I3(n62726), 
            .O(n69910));
    defparam i53735_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i535_4_lut (.I0(n69910), .I1(n44_adj_5259), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 i47986_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n64151));
    defparam i47986_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5257), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_3_lut_4_lut_adj_1088 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n62370));
    defparam i1_3_lut_4_lut_adj_1088.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7342_4_lut (.I0(n960), .I1(n11848), .I2(n21444), .I3(baudrate[3]), 
            .O(n21446));   // verilog/uart_rx.v(119[33:55])
    defparam i7342_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8877[20]), .I3(n294[1]), .O(n41_adj_5344));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8877[19]), .I3(n294[1]), .O(n39_adj_5345));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8877[14]), .I3(n294[1]), .O(n29_adj_5346));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8877[15]), .I3(n294[1]), .O(n31_adj_5347));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8877[11]), .I3(n294[1]), .O(n23_adj_5348));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8877[12]), .I3(n294[1]), .O(n25_adj_5349));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8877[16]), .I3(n294[1]), .O(n33_adj_5350));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5256), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8461[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8877[17]), .I3(n294[1]), .O(n35_adj_5351));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8877[18]), .I3(n294[1]), .O(n37_adj_5352));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8877[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8877[22]), .I3(n294[1]), .O(n45_adj_5353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8487[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8877[21]), .I3(n294[1]), .O(n43_adj_5354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8877[5]), .I3(n294[1]), .O(n11_adj_5355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8877[6]), .I3(n294[1]), .O(n13_adj_5356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8877[7]), .I3(n294[1]), .O(n15_adj_5357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_adj_1089 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n63852));
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8877[13]), .I3(n294[1]), .O(n27_adj_5358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8877[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n63754));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n63756));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8877[8]), .I3(n294[1]), .O(n17_adj_5359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8877[9]), .I3(n294[1]), .O(n19_adj_5360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8877[10]), .I3(n294[1]), .O(n21_adj_5361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i51811_4_lut (.I0(n27_adj_5358), .I1(n15_adj_5357), .I2(n13_adj_5356), 
            .I3(n11_adj_5355), .O(n67985));
    defparam i51811_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i43829_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n59955));
    defparam i43829_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i54478_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n26049), .I3(n48_adj_5274), .O(n294[8]));
    defparam i54478_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51829_4_lut (.I0(n21_adj_5361), .I1(n19_adj_5360), .I2(n17_adj_5359), 
            .I3(n9), .O(n68003));
    defparam i51829_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5354), .I3(GND_net), .O(n16_adj_5362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51756_2_lut (.I0(n43_adj_5354), .I1(n19_adj_5360), .I2(GND_net), 
            .I3(GND_net), .O(n67930));
    defparam i51756_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5359), .I3(GND_net), .O(n8_adj_5363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5362), .I1(baudrate[22]), 
            .I2(n45_adj_5353), .I3(GND_net), .O(n24_adj_5364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8877[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51844_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n68018));
    defparam i51844_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i48006_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n64171));
    defparam i48006_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i52605_4_lut (.I0(n13_adj_5356), .I1(n11_adj_5355), .I2(n9), 
            .I3(n68018), .O(n68780));
    defparam i52605_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52601_4_lut (.I0(n19_adj_5360), .I1(n17_adj_5359), .I2(n15_adj_5357), 
            .I3(n68780), .O(n68776));
    defparam i52601_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48117_4_lut (.I0(n64171), .I1(n63384), .I2(n63756), .I3(baudrate[9]), 
            .O(n64282));
    defparam i48117_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53498_4_lut (.I0(n25_adj_5349), .I1(n23_adj_5348), .I2(n21_adj_5361), 
            .I3(n68776), .O(n69673));
    defparam i53498_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52938_4_lut (.I0(n31_adj_5347), .I1(n29_adj_5346), .I2(n27_adj_5358), 
            .I3(n69673), .O(n69113));
    defparam i52938_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53577_4_lut (.I0(n37_adj_5352), .I1(n35_adj_5351), .I2(n33_adj_5350), 
            .I3(n69113), .O(n69752));
    defparam i53577_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5350), .I3(GND_net), .O(n12_adj_5365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n62402), .I3(n48_adj_5366), .O(n4_adj_5367));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_4_lut_adj_1092 (.I0(baudrate[17]), .I1(n64187), .I2(baudrate[2]), 
            .I3(n44071), .O(n62318));
    defparam i1_4_lut_adj_1092.LUT_INIT = 16'h0100;
    SB_LUT4 i52984_3_lut (.I0(n4_adj_5367), .I1(baudrate[13]), .I2(n27_adj_5358), 
            .I3(GND_net), .O(n69159));   // verilog/uart_rx.v(119[33:55])
    defparam i52984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52985_3_lut (.I0(n69159), .I1(baudrate[14]), .I2(n29_adj_5346), 
            .I3(GND_net), .O(n69160));   // verilog/uart_rx.v(119[33:55])
    defparam i52985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47822_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n26049), .I3(baudrate[15]), .O(n63984));
    defparam i47822_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1093 (.I0(n64236), .I1(n62318), .I2(n26049), 
            .I3(n64151), .O(n61397));
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'h0004;
    SB_LUT4 i51803_2_lut (.I0(n33_adj_5350), .I1(n15_adj_5357), .I2(GND_net), 
            .I3(GND_net), .O(n67977));
    defparam i51803_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5356), .I3(GND_net), .O(n10_adj_5368));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5365), .I1(baudrate[17]), 
            .I2(n35_adj_5351), .I3(GND_net), .O(n30_adj_5369));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1094 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n44073), .O(n62642));
    defparam i1_4_lut_adj_1094.LUT_INIT = 16'h0100;
    SB_LUT4 i51805_4_lut (.I0(n33_adj_5350), .I1(n31_adj_5347), .I2(n29_adj_5346), 
            .I3(n67985), .O(n67979));
    defparam i51805_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53460_4_lut (.I0(n30_adj_5369), .I1(n10_adj_5368), .I2(n35_adj_5351), 
            .I3(n67977), .O(n69635));   // verilog/uart_rx.v(119[33:55])
    defparam i53460_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1095 (.I0(n62642), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n62660));
    defparam i1_4_lut_adj_1095.LUT_INIT = 16'h0002;
    SB_LUT4 i52241_3_lut (.I0(n69160), .I1(baudrate[15]), .I2(n31_adj_5347), 
            .I3(GND_net), .O(n68415));   // verilog/uart_rx.v(119[33:55])
    defparam i52241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53650_4_lut (.I0(n68415), .I1(n69635), .I2(n35_adj_5351), 
            .I3(n67979), .O(n69825));   // verilog/uart_rx.v(119[33:55])
    defparam i53650_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53651_3_lut (.I0(n69825), .I1(baudrate[18]), .I2(n37_adj_5352), 
            .I3(GND_net), .O(n69826));   // verilog/uart_rx.v(119[33:55])
    defparam i53651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5370));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48129_4_lut (.I0(n64228), .I1(n64151), .I2(n64155), .I3(n64064), 
            .O(n64294));
    defparam i48129_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52994_3_lut (.I0(n6_adj_5370), .I1(baudrate[10]), .I2(n21_adj_5361), 
            .I3(GND_net), .O(n69169));   // verilog/uart_rx.v(119[33:55])
    defparam i52994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(n64282), .I1(n64294), .I2(n59955), 
            .I3(n62660), .O(n60673));
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(n62884), .I1(n62880), .I2(n62882), 
            .I3(n64064), .O(n62902));
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'hfffe;
    SB_LUT4 i47821_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n26049), .I3(GND_net), .O(n60167));
    defparam i47821_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_1098 (.I0(n64187), .I1(n62888), .I2(n62890), 
            .I3(n62886), .O(n62904));
    defparam i1_4_lut_adj_1098.LUT_INIT = 16'hfffe;
    SB_LUT4 i52995_3_lut (.I0(n69169), .I1(baudrate[11]), .I2(n23_adj_5348), 
            .I3(GND_net), .O(n69170));   // verilog/uart_rx.v(119[33:55])
    defparam i52995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51784_4_lut (.I0(n43_adj_5354), .I1(n25_adj_5349), .I2(n23_adj_5348), 
            .I3(n68003), .O(n67958));
    defparam i51784_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53135_4_lut (.I0(n24_adj_5364), .I1(n8_adj_5363), .I2(n45_adj_5353), 
            .I3(n67930), .O(n69310));   // verilog/uart_rx.v(119[33:55])
    defparam i53135_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52239_3_lut (.I0(n69170), .I1(baudrate[12]), .I2(n25_adj_5349), 
            .I3(GND_net), .O(n68413));   // verilog/uart_rx.v(119[33:55])
    defparam i52239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1099 (.I0(n62904), .I1(n26052), .I2(n62902), 
            .I3(GND_net), .O(n25994));
    defparam i1_3_lut_adj_1099.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n60673), .I1(baudrate[2]), 
            .I2(n61397), .I3(GND_net), .O(n48_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53594_3_lut (.I0(n69826), .I1(baudrate[19]), .I2(n39_adj_5345), 
            .I3(GND_net), .O(n69769));   // verilog/uart_rx.v(119[33:55])
    defparam i53594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51786_4_lut (.I0(n43_adj_5354), .I1(n41_adj_5344), .I2(n39_adj_5345), 
            .I3(n69752), .O(n67960));
    defparam i51786_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47816_2_lut (.I0(baudrate[17]), .I1(n26049), .I2(GND_net), 
            .I3(GND_net), .O(n63978));
    defparam i47816_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53535_4_lut (.I0(n68413), .I1(n69310), .I2(n45_adj_5353), 
            .I3(n67958), .O(n69710));   // verilog/uart_rx.v(119[33:55])
    defparam i53535_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52247_3_lut (.I0(n69769), .I1(baudrate[20]), .I2(n41_adj_5344), 
            .I3(GND_net), .O(n68421));   // verilog/uart_rx.v(119[33:55])
    defparam i52247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54507_2_lut (.I0(n48_adj_5258), .I1(n25994), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i54507_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i53968_2_lut (.I0(n48_adj_5260), .I1(n26011), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i53968_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1100 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n62330));
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8877[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53537_4_lut (.I0(n68421), .I1(n69710), .I2(n45_adj_5353), 
            .I3(n67960), .O(n69712));   // verilog/uart_rx.v(119[33:55])
    defparam i53537_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1101 (.I0(n63958), .I1(n63802), .I2(n62330), 
            .I3(n63800), .O(n62338));
    defparam i1_4_lut_adj_1101.LUT_INIT = 16'hfffe;
    SB_LUT4 i54232_4_lut (.I0(n62338), .I1(n69712), .I2(baudrate[23]), 
            .I3(n3253), .O(n61327));   // verilog/uart_rx.v(119[33:55])
    defparam i54232_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 i1_4_lut_adj_1102 (.I0(n63766), .I1(n63852), .I2(baudrate[16]), 
            .I3(n44071), .O(n62968));
    defparam i1_4_lut_adj_1102.LUT_INIT = 16'h0100;
    SB_LUT4 i51883_3_lut (.I0(n60673), .I1(n61397), .I2(baudrate[2]), 
            .I3(GND_net), .O(n66965));   // verilog/uart_rx.v(119[33:55])
    defparam i51883_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i51688_4_lut (.I0(n59955), .I1(n62968), .I2(n63768), .I3(n63380), 
            .O(n66966));   // verilog/uart_rx.v(119[33:55])
    defparam i51688_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n66966), .I1(n66965), .I2(n294[21]), 
            .I3(n63978), .O(n59901));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 div_37_i534_3_lut (.I0(n59901), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n59905));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53974_2_lut (.I0(n48_adj_5267), .I1(n26014), .I2(GND_net), 
            .I3(GND_net), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i53974_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i7334_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21434));   // verilog/uart_rx.v(119[33:55])
    defparam i7334_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i47990_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n64155));
    defparam i47990_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5659_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n11684), .I3(n21436), 
            .O(n46_adj_5371));   // verilog/uart_rx.v(119[33:55])
    defparam i5659_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i639_4_lut (.I0(n59905), .I1(n294[19]), .I2(n46_adj_5371), 
            .I3(baudrate[4]), .O(n59907));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51193_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n67367));
    defparam i51193_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8851[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8851[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51171_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n67345));
    defparam i51171_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8851[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5372));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8851[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5373));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8851[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5830_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n11855), .I3(n21446), 
            .O(n46_adj_5374));   // verilog/uart_rx.v(119[33:55])
    defparam i5830_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5375));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i742_4_lut (.I0(n59907), .I1(n294[18]), .I2(n46_adj_5374), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 i1_2_lut_4_lut_adj_1103 (.I0(n69300), .I1(baudrate[21]), .I2(n3046), 
            .I3(n62400), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1103.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8851[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5376));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8851[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54499_2_lut_4_lut (.I0(n69300), .I1(baudrate[21]), .I2(n3046), 
            .I3(n26081), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i54499_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8461[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8487[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8851[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5377));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5378));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5379));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51158_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n67332));
    defparam i51158_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8851[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8851[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5380));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51128_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n67302));
    defparam i51128_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5381));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8851[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8851[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53036_3_lut (.I0(n34_adj_5255), .I1(baudrate[5]), .I2(n41_adj_5235), 
            .I3(GND_net), .O(n69211));   // verilog/uart_rx.v(119[33:55])
    defparam i53036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53037_3_lut (.I0(n69211), .I1(baudrate[6]), .I2(n43_adj_5236), 
            .I3(GND_net), .O(n69212));   // verilog/uart_rx.v(119[33:55])
    defparam i53037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5382));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8851[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52342_4_lut (.I0(n43_adj_5236), .I1(n41_adj_5235), .I2(n39_adj_5237), 
            .I3(n67626), .O(n68516));
    defparam i52342_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8851[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5383));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5384));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5244), .I1(baudrate[4]), 
            .I2(n39_adj_5237), .I3(GND_net), .O(n38_adj_5385));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8851[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8851[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52183_3_lut (.I0(n69212), .I1(baudrate[7]), .I2(n45_adj_5377), 
            .I3(GND_net), .O(n68357));   // verilog/uart_rx.v(119[33:55])
    defparam i52183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8851[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53062_4_lut (.I0(n68357), .I1(n38_adj_5385), .I2(n45_adj_5377), 
            .I3(n68516), .O(n69237));   // verilog/uart_rx.v(119[33:55])
    defparam i53062_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8851[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5386));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5387));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53063_3_lut (.I0(n69237), .I1(baudrate[8]), .I2(n1408), .I3(GND_net), 
            .O(n48_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam i53063_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5388));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5389));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n63800));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63958));
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'heeee;
    SB_LUT4 i51084_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n67258));
    defparam i51084_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1106 (.I0(n63962), .I1(n63964), .I2(n63800), 
            .I3(n63960), .O(n26061));
    defparam i1_4_lut_adj_1106.LUT_INIT = 16'hfffe;
    SB_LUT4 i50974_4_lut (.I0(n29_adj_5389), .I1(n17_adj_5388), .I2(n15_adj_5387), 
            .I3(n13_adj_5386), .O(n67148));
    defparam i50974_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8487[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51905_4_lut (.I0(n11_adj_5383), .I1(n9_adj_5382), .I2(n3171), 
            .I3(baudrate[2]), .O(n68079));
    defparam i51905_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i52641_4_lut (.I0(n17_adj_5388), .I1(n15_adj_5387), .I2(n13_adj_5386), 
            .I3(n68079), .O(n68816));
    defparam i52641_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52639_4_lut (.I0(n23_adj_5381), .I1(n21_adj_5380), .I2(n19_adj_5384), 
            .I3(n68816), .O(n68814));
    defparam i52639_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8513[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50976_4_lut (.I0(n29_adj_5389), .I1(n27_adj_5379), .I2(n25_adj_5378), 
            .I3(n68814), .O(n67150));
    defparam i50976_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5390));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8539[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8565[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53197_3_lut (.I0(n6_adj_5390), .I1(baudrate[13]), .I2(n29_adj_5389), 
            .I3(GND_net), .O(n69372));   // verilog/uart_rx.v(119[33:55])
    defparam i53197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8565[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5391));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5253), .I1(baudrate[17]), 
            .I2(n37_adj_5375), .I3(GND_net), .O(n32_adj_5392));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53198_3_lut (.I0(n69372), .I1(baudrate[14]), .I2(n31_adj_5373), 
            .I3(GND_net), .O(n69373));   // verilog/uart_rx.v(119[33:55])
    defparam i53198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51881_4_lut (.I0(n35_adj_5376), .I1(n33_adj_5372), .I2(n31_adj_5373), 
            .I3(n67148), .O(n68055));
    defparam i51881_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53452_4_lut (.I0(n32_adj_5392), .I1(n12_adj_5252), .I2(n37_adj_5375), 
            .I3(n68050), .O(n69627));   // verilog/uart_rx.v(119[33:55])
    defparam i53452_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53134_3_lut (.I0(n69373), .I1(baudrate[15]), .I2(n33_adj_5372), 
            .I3(GND_net), .O(n30_adj_5393));   // verilog/uart_rx.v(119[33:55])
    defparam i53134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5394));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53199_3_lut (.I0(n8_adj_5251), .I1(baudrate[10]), .I2(n23_adj_5381), 
            .I3(GND_net), .O(n69374));   // verilog/uart_rx.v(119[33:55])
    defparam i53199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5395));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53200_3_lut (.I0(n69374), .I1(baudrate[11]), .I2(n25_adj_5378), 
            .I3(GND_net), .O(n69375));   // verilog/uart_rx.v(119[33:55])
    defparam i53200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51893_4_lut (.I0(n25_adj_5378), .I1(n23_adj_5381), .I2(n21_adj_5380), 
            .I3(n67158), .O(n68067));
    defparam i51893_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53131_3_lut (.I0(n10_adj_5254), .I1(baudrate[9]), .I2(n21_adj_5380), 
            .I3(GND_net), .O(n69306));   // verilog/uart_rx.v(119[33:55])
    defparam i53131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8565[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53130_3_lut (.I0(n69375), .I1(baudrate[12]), .I2(n27_adj_5379), 
            .I3(GND_net), .O(n24_adj_5396));   // verilog/uart_rx.v(119[33:55])
    defparam i53130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52956_4_lut (.I0(n35_adj_5376), .I1(n33_adj_5372), .I2(n31_adj_5373), 
            .I3(n67150), .O(n69131));
    defparam i52956_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51412_4_lut (.I0(n35_adj_5395), .I1(n33_adj_5394), .I2(n31_adj_5391), 
            .I3(n29_adj_5397), .O(n67586));
    defparam i51412_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32), .I1(baudrate[9]), 
            .I2(n43_adj_5329), .I3(GND_net), .O(n40_adj_5398));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5399));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53026_3_lut (.I0(n28_adj_5399), .I1(baudrate[5]), .I2(n35_adj_5395), 
            .I3(GND_net), .O(n69201));   // verilog/uart_rx.v(119[33:55])
    defparam i53026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53027_3_lut (.I0(n69201), .I1(baudrate[6]), .I2(n37_adj_5326), 
            .I3(GND_net), .O(n69202));   // verilog/uart_rx.v(119[33:55])
    defparam i53027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51408_4_lut (.I0(n41_adj_5330), .I1(n39_adj_5327), .I2(n37_adj_5326), 
            .I3(n67586), .O(n67582));
    defparam i51408_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53432_4_lut (.I0(n40_adj_5398), .I1(n30), .I2(n43_adj_5329), 
            .I3(n67580), .O(n69607));   // verilog/uart_rx.v(119[33:55])
    defparam i53432_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53646_4_lut (.I0(n30_adj_5393), .I1(n69627), .I2(n37_adj_5375), 
            .I3(n68055), .O(n69821));   // verilog/uart_rx.v(119[33:55])
    defparam i53646_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53317_4_lut (.I0(n24_adj_5396), .I1(n69306), .I2(n27_adj_5379), 
            .I3(n68067), .O(n69492));   // verilog/uart_rx.v(119[33:55])
    defparam i53317_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53716_4_lut (.I0(n69492), .I1(n69821), .I2(n37_adj_5375), 
            .I3(n69131), .O(n69891));   // verilog/uart_rx.v(119[33:55])
    defparam i53716_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52199_3_lut (.I0(n69202), .I1(baudrate[7]), .I2(n39_adj_5327), 
            .I3(GND_net), .O(n68373));   // verilog/uart_rx.v(119[33:55])
    defparam i52199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53717_3_lut (.I0(n69891), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n69892));   // verilog/uart_rx.v(119[33:55])
    defparam i53717_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53707_3_lut (.I0(n69892), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n69882));   // verilog/uart_rx.v(119[33:55])
    defparam i53707_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53640_4_lut (.I0(n68373), .I1(n69607), .I2(n43_adj_5329), 
            .I3(n67582), .O(n69815));   // verilog/uart_rx.v(119[33:55])
    defparam i53640_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53641_3_lut (.I0(n69815), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n69816));   // verilog/uart_rx.v(119[33:55])
    defparam i53641_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53608_3_lut (.I0(n69816), .I1(baudrate[11]), .I2(n1831), 
            .I3(GND_net), .O(n48_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam i53608_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53526_3_lut (.I0(n69882), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n69701));   // verilog/uart_rx.v(119[33:55])
    defparam i53526_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n62384), .I1(n48_adj_5277), .I2(GND_net), 
            .I3(GND_net), .O(n1977));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h2222;
    SB_LUT4 i53527_3_lut (.I0(n69701), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n69702));   // verilog/uart_rx.v(119[33:55])
    defparam i53527_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52237_3_lut (.I0(n69702), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5366));   // verilog/uart_rx.v(119[33:55])
    defparam i52237_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51064_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n67238));
    defparam i51064_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51008_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n67182));
    defparam i51008_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51029_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n67203));
    defparam i51029_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8851[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8851[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (enable_slow_N_4340, ready_prev, clk16MHz, n6195, \state[2] , 
            GND_net, n30024, rw, n58524, data_ready, n30015, ID, 
            \state[0] , \state[1] , n58352, n30804, n30803, n30802, 
            n30801, n30800, n30799, n30798, n30797, baudrate, n30796, 
            n30795, n30794, n30793, n30792, n30791, n30790, n30772, 
            n30771, n30770, n30769, n30768, n30767, n30766, n30765, 
            n3, n6878, n11, \state[2]_adj_5 , \state[3] , n6, \state_7__N_4253[3] , 
            \state_7__N_4045[0] , \state[1]_adj_6 , \state[0]_adj_7 , 
            n59067, n61238, n59065, n5, n25956, data, n4, n49984, 
            n62253, VCC_net, sda_enable, sda_out, scl_enable, n62, 
            \state_7__N_4237[0] , \saved_addr[0] , n30054, n30049, n30047, 
            n30042, n30041, n11_adj_8, n30841, n8, n29813, n10, 
            n4_adj_9, n44006, n25984, scl) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output enable_slow_N_4340;
    output ready_prev;
    input clk16MHz;
    output [0:0]n6195;
    output \state[2] ;
    input GND_net;
    input n30024;
    output rw;
    input n58524;
    output data_ready;
    input n30015;
    output [7:0]ID;
    output \state[0] ;
    output \state[1] ;
    input n58352;
    input n30804;
    input n30803;
    input n30802;
    input n30801;
    input n30800;
    input n30799;
    input n30798;
    input n30797;
    output [31:0]baudrate;
    input n30796;
    input n30795;
    input n30794;
    input n30793;
    input n30792;
    input n30791;
    input n30790;
    input n30772;
    input n30771;
    input n30770;
    input n30769;
    input n30768;
    input n30767;
    input n30766;
    input n30765;
    output n3;
    output n6878;
    output n11;
    output \state[2]_adj_5 ;
    output \state[3] ;
    output n6;
    input \state_7__N_4253[3] ;
    input \state_7__N_4045[0] ;
    output \state[1]_adj_6 ;
    output \state[0]_adj_7 ;
    output n59067;
    output n61238;
    output n59065;
    output n5;
    output n25956;
    output [7:0]data;
    output n4;
    output n49984;
    output n62253;
    input VCC_net;
    output sda_enable;
    output sda_out;
    output scl_enable;
    input n62;
    output \state_7__N_4237[0] ;
    output \saved_addr[0] ;
    input n30054;
    input n30049;
    input n30047;
    input n30042;
    input n30041;
    output n11_adj_8;
    input n30841;
    input n8;
    input n29813;
    output n10;
    output n4_adj_9;
    output n44006;
    output n25984;
    output scl;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire enable;
    wire [15:0]delay_counter_15__N_4083;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    wire [15:0]n5403;
    
    wire n51537, n51536, n51535, n51534, n51533, n7100, n51532, 
        n50082, n7099, n51531, n7098, n51530, n7097, n51529, n7096, 
        n51528, n51527, n7094, n51526, n51525, n51524, n51523, 
        n28101, n50099;
    wire [2:0]n17;
    
    wire n28171;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n29526, n54052, n59008, n58344, data_ready_N_4155, n30789, 
        n30788, n30787, n30786, n30785, n30784, n30783, n30782, 
        n30781, n30780, n30779, n30778, n30777, n30776, n30775, 
        n30774, n59009, n59068, n25838;
    wire [7:0]state_7__N_4012;
    
    wire n61958, n14, n13, n14_adj_5114, n15, n9, n65, n10_c, 
        n44000, n49980, n15_adj_5116, n67026, n44045, n28163, n43931, 
        n4_c, n58508, n48, n30053, n4_adj_5120, n67134;
    
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4340));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n6195[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1121_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5403[5]), 
            .I3(n51537), .O(delay_counter_15__N_4083[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1121_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5403[5]), 
            .I3(n51536), .O(delay_counter_15__N_4083[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_16 (.CI(n51536), .I0(delay_counter[14]), .I1(n5403[5]), 
            .CO(n51537));
    SB_LUT4 add_1121_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5403[5]), 
            .I3(n51535), .O(delay_counter_15__N_4083[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_15 (.CI(n51535), .I0(delay_counter[13]), .I1(n5403[5]), 
            .CO(n51536));
    SB_LUT4 add_1121_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5403[5]), 
            .I3(n51534), .O(delay_counter_15__N_4083[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_14 (.CI(n51534), .I0(delay_counter[12]), .I1(n5403[5]), 
            .CO(n51535));
    SB_LUT4 add_1121_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5403[5]), 
            .I3(n51533), .O(delay_counter_15__N_4083[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_13 (.CI(n51533), .I0(delay_counter[11]), .I1(n5403[5]), 
            .CO(n51534));
    SB_LUT4 add_1121_12_lut (.I0(n50082), .I1(delay_counter[10]), .I2(n5403[5]), 
            .I3(n51532), .O(n7100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_12 (.CI(n51532), .I0(delay_counter[10]), .I1(n5403[5]), 
            .CO(n51533));
    SB_LUT4 add_1121_11_lut (.I0(n50082), .I1(delay_counter[9]), .I2(n5403[5]), 
            .I3(n51531), .O(n7099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_11 (.CI(n51531), .I0(delay_counter[9]), .I1(n5403[5]), 
            .CO(n51532));
    SB_LUT4 add_1121_10_lut (.I0(n50082), .I1(delay_counter[8]), .I2(n5403[5]), 
            .I3(n51530), .O(n7098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_10 (.CI(n51530), .I0(delay_counter[8]), .I1(n5403[5]), 
            .CO(n51531));
    SB_LUT4 add_1121_9_lut (.I0(n50082), .I1(delay_counter[7]), .I2(n5403[5]), 
            .I3(n51529), .O(n7097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_9 (.CI(n51529), .I0(delay_counter[7]), .I1(n5403[5]), 
            .CO(n51530));
    SB_LUT4 add_1121_8_lut (.I0(n50082), .I1(delay_counter[6]), .I2(n5403[5]), 
            .I3(n51528), .O(n7096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_8 (.CI(n51528), .I0(delay_counter[6]), .I1(n5403[5]), 
            .CO(n51529));
    SB_LUT4 add_1121_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5403[5]), 
            .I3(n51527), .O(delay_counter_15__N_4083[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_7 (.CI(n51527), .I0(delay_counter[5]), .I1(n5403[5]), 
            .CO(n51528));
    SB_LUT4 add_1121_6_lut (.I0(n50082), .I1(delay_counter[4]), .I2(n5403[5]), 
            .I3(n51526), .O(n7094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1121_6 (.CI(n51526), .I0(delay_counter[4]), .I1(n5403[5]), 
            .CO(n51527));
    SB_LUT4 add_1121_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5403[5]), 
            .I3(n51525), .O(delay_counter_15__N_4083[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_5 (.CI(n51525), .I0(delay_counter[3]), .I1(n5403[5]), 
            .CO(n51526));
    SB_LUT4 add_1121_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5403[5]), 
            .I3(n51524), .O(delay_counter_15__N_4083[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_4 (.CI(n51524), .I0(delay_counter[2]), .I1(n5403[5]), 
            .CO(n51525));
    SB_LUT4 add_1121_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5403[5]), 
            .I3(n51523), .O(delay_counter_15__N_4083[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_3 (.CI(n51523), .I0(delay_counter[1]), .I1(n5403[5]), 
            .CO(n51524));
    SB_LUT4 add_1121_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5403[5]), 
            .I3(GND_net), .O(delay_counter_15__N_4083[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1121_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1121_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5403[5]), 
            .CO(n51523));
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28101), 
            .D(delay_counter_15__N_4083[5]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28101), 
            .D(n7096), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28101), 
            .D(n7097), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28101), 
            .D(n7098), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28101), 
            .D(n7099), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n28101), .D(n7100), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n28101), .D(delay_counter_15__N_4083[11]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n28101), .D(delay_counter_15__N_4083[12]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n28101), .D(delay_counter_15__N_4083[13]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n28101), .D(delay_counter_15__N_4083[14]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n28101), .D(delay_counter_15__N_4083[15]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n30024));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n58524));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n30015));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2055__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n28171), .D(n17[1]), .R(n29526));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2055__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n28171), .D(n17[2]), .R(n29526));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2055__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n28171), .D(n54052), .R(n29526));   // verilog/eeprom.v(68[25:39])
    SB_LUT4 i1_3_lut_4_lut (.I0(enable_slow_N_4340), .I1(ready_prev), .I2(\state[2] ), 
            .I3(n59008), .O(n58344));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf2f0;
    SB_LUT4 i53765_2_lut_3_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(GND_net), .O(data_ready_N_4155));   // verilog/eeprom.v(71[5:15])
    defparam i53765_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF state_i0 (.Q(\state[0] ), .C(clk16MHz), .D(n58352));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30804));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30803));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30802));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30801));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30800));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30798));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30797));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30796));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30795));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30794));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30793));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30792));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30791));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30790));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30789));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30788));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30786));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n30785));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n30784));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n30783));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n30782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30781));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30780));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30779));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30778));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30777));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30776));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30775));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30774));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30772));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30771));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30770));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30769));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30768));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30767));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30766));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30765));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i13_2_lut (.I0(\state[2] ), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n50082));
    defparam i13_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(n59009), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n59068));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i53783_2_lut (.I0(n25838), .I1(enable_slow_N_4340), .I2(GND_net), 
            .I3(GND_net), .O(n5403[5]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i53783_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n58344), .R(data_ready_N_4155));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n61958), .D(state_7__N_4012[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i6_4_lut (.I0(delay_counter[10]), .I1(delay_counter[6]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n14));   // verilog/eeprom.v(55[12:28])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[4]), .I1(delay_counter[2]), .I2(delay_counter[0]), 
            .I3(delay_counter[5]), .O(n13));   // verilog/eeprom.v(55[12:28])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_978 (.I0(delay_counter[1]), .I1(n13), .I2(delay_counter[13]), 
            .I3(n14), .O(n14_adj_5114));   // verilog/eeprom.v(55[12:28])
    defparam i5_4_lut_adj_978.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_979 (.I0(delay_counter[9]), .I1(delay_counter[3]), 
            .I2(delay_counter[7]), .I3(delay_counter[11]), .O(n15));   // verilog/eeprom.v(55[12:28])
    defparam i6_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(delay_counter[15]), .I2(n14_adj_5114), 
            .I3(delay_counter[14]), .O(n25838));   // verilog/eeprom.v(55[12:28])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1507_Mux_0_i3_4_lut (.I0(\state[0] ), .I1(enable_slow_N_4340), 
            .I2(\state[1] ), .I3(n25838), .O(n6195[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1507_Mux_0_i3_4_lut.LUT_INIT = 16'h0a4a;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28101), 
            .D(delay_counter_15__N_4083[1]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28101), 
            .D(delay_counter_15__N_4083[2]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28101), 
            .D(delay_counter_15__N_4083[3]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28101), 
            .D(n7094), .S(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28101), 
            .D(delay_counter_15__N_4083[0]), .R(n50099));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i53743_4_lut (.I0(n6878), .I1(n11), .I2(n9), .I3(\state[2]_adj_5 ), 
            .O(n65));
    defparam i53743_4_lut.LUT_INIT = 16'h222a;
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n25838), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[2] ), .I1(n3), .I2(\state[1] ), 
            .I3(\state[0] ), .O(state_7__N_4012[1]));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'ha5f2;
    SB_LUT4 i1_4_lut_4_lut_adj_980 (.I0(\state[2] ), .I1(n3), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n50099));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_4_lut_adj_980.LUT_INIT = 16'h0052;
    SB_LUT4 i25_4_lut_4_lut (.I0(\state[2] ), .I1(n3), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n28101));   // verilog/eeprom.v(27[11:16])
    defparam i25_4_lut_4_lut.LUT_INIT = 16'h0552;
    SB_LUT4 i1_4_lut (.I0(n10_c), .I1(n9), .I2(\state_7__N_4253[3] ), 
            .I3(n44000), .O(n49980));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut.LUT_INIT = 16'h1511;
    SB_LUT4 i5914_4_lut (.I0(n15_adj_5116), .I1(n67026), .I2(n44045), 
            .I3(\state_7__N_4253[3] ), .O(n28163));   // verilog/eeprom.v(38[3] 80[10])
    defparam i5914_4_lut.LUT_INIT = 16'h353f;
    SB_LUT4 i29637_2_lut (.I0(enable_slow_N_4340), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n43931));
    defparam i29637_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_4_lut (.I0(\state_7__N_4045[0] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n29526));   // verilog/eeprom.v(68[25:39])
    defparam i2_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_981 (.I0(\state[2] ), .I1(\state_7__N_4045[0] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n28171));
    defparam i1_4_lut_adj_981.LUT_INIT = 16'h5004;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[1]_adj_6 ), .I1(\state[2]_adj_5 ), 
            .I2(\state[0]_adj_7 ), .I3(\state[3] ), .O(n59067));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36849_2_lut_3_lut_4_lut (.I0(enable_slow_N_4340), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i36849_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(byte_counter[2]), .I1(n59009), .I2(byte_counter[0]), 
            .I3(byte_counter[1]), .O(n61238));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(byte_counter[2]), .I1(n59009), .I2(byte_counter[1]), 
            .I3(byte_counter[0]), .O(n59065));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i36856_3_lut_4_lut (.I0(n43931), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i36856_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i51052_4_lut_4_lut (.I0(\state[1]_adj_6 ), .I1(\state[2]_adj_5 ), 
            .I2(\state[0]_adj_7 ), .I3(n4_c), .O(n67026));   // verilog/eeprom.v(55[12:28])
    defparam i51052_4_lut_4_lut.LUT_INIT = 16'hffc1;
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[1]_adj_6 ), .I1(\state[2]_adj_5 ), 
            .I2(\state[0]_adj_7 ), .I3(GND_net), .O(n5));   // verilog/eeprom.v(55[12:28])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n59008));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(ready_prev), .I1(n59008), .I2(\state[2] ), .I3(n59067), 
            .O(n59009));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_adj_983 (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n25956));   // verilog/eeprom.v(38[3] 80[10])
    defparam i1_2_lut_adj_983.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut (.I0(\state_7__N_4253[3] ), .I1(data[4]), .I2(n4), 
            .I3(n49984), .O(n58508));   // verilog/i2c_controller.v(33[12:17])
    defparam i11_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35708_3_lut (.I0(n48), .I1(\state_7__N_4253[3] ), .I2(data[6]), 
            .I3(GND_net), .O(n30053));   // verilog/i2c_controller.v(33[12:17])
    defparam i35708_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i29748_3_lut_4_lut (.I0(\state[2]_adj_5 ), .I1(\state[3] ), 
            .I2(\state[0]_adj_7 ), .I3(GND_net), .O(n44045));
    defparam i29748_3_lut_4_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_984 (.I0(enable_slow_N_4340), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(GND_net), .O(n54052));
    defparam i1_2_lut_3_lut_adj_984.LUT_INIT = 16'hd2d2;
    SB_LUT4 i16375_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[7]), 
            .I3(baudrate[15]), .O(n30782));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16376_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[6]), 
            .I3(baudrate[14]), .O(n30783));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16377_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[5]), 
            .I3(baudrate[13]), .O(n30784));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16378_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[4]), 
            .I3(baudrate[12]), .O(n30785));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16379_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[3]), 
            .I3(baudrate[11]), .O(n30786));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16380_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[2]), 
            .I3(baudrate[10]), .O(n30787));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16381_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[1]), 
            .I3(baudrate[9]), .O(n30788));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16382_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[0]), 
            .I3(baudrate[8]), .O(n30789));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_985 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(byte_counter[2]), .I3(n59009), .O(n62253));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut_adj_985.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_986 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(byte_counter[2]), .I3(GND_net), .O(n3));   // verilog/eeprom.v(68[25:39])
    defparam i1_2_lut_3_lut_adj_986.LUT_INIT = 16'he0e0;
    SB_LUT4 i16367_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30774));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16368_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30775));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16368_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16369_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30776));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16370_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30777));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16370_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16371_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30778));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16371_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16372_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30779));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16372_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16373_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30780));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16373_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16374_3_lut_4_lut (.I0(byte_counter[0]), .I1(n59068), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30781));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16374_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_987 (.I0(\state[2] ), .I1(\state[1] ), .I2(\state_7__N_4045[0] ), 
            .I3(\state[0] ), .O(n4_adj_5120));
    defparam i1_4_lut_adj_987.LUT_INIT = 16'hbbba;
    SB_LUT4 i51825_4_lut (.I0(n5), .I1(n25838), .I2(\state[1] ), .I3(\state[3] ), 
            .O(n67134));
    defparam i51825_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut_adj_988 (.I0(n67134), .I1(n4_adj_5120), .I2(n43931), 
            .I3(\state[0] ), .O(n61958));
    defparam i2_4_lut_adj_988.LUT_INIT = 16'hcfee;
    i2c_controller i2c (.VCC_net(VCC_net), .GND_net(GND_net), .sda_enable(sda_enable), 
            .sda_out(sda_out), .clk16MHz(clk16MHz), .scl_enable(scl_enable), 
            .n6878(n6878), .\state[1] (\state[1]_adj_6 ), .n65(n65), .n62(n62), 
            .\state[2] (\state[2]_adj_5 ), .\state_7__N_4237[0] (\state_7__N_4237[0] ), 
            .\state[3] (\state[3] ), .\state[0] (\state[0]_adj_7 ), .\saved_addr[0] (\saved_addr[0] ), 
            .n30054(n30054), .data({data}), .n30053(n30053), .n30049(n30049), 
            .n58508(n58508), .n30047(n30047), .n30042(n30042), .n30041(n30041), 
            .n28163(n28163), .n49980(n49980), .\state_7__N_4253[3] (\state_7__N_4253[3] ), 
            .n11(n11_adj_8), .enable(enable), .n30841(n30841), .n8(n8), 
            .enable_slow_N_4340(enable_slow_N_4340), .n9(n9), .n10(n10_c), 
            .n29813(n29813), .n10_adj_1(n10), .n44000(n44000), .n11_adj_2(n11), 
            .n4(n4_c), .n4_adj_3(n4_adj_9), .n4_adj_4(n4), .n44006(n44006), 
            .n48(n48), .n25984(n25984), .n49984(n49984), .scl(scl), 
            .n15(n15_adj_5116)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (VCC_net, GND_net, sda_enable, sda_out, clk16MHz, 
            scl_enable, n6878, \state[1] , n65, n62, \state[2] , 
            \state_7__N_4237[0] , \state[3] , \state[0] , \saved_addr[0] , 
            n30054, data, n30053, n30049, n58508, n30047, n30042, 
            n30041, n28163, n49980, \state_7__N_4253[3] , n11, enable, 
            n30841, n8, enable_slow_N_4340, n9, n10, n29813, n10_adj_1, 
            n44000, n11_adj_2, n4, n4_adj_3, n4_adj_4, n44006, n48, 
            n25984, n49984, scl, n15) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    output sda_enable;
    output sda_out;
    input clk16MHz;
    output scl_enable;
    output n6878;
    output \state[1] ;
    input n65;
    input n62;
    output \state[2] ;
    output \state_7__N_4237[0] ;
    output \state[3] ;
    output \state[0] ;
    output \saved_addr[0] ;
    input n30054;
    output [7:0]data;
    input n30053;
    input n30049;
    input n58508;
    input n30047;
    input n30042;
    input n30041;
    input n28163;
    input n49980;
    input \state_7__N_4253[3] ;
    output n11;
    input enable;
    input n30841;
    input n8;
    output enable_slow_N_4340;
    output n9;
    output n10;
    input n29813;
    output n10_adj_1;
    output n44000;
    output n11_adj_2;
    output n4;
    output n4_adj_3;
    output n4_adj_4;
    output n44006;
    output n48;
    output n25984;
    output n49984;
    output scl;
    output n15;
    
    wire i2c_clk /* synthesis SET_AS_NETWORK=\eeprom/i2c/i2c_clk, is_clock=1 */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n52834, n52835, sda_out_adj_5102, n52833, n52832, n52831, 
        i2c_clk_N_4326, n52830, scl_enable_N_4327, n52829;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n52828, n52827, n52826, n52825, n5, n47, n52824, enable_slow_N_4339, 
        n28158, n62148, n60874, n28, n69912, n11_c, n59979, n28145;
    wire [1:0]n6942;
    
    wire n71151, n58372, n28147, n29502, n4_c, n10_c, n9_adj_5105, 
        n61051, n10_adj_5107, n12, n6871, state_7__N_4236, n43912, 
        n11_adj_5109, n11_adj_5110;
    
    SB_LUT4 counter_2067_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n52834), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_8 (.CI(n52834), .I0(VCC_net), .I1(counter[6]), 
            .CO(n52835));
    SB_LUT4 i2499_2_lut (.I0(sda_out_adj_5102), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2067_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n52833), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_7 (.CI(n52833), .I0(VCC_net), .I1(counter[5]), 
            .CO(n52834));
    SB_LUT4 counter_2067_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n52832), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_6 (.CI(n52832), .I0(VCC_net), .I1(counter[4]), 
            .CO(n52833));
    SB_LUT4 counter_2067_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n52831), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_5 (.CI(n52831), .I0(VCC_net), .I1(counter[3]), 
            .CO(n52832));
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4326));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 counter_2067_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n52830), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4327));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_CARRY counter_2067_add_4_4 (.CI(n52830), .I0(VCC_net), .I1(counter[2]), 
            .CO(n52831));
    SB_LUT4 counter_2067_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n52829), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_3 (.CI(n52829), .I0(VCC_net), .I1(counter[1]), 
            .CO(n52830));
    SB_LUT4 counter_2067_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2067_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52829));
    SB_LUT4 counter2_2065_2066_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n52828), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2065_2066_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n52827), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2065_2066_add_4_6 (.CI(n52827), .I0(GND_net), .I1(counter2[4]), 
            .CO(n52828));
    SB_LUT4 counter2_2065_2066_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n52826), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2065_2066_add_4_5 (.CI(n52826), .I0(GND_net), .I1(counter2[3]), 
            .CO(n52827));
    SB_LUT4 counter2_2065_2066_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n52825), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6878), .D(n5), 
            .S(n65));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6878), .D(n62), 
            .S(n47));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_CARRY counter2_2065_2066_add_4_4 (.CI(n52825), .I0(GND_net), .I1(counter2[2]), 
            .CO(n52826));
    SB_LUT4 counter2_2065_2066_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n52824), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2065_2066_add_4_3 (.CI(n52824), .I0(GND_net), .I1(counter2[1]), 
            .CO(n52825));
    SB_LUT4 counter2_2065_2066_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2065_2066_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2065_2066_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n52824));
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4237[0] ), .C(clk16MHz), .E(n28158), 
            .D(enable_slow_N_4339));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6878), .D(n62148), 
            .S(n60874));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i53737_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n69912));
    defparam i53737_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_968 (.I0(n11_c), .I1(n69912), .I2(n28), .I3(n59979), 
            .O(n28145));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1809_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6942[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1809_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i3_4_lut (.I0(n6942[1]), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(\state[2] ), .O(n71151));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i3_4_lut_adj_969 (.I0(n11_c), .I1(n59979), .I2(\state[3] ), 
            .I3(\state[1] ), .O(n58372));
    defparam i3_4_lut_adj_969.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_970 (.I0(n11_c), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n59979), .O(n28147));
    defparam i1_4_lut_adj_970.LUT_INIT = 16'h0a22;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n30054));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30053));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n30049));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n58508));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n30047));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30042));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n30041));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2065_2066__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2065_2066__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2065_2066__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2065_2066__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2065_2066__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_2067__i0 (.Q(counter[0]), .C(i2c_clk), .E(n28163), 
            .D(n37[0]), .S(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFSR counter2_2065_2066__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29502));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_2067__i1 (.Q(counter[1]), .C(i2c_clk), .E(n28163), 
            .D(n37[1]), .S(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESS counter_2067__i2 (.Q(counter[2]), .C(i2c_clk), .E(n28163), 
            .D(n37[2]), .S(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESR counter_2067__i3 (.Q(counter[3]), .C(i2c_clk), .E(n28163), 
            .D(n37[3]), .R(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESR counter_2067__i4 (.Q(counter[4]), .C(i2c_clk), .E(n28163), 
            .D(n37[4]), .R(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESR counter_2067__i5 (.Q(counter[5]), .C(i2c_clk), .E(n28163), 
            .D(n37[5]), .R(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESR counter_2067__i6 (.Q(counter[6]), .C(i2c_clk), .E(n28163), 
            .D(n37[6]), .R(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_DFFESR counter_2067__i7 (.Q(counter[7]), .C(i2c_clk), .E(n28163), 
            .D(n37[7]), .R(n49980));   // verilog/i2c_controller.v(113[18:32])
    SB_LUT4 i1_4_lut_adj_971 (.I0(\state_7__N_4253[3] ), .I1(n11), .I2(n11_c), 
            .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_971.LUT_INIT = 16'h2a2f;
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30841));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i53775_2_lut (.I0(\state_7__N_4237[0] ), .I1(enable_slow_N_4340), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4339));   // verilog/i2c_controller.v(62[6:32])
    defparam i53775_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_310_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_310_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n29502));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29502), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4326));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_308_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(44[32:47])
    defparam equal_308_i10_2_lut.LUT_INIT = 16'heeee;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29813));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 state_7__I_0_139_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5105));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_139_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n28147), 
            .D(n61051), .S(n58372));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_5102), .C(i2c_clk), .E(n28145), 
            .D(n71151), .S(n58372));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_1));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5107));   // verilog/i2c_controller.v(143[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_1), 
            .O(n6871));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29705_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n44000));
    defparam i29705_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53759_4_lut (.I0(state_7__N_4236), .I1(n6871), .I2(n11_adj_2), 
            .I3(n43912), .O(n6878));
    defparam i53759_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n11_adj_5109), .I1(n11), .I2(\state_7__N_4253[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h5755;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5110));   // verilog/i2c_controller.v(139[9:14])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i53801_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4340));   // verilog/i2c_controller.v(44[32:47])
    defparam i53801_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(scl_enable_N_4327));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 counter_2067_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n52835), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2067_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\state[3] ), .I1(n6871), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'hbbbb;
    SB_LUT4 i30425_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n59979));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i30425_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_390_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_390_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_388_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_388_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i29711_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n44006));
    defparam i29711_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(n9_adj_5105), .I1(n10_adj_5107), .I2(counter[0]), 
            .I3(n44006), .O(n48));   // verilog/i2c_controller.v(151[5:14])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9_adj_5105), .I1(n10_adj_5107), .I2(counter[0]), 
            .I3(GND_net), .O(n25984));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i53785_3_lut_4_lut (.I0(n9_adj_5105), .I1(n10_adj_5107), .I2(n11_adj_5110), 
            .I3(n6878), .O(n47));   // verilog/i2c_controller.v(151[5:14])
    defparam i53785_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut_adj_974 (.I0(n9_adj_5105), .I1(n10_adj_5107), 
            .I2(counter[0]), .I3(GND_net), .O(n49984));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_974.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9_adj_5105), .O(n62148));   // verilog/i2c_controller.v(139[9:14])
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'hf0f4;
    SB_LUT4 i29655_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i29655_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_145_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_5109));   // verilog/i2c_controller.v(161[5:14])
    defparam state_7__I_0_145_i11_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i30328_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(state_7__N_4236));
    defparam i30328_3_lut_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 state_7__I_0_139_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_2));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_139_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i30317_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n43912));
    defparam i30317_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 state_7__I_0_140_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(117[5:13])
    defparam state_7__I_0_140_i11_2_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 equal_310_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_310_i11_2_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_adj_976 (.I0(enable), .I1(\state_7__N_4237[0] ), 
            .I2(enable_slow_N_4340), .I3(GND_net), .O(n28158));
    defparam i1_2_lut_3_lut_adj_976.LUT_INIT = 16'haeae;
    SB_LUT4 i54358_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6878), .O(n60874));
    defparam i54358_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 state_7__I_0_143_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_c));   // verilog/i2c_controller.v(143[5:14])
    defparam state_7__I_0_143_i11_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_977 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n61051));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_977.LUT_INIT = 16'h1110;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[14] , \PID_CONTROLLER.integral_23__N_3844[1] , 
            GND_net, \Ki[15] , \Ki[6] , \PID_CONTROLLER.integral_23__N_3844[7] , 
            \Ki[7] , \Ki[8] , \Ki[9] , \Kp[11] , \Ki[10] , \Ki[1] , 
            \PID_CONTROLLER.integral_23__N_3844[0] , \Ki[0] , \Ki[2] , 
            \Ki[11] , \Ki[3] , \Ki[12] , \Ki[13] , \Kp[12] , \Ki[4] , 
            \Kp[13] , \Ki[5] , \Kp[1] , \Kp[0] , \Kp[14] , \Kp[15] , 
            \Kp[2] , \Kp[3] , \Kp[4] , \Kp[5] , deadband, \Kp[6] , 
            \Kp[7] , \Kp[8] , n379, \PID_CONTROLLER.integral_23__N_3844[6] , 
            n4, control_update, \PID_CONTROLLER.integral_23__N_3844[5] , 
            n181, IntegralLimit, n155, \PID_CONTROLLER.integral_23__N_3844[15] , 
            \PID_CONTROLLER.integral_23__N_3844[14] , clk16MHz, \PID_CONTROLLER.integral_23__N_3844[16] , 
            VCC_net, \PID_CONTROLLER.integral , \Kp[9] , \PID_CONTROLLER.integral_23__N_3844[4] , 
            PWMLimit, duty, reset, n149, n136, \PID_CONTROLLER.integral_23__N_3844[22] , 
            \PID_CONTROLLER.integral_23__N_3844[21] , n11, \PID_CONTROLLER.integral_23__N_3844[3] , 
            \Kp[10] , \PID_CONTROLLER.integral_23__N_3844[20] , setpoint, 
            \motor_state[23] , \PID_CONTROLLER.integral_23__N_3844[19] , 
            \PID_CONTROLLER.integral_23__N_3844[17] , n6, n37023, \PID_CONTROLLER.integral_23__N_3844[13] , 
            \motor_state[22] , \PID_CONTROLLER.integral_23__N_3844[23] , 
            n20625, n37, n20626, \motor_state[21] , \PID_CONTROLLER.integral_23__N_3844[12] , 
            n188, \motor_state[20] , \PID_CONTROLLER.integral_23__N_3844[11] , 
            \motor_state[19] , \motor_state[18] , \motor_state[17] , \PID_CONTROLLER.integral_23__N_3844[2] , 
            \motor_state[16] , \motor_state[15] , \motor_state[14] , n10, 
            \motor_state[12] , n51273, \motor_state[11] , \motor_state[10] , 
            \motor_state[9] , \motor_state[8] , \motor_state[7] , \motor_state[6] , 
            \motor_state[5] , \PID_CONTROLLER.integral_23__N_3844[10] , 
            \motor_state[4] , \motor_state[3] , \motor_state[2] , \motor_state[1] , 
            n34987, \motor_state[0] , \PID_CONTROLLER.integral_23__N_3844[9] , 
            \PID_CONTROLLER.integral_23__N_3844[8] , n30012, n30827, n30826, 
            n30825, n30824, n30823, n30822, n30821, n30820, n30819, 
            n30818, n30817, n30816, n30815, n30814, n30813, n30812, 
            n30811, n30810, n30809, n30808, n30807, n30806, n30805, 
            n219, n405, n38, n28, n110, n20576, n20577, n56) /* synthesis syn_module_defined=1 */ ;
    input \Ki[14] ;
    output \PID_CONTROLLER.integral_23__N_3844[1] ;
    input GND_net;
    input \Ki[15] ;
    input \Ki[6] ;
    output \PID_CONTROLLER.integral_23__N_3844[7] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Kp[11] ;
    input \Ki[10] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.integral_23__N_3844[0] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[11] ;
    input \Ki[3] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Kp[12] ;
    input \Ki[4] ;
    input \Kp[13] ;
    input \Ki[5] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input [23:0]deadband;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    output n379;
    output \PID_CONTROLLER.integral_23__N_3844[6] ;
    input n4;
    output control_update;
    output \PID_CONTROLLER.integral_23__N_3844[5] ;
    output n181;
    input [23:0]IntegralLimit;
    output n155;
    output \PID_CONTROLLER.integral_23__N_3844[15] ;
    output \PID_CONTROLLER.integral_23__N_3844[14] ;
    input clk16MHz;
    output \PID_CONTROLLER.integral_23__N_3844[16] ;
    input VCC_net;
    output [23:0]\PID_CONTROLLER.integral ;
    input \Kp[9] ;
    output \PID_CONTROLLER.integral_23__N_3844[4] ;
    input [23:0]PWMLimit;
    output [23:0]duty;
    input reset;
    output n149;
    output n136;
    output \PID_CONTROLLER.integral_23__N_3844[22] ;
    output \PID_CONTROLLER.integral_23__N_3844[21] ;
    input n11;
    output \PID_CONTROLLER.integral_23__N_3844[3] ;
    input \Kp[10] ;
    output \PID_CONTROLLER.integral_23__N_3844[20] ;
    input [23:0]setpoint;
    input \motor_state[23] ;
    output \PID_CONTROLLER.integral_23__N_3844[19] ;
    output \PID_CONTROLLER.integral_23__N_3844[17] ;
    input n6;
    input n37023;
    output \PID_CONTROLLER.integral_23__N_3844[13] ;
    input \motor_state[22] ;
    output \PID_CONTROLLER.integral_23__N_3844[23] ;
    output n20625;
    input n37;
    output n20626;
    input \motor_state[21] ;
    input \PID_CONTROLLER.integral_23__N_3844[12] ;
    output n188;
    input \motor_state[20] ;
    output \PID_CONTROLLER.integral_23__N_3844[11] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    output \PID_CONTROLLER.integral_23__N_3844[2] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input n10;
    input \motor_state[12] ;
    output n51273;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    output \PID_CONTROLLER.integral_23__N_3844[10] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    output n34987;
    input \motor_state[0] ;
    output \PID_CONTROLLER.integral_23__N_3844[9] ;
    output \PID_CONTROLLER.integral_23__N_3844[8] ;
    input n30012;
    input n30827;
    input n30826;
    input n30825;
    input n30824;
    input n30823;
    input n30822;
    input n30821;
    input n30820;
    input n30819;
    input n30818;
    input n30817;
    input n30816;
    input n30815;
    input n30814;
    input n30813;
    input n30812;
    input n30811;
    input n30810;
    input n30809;
    input n30808;
    input n30807;
    input n30806;
    input n30805;
    output n219;
    output n405;
    input n38;
    output n28;
    input n110;
    input n20576;
    input n20577;
    input n56;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n1026, n1099, n460, n533, n606, n679;
    wire [23:0]n356;
    wire [23:0]n382;
    
    wire n71255, n67829, n69071;
    wire [23:0]n1;
    
    wire n828, n71281, n752, n69657, n74, n5, n147, n825, n220, 
        n71246, n898, n971, n1044, n901, n293, n974, n1117, 
        n366_adj_4560, n119, n50, n1047, n1120, n69841, n192, 
        n71243, n265, n338, n19, n10_c, n411, n11_c, n9, n68794, 
        n484, n17, n15, n13, n69123, n439, n512, n557, n585, 
        n658, n23, n21, n69121, n630, n29, n27, n25, n67956, 
        n731, n804, n66952, n6_c, n69326, n35, n14, n12, n37_c, 
        n32, n92, n877, n23_adj_4561, n165, n950, n1023, n1096, 
        n67921, n31, n69327, n33, n67899, n67877, n69581, n68182, 
        n6_adj_4562, n238, n69322, n69323, n69320, n69321, n71251, 
        n68690, n67817, n71277, n30, n10_adj_4563, n67815, n69583, 
        n68192, n69807, n69808, n69796, n71265, n68698, n67801, 
        n24, n8, n71241, n67799, n69175, n68190, n67807, n311, 
        n384_adj_4564, n457, n69484, n68198, n8_adj_4565, n530, 
        n69328, n69329, n603, n68013, n68764, n69171, n676, n749, 
        n68180, n69436, n69805, n69420, n822, n69885, n895, n968, 
        n69886, n69719, n69629, n69630, n1041, n69695, n63914, 
        n47, n62203, n1114, n89, n20, n162, n235, n308, n381, 
        n454, n527, n600, n673, n746, n819, n892, n965;
    wire [23:0]n130;
    wire [23:0]n182;
    wire [23:0]n207;
    
    wire n116, n47_adj_4566, n119_adj_4567, counter_31__N_3843, n189, 
        n50_adj_4568, n1038, n74_adj_4569;
    wire [23:0]n1_adj_5099;
    
    wire n51539, n5_adj_4571, n1111, n51540, n51538, n192_adj_4573, 
        n116_adj_4574, n47_adj_4575, n189_adj_4576, n262, n265_adj_4577, 
        n335, n408, n481, n51458, n51459, n338_adj_4579, n554, 
        n411_adj_4580, n627, n51457, n700, n86;
    wire [18:0]n15358;
    wire [17:0]n16118;
    
    wire n51912;
    wire [23:0]n436;
    
    wire n12030, n28308, n17_adj_4582, n12028;
    wire [23:0]n49;
    
    wire n51911, n484_adj_4583, n28303, n28298, n159, n51910, n232, 
        n28293, n305, n51456, n378_adj_4585, n28288, n77, n8_adj_4586, 
        n557_adj_4587, n28283, n150, n28278, n630_adj_4589, n451, 
        n28273, n95, n26, n168, n28268, n51909, n262_adj_4591, 
        n51455, n28263, n335_adj_4592, n1108, n51908, n223, n241, 
        n28258, n147_adj_4593, n314, n28253, n408_adj_4595, n524, 
        n387_adj_4596, n220_adj_4597, n28248, n28243, n597, n670, 
        n296, n460_adj_4598, n28238, n1035, n51907, n743, n481_adj_4599, 
        n293_adj_4600, n533_adj_4601, n816, n28233, n28228, n962, 
        n51906, n889, n51905, n816_adj_4602, n51904, n743_adj_4603, 
        n51903, n51454, n670_adj_4605, n51902, n51453, n554_adj_4606, 
        n597_adj_4607, n51901, n627_adj_4608, n41, n51452, n51451, 
        n889_adj_4610, n28223, n39, n45, n524_adj_4611, n51900, 
        n451_adj_4612, n51899, n51450, n43, n37_adj_4613, n23_adj_4614, 
        n369_adj_4615, n378_adj_4616, n51898, n25_adj_4617, n41_adj_4618, 
        n28218, n305_adj_4619, n51897, n232_adj_4620, n51896, n39_adj_4621, 
        n45_adj_4622, n43_adj_4624, n29_adj_4625, n37_adj_4626, n31_adj_4627, 
        n29_adj_4628, n35_adj_4629, n33_adj_4630, n31_adj_4631, n606_adj_4632, 
        n51449, n28213, n962_adj_4634, n9_adj_4635, n23_adj_4636, 
        n25_adj_4638, n159_adj_4639, n51895, n17_adj_4640, n1035_adj_4641, 
        n51448, n28208, n17_adj_4642, n86_adj_4643, n19_adj_4645, 
        n35_adj_4646, n21_adj_4647, n13_adj_4648;
    wire [1:0]n20670;
    
    wire n442_adj_4649, n515, n28203, n1108_adj_4650, n51447, n51027, 
        n15_adj_4651, n27_adj_4652, n67535, n67520, n12_adj_4654;
    wire [10:0]n19534;
    wire [9:0]n19798;
    
    wire n840, n51675, n10_adj_4655, n30_adj_4656, n33_adj_4657, n11_adj_4658, 
        n13_adj_4659, n15_adj_4660, n27_adj_4661, n67578, n68472, 
        n9_adj_4662, n68458, n767, n51674, n69571, n17_adj_4663, 
        n588, n679_adj_4664, n28198, n68951, n19_adj_4666, n83, 
        n51446, n14_adj_4667, n752_adj_4668, n156, n229, n302, n661;
    wire [2:0]n20653;
    
    wire n51191, n69705, n16, n6_adj_4669, n68965, n375_adj_4670, 
        n448_adj_4671, n21_adj_4672, n521, n694, n51673, n67713, 
        n68966, n51445, n621, n51672;
    wire [0:0]n12063;
    wire [21:0]n12570;
    
    wire n52069;
    wire [47:0]n257;
    
    wire n52068, n67707, n12_adj_4673, n8_adj_4674, n24_adj_4675, 
        n10_adj_4676, n594, n30_adj_4677, n667, n825_adj_4678, n67478, 
        n67443, n69161, n68168, n4_adj_4679, n68963, n68964, n67503, 
        n67729, n68608, n67499, n69370, n68602, n69641, n4_adj_4680;
    wire [3:0]n20622;
    
    wire n69021, n6_adj_4681, n734, n69742, n740, n51223, n68170, 
        n69799, n813, n69800, n69715, n6_adj_4682, n69249, n67480, 
        n16_adj_4683, n69478, n886, n68176, n69689, n548, n51671, 
        n959, n39_adj_4684, n41_adj_4685, n25_adj_4686, n45_adj_4687, 
        n1032, n23_adj_4688, n43_adj_4689, n8_adj_4690, n898_adj_4691, 
        n29_adj_4693, n31_adj_4694, n24_adj_4695, n35_adj_4697, n33_adj_4698, 
        n11_adj_4699, n125_adj_4700, n1105, n198, n13_adj_4702, n69250, 
        n15_adj_4703, n52067, n67678, n27_adj_4704, n9_adj_4705, n271, 
        n67676, n69179, n68210, n807, n344, n475, n51670, n417;
    wire [4:0]n20573;
    
    wire n41_adj_4711, n17_adj_4713, n19_adj_4714, n21_adj_4715, n67400, 
        n67369, n4_adj_4717, n52066, n12_adj_4718, n10_adj_4719, n69247, 
        n30_adj_4720, n51444, n69248, n67435, n68305, n402, n51669, 
        n67698, n971_adj_4721, n490, n880, n63894, n63898, n63896, 
        n68291, n113_adj_4722, n44_adj_4723, n63904, n4_adj_4724, 
        n8_adj_4725, n69512, n61143, n68874, n69681, n16_adj_4727, 
        n186_adj_4728, n6_adj_4729, n68957, n67696, n69611, n51443, 
        n68212, n259, n1044_adj_4732, n183, n68958, n107_adj_4733, 
        n38_adj_4734, n8_adj_4736, n24_adj_4738, n256, n69817, n69818, 
        n1117_adj_4739, n180, n52065, n69781, n329, n253, n402_adj_4743, 
        n326, n68037, n68033, n69167, n68178, n4_adj_4745, n67682, 
        n399, n69488, n68218, n332, n472, n953, n69424, n545, 
        n475_adj_4749, n69425, n67241, n113_adj_4750, n44_adj_4751, 
        n186_adj_4752, n67232, n69717, n69164, n37361, n69863, n69864, 
        n69824;
    wire [23:0]n1_adj_5100;
    
    wire n259_adj_4754, n69699, n69700, n409, n68041, n69691, n618, 
        n28153, n332_adj_4755, n40_adj_4756, n405_c, n69693, n405_adj_4757, 
        n691, n548_adj_4759, n478, n700_adj_4760, n478_adj_4761, n621_adj_4762, 
        n551, n694_adj_4763, n624, n764, n551_adj_4764, n51442, 
        n767_adj_4765, n697, n840_adj_4766, n770, n837, n107_adj_4767, 
        n83_adj_4768, n14_adj_4769, n156_adj_4770, n89_adj_4772, n20_adj_4773, 
        n162_adj_4774, n180_adj_4775, n1026_adj_4776, n229_adj_4777, 
        n253_adj_4778, n326_adj_4779, n302_adj_4780, n375_adj_4781, 
        n366_adj_4783, n624_adj_4784, n448_adj_4785, n697_adj_4786, 
        n329_adj_4787, n51668, n521_adj_4788, n594_adj_4789, n256_adj_4790, 
        n51667, n667_adj_4791, n740_adj_4792, n813_adj_4793, n399_adj_4794, 
        n886_adj_4795, n52064, n910;
    wire [16:0]n16802;
    
    wire n51880, n770_adj_4796, n51441, n52063, n183_adj_4798, n51666, 
        n959_adj_4799, n51879, n1032_adj_4800, n51440, n1105_adj_4803, 
        n41_adj_4804, n110_adj_4805, n51878, n52062, n51439, n1096_adj_4807, 
        n52061, n1111_adj_4808, n51877, n1038_adj_4809, n51876, n965_adj_4812, 
        n51875, n1023_adj_4814, n52060, n472_adj_4816, n892_adj_4817, 
        n51874, n80, n11_adj_4819, n51438, n545_adj_4820, n104, 
        n819_adj_4822, n51873, n35_adj_4823, n153_adj_4824, n746_adj_4826, 
        n51872, n177, n618_adj_4827, n250, n950_adj_4829, n52059, 
        n691_adj_4831, n877_adj_4834, n52058, n673_adj_4835, n51871, 
        n764_adj_4836, n51437, n804_adj_4837, n52057, n51436, n731_adj_4838, 
        n52056, n600_adj_4839, n51870, n527_adj_4840, n51869, n837_adj_4841, 
        n910_adj_4842, n323, n658_adj_4844, n52055, n51435, n454_adj_4848, 
        n51868, n396_adj_4849, n51434, n381_adj_4850, n51867, n469, 
        n308_adj_4851, n51866, n125_adj_4852, n56_adj_4853, n542, 
        n585_adj_4855, n52054, n51433, n198_adj_4857, n51432, n512_adj_4858, 
        n52053, n439_adj_4859, n52052, n235_adj_4861, n51865, n615, 
        n52051, n51864, n688, n761, n51431;
    wire [8:0]n20117;
    wire [7:0]n20278;
    
    wire n51863, n271_adj_4864, n51862;
    wire [23:0]n1_adj_5101;
    
    wire n51861, n51430, n834, n907, n51429, n51428, n52050, n980, 
        n51860, n52049, n344_adj_4867, n51859;
    wire [47:0]n306;
    
    wire n52048, n51858, n51857, n417_adj_4877;
    wire [3:0]n20598;
    
    wire n6_adj_4878;
    wire [4:0]n20538;
    
    wire n51427, n80_adj_4879, n11_adj_4880, n204_adj_4881, n226;
    wire [1:0]n20662;
    
    wire n131_adj_4882, n62_adj_4883, n490_adj_4884, n63928, n63930, 
        n210, n63934, n51257, n63938, n8_adj_4885, n6_adj_4886, 
        n4_adj_4887, n61880, n51856, n104_adj_4888, n35_adj_4889, 
        n51426, n122_adj_4891, n53, n153_adj_4892, n195_adj_4893, 
        n177_adj_4895, n268, n226_adj_4897, n250_adj_4899, n341, n414, 
        n299_adj_4901, n372_adj_4903, n323_adj_4904, n487, n560, n101, 
        n32_adj_4906, n445_adj_4907, n396_adj_4908, n174, n247, n51425, 
        n320, n518, n393_adj_4911, n466, n591, n539, n612, n664, 
        n51424, n737, n685, n758, n469_adj_4916, n831, n51423, 
        n810, n904, n883, n977, n299_adj_4919, n1050, n956, n1029, 
        n1102, n542_adj_4920, n1099_adj_4921, n615_adj_4922, n688_adj_4923, 
        n761_adj_4924, n834_adj_4925, n907_adj_4926, n980_adj_4927, 
        n101_adj_4928, n32_adj_4929, n174_adj_4930, n247_adj_4931, n320_adj_4932, 
        n393_adj_4933, n466_adj_4934, n539_adj_4935, n98, n29_adj_4936, 
        n612_adj_4937, n685_adj_4938, n758_adj_4939;
    wire [15:0]n17414;
    
    wire n51842, n51841, n1114_adj_4940, n51840, n831_adj_4941, n904_adj_4942, 
        n977_adj_4943, n1050_adj_4944, n122_adj_4945, n53_adj_4946, 
        n195_adj_4947, n268_adj_4948, n341_adj_4949, n414_adj_4950, 
        n487_adj_4951, n560_adj_4952, n98_adj_4953, n29_adj_4954, n171, 
        n244, n1041_adj_4955, n51839, n171_adj_4956, n317, n390_adj_4957, 
        n463, n968_adj_4958, n51838, n244_adj_4959, n536, n317_adj_4960, 
        n390_adj_4961, n895_adj_4962, n51837, n822_adj_4963, n51836, 
        n609, n463_adj_4964, n682, n755, n536_adj_4965, n828_adj_4966, 
        n901_adj_4967, n974_adj_4968, n1047_adj_4969, n609_adj_4970, 
        n1120_adj_4971, n95_adj_4972, n26_adj_4973, n168_adj_4974, n749_adj_4975, 
        n51835, n241_adj_4976, n682_adj_4977, n314_adj_4978, n755_adj_4979, 
        n387_adj_4980, n372_adj_4981, n676_adj_4982, n51834, n603_adj_4983, 
        n51833, n530_adj_4984, n51832, n457_adj_4985, n51831, n384_adj_4986, 
        n51830, n311_adj_4987, n51829, n238_adj_4988, n51828;
    wire [31:0]n51;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n165_adj_5015, n51827;
    wire [20:0]n13590;
    
    wire n52029, n23_adj_5016, n92_adj_5017, n52028, n52027, n52026, 
        n445_adj_5018, n52025;
    wire [0:0]n12598;
    wire [21:0]n13105;
    
    wire n53109, n53108, n53107, n53106, n53105, n53104, n53103, 
        n53102, n53101, n53100, n53099, n53098, n53097, n53096, 
        n53095, n53094, n53093, n53092, n53091, n53090, n53089, 
        n53088;
    wire [20:0]n14074;
    
    wire n53087, n53086, n53085, n53084, n53083, n53082, n53081, 
        n53080, n53079, n953_adj_5024, n53078, n880_adj_5025, n53077, 
        n807_adj_5026, n53076, n734_adj_5027, n53075, n661_adj_5028, 
        n53074, n588_adj_5029, n53073, n515_adj_5030, n53072, n442_adj_5031, 
        n53071, n369_adj_5032, n53070, n296_adj_5033, n53069, n223_adj_5034, 
        n53068, n150_adj_5035, n53067, n12_adj_5036, n8_adj_5037, 
        n77_adj_5038, n11_adj_5039, n62077, n18_adj_5040, n10_adj_5041, 
        n16_adj_5042, n15_adj_5043, n24_adj_5044, n23_adj_5045;
    wire [19:0]n14958;
    
    wire n53066, n53065, n25_adj_5046, n53064, n53063, n53062, n53061, 
        n52024, n1102_adj_5047, n53060, n1029_adj_5048, n53059, n956_adj_5049, 
        n53058, n883_adj_5050, n53057, n810_adj_5051, n53056, n737_adj_5052, 
        n53055, n51491, n664_adj_5053, n53054, n591_adj_5054, n53053, 
        n518_adj_5056, n53052, n53051, n52733, n52732, n52731, n52730, 
        n53050, n52729, n52023, n52022, n51490, n53049, n52728, 
        n53048, n53047, n52727, n51489;
    wire [8:0]n20018;
    
    wire n53046, n53045, n53044, n52021, n52726, n53043, n53042, 
        n53041, n51488, n52020, n53040;
    wire [14:0]n17958;
    
    wire n51814, n51813, n51487, n51812, n53039, n53038, n52019;
    wire [18:0]n15757;
    
    wire n53037, n53036, n53035, n51811, n53034, n53033, n52018, 
        n53032, n51810, n53031, n52725, n53030, n53029, n53028, 
        n53027, n52017, n51809, n53026, n52724, n53025, n53024, 
        n53023, n53022, n52016, n53021, n53020, n52723, n53019, 
        n51808;
    wire [17:0]n16478;
    
    wire n53018, n52722, n53017, n53016, n51807, n53015, n52015, 
        n52721, n53014, n52014, n52013, n53013, n52720, n53012, 
        n51806, n52012, n53011, n52719, n53010, n51486, n51805, 
        n52718, n53009, n51804, n52011, n53008, n53007, n51803, 
        n52717, n53006, n51485, n51802, n51484, n51801, n52010, 
        n51800, n52716, n53005, n51483;
    wire [6:0]n20405;
    
    wire n51799, n52009, n51798, n53004, n53003, n53002, n52715, 
        n53001, n51797, n52714;
    wire [7:0]n20198;
    
    wire n53000, n52999, n51796, n52713, n52998, n51795, n52997, 
        n52996, n52995, n51794, n52994, n52993, n52712;
    wire [16:0]n17125;
    
    wire n52992, n52991, n51482, n51793, n52990, n52989, n52988, 
        n52711, n52987, n52986, n52985, n52710, n52984, n52983, 
        n52709, n52982, n52708, n52981, n52980, n51481, n52979, 
        n52707, n52978, n52706, n52977, n52705, n52704, n52976, 
        n52703;
    wire [15:0]n17702;
    
    wire n52975, n52974, n52973, n52972, n52971, n52970, n52969, 
        n52968, n52967, n52966, n52965, n52964, n52963, n52962, 
        n52961, n52960;
    wire [6:0]n20342;
    
    wire n52959, n52958, n52957, n52956, n52955, n52954, n52953;
    wire [13:0]n18438;
    
    wire n51781, n51780;
    wire [14:0]n18213;
    
    wire n52952, n51480, n52951, n51779, n51778, n52950, n51479, 
        n52949, n52948, n52947, n52946, n51777, n52945, n52944, 
        n52943, n52942, n52941, n51776, n52940, n51775, n52939, 
        n52938, n51478;
    wire [13:0]n18662;
    
    wire n52937, n51774, n52936, n52935, n52934, n52933, n51773, 
        n52932, n52931, n51477, n51772, n52930, n51771;
    wire [19:0]n14518;
    
    wire n51991, n51770, n52929, n51769, n51990, n52928, n51476, 
        n52927, n52926, n51768, n52925, n51989, n52924;
    wire [5:0]n20454;
    
    wire n52923, n52922, n52921, n52920, n52919, n39_adj_5059, n41_adj_5060, 
        n45_adj_5061, n52918, n43_adj_5062, n23_adj_5063;
    wire [12:0]n19053;
    
    wire n52917, n52916, n25_adj_5065, n52915, n52914, n52913, n52912, 
        n52911, n52910, n52909, n29_adj_5066, n31_adj_5067, n37_adj_5068, 
        n35_adj_5069, n52908, n52907, n52906, n33_adj_5070, n11_adj_5071, 
        n51988, n52905;
    wire [11:0]n19390;
    
    wire n52904, n13_adj_5072, n15_adj_5073, n51987, n52903, n52902, 
        n52901, n52900, n27_adj_5074, n9_adj_5075, n52899, n51475, 
        n51986, n52898, n51985, n51984, n51474, n51983;
    wire [12:0]n18858;
    
    wire n51757, n51756, n51982, n51606, n51755, n51981, n51754, 
        n51605, n52897, n51753, n51604, n51752, n51980, n51603, 
        n51979, n51751, n51602, n17_adj_5076, n51750, n51601, n51978, 
        n51749, n51748, n51473, n51977, n51747, n51472, n51600, 
        n51746, n51599, n51745, n52896, n51976, n19_adj_5077, n51598;
    wire [5:0]n20502;
    
    wire n51744, n51743, n52895, n51975, n51471, n51597, n21_adj_5078, 
        n51974, n51742, n51596, n51741, n52894, n51595, n51973, 
        n51594, n51740, n52893, n51593, n51739, n51972, n51592, 
        n52892, n67772, n52891, n51470, n51591, n51469, n51590, 
        n51589, n51588, n51587, n51586, n51585, n51584, n52890;
    wire [11:0]n19222;
    
    wire n51729, n51728, n51727, n52889, n51468, n51726, n51725, 
        n51467, n51583, n51582, n51724, n51581, n52888, n51580, 
        n51723, n51579, n51722, n51721, n51578, n51466, n51577, 
        n51720;
    wire [10:0]n19677;
    
    wire n52887, n52886, n52885, n51576, n52884, n51575, n51465, 
        n51719, n51574, n52883, n51718, n51464, n51573, n51572, 
        n52882, n51463, n51571, n51955, n52881, n51462, n51570, 
        n51954, n51569, n51953, n51568, n51952, n51461, n51951, 
        n51567, n67758, n51566, n51950, n51565, n51564, n51949, 
        n51948, n51563, n51709, n51947, n52880, n51946, n51945, 
        n51944, n51943, n51942, n51941, n51562, n51940, n51939, 
        n52879, n52878, n51938, n52877, n51561, n51937, n51708;
    wire [9:0]n19918;
    
    wire n51936, n52876, n51935, n52875, n51707, n51934, n52874, 
        n51933, n52873, n51932, n52872, n51706, n51931, n51930, 
        n51705, n51929, n51928, n51560, n51559, n52871, n51704, 
        n51460, n51558, n51703, n51557, n51702, n51556, n51555, 
        n51701, n51554, n52870, n51553, n51700, n51552, n52869, 
        n51551, n51699, n52868, n51550, n51549, n52867, n51548, 
        n51547, n51698, n51697, n51546, n51545, n51696, n51544, 
        n51543, n51542, n12_adj_5086, n10_adj_5087, n30_adj_5088, 
        n67793, n68658, n68650, n69651, n69043, n69744, n16_adj_5089, 
        n6_adj_5090, n69312, n69313, n8_adj_5091, n24_adj_5092, n67733, 
        n67731, n69177, n68200, n4_adj_5093, n51695, n69302, n69303, 
        n67750, n67744, n69597, n68202, n69813, n69814, n69789, 
        n67735, n69486, n68208, n69697, n51694, n51541, n67845, 
        n68706, n71257, n12_adj_5095, n67837, n68702, n71270, n16_adj_5096, 
        n67849, n71296, n67847, n71289, n69077, n71292, n68704, 
        n69432, n4_adj_5097, n51141;
    wire [2:0]n20638;
    
    wire n4_adj_5098, n51002;
    
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i29_rep_146_2_lut (.I0(n356[14]), .I1(n382[14]), 
            .I2(GND_net), .I3(GND_net), .O(n71255));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i29_rep_146_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52896_4_lut (.I0(n356[15]), .I1(n71255), .I2(n382[15]), .I3(n67829), 
            .O(n69071));
    defparam i52896_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i33_rep_172_2_lut (.I0(n356[16]), .I1(n382[16]), 
            .I2(GND_net), .I3(GND_net), .O(n71281));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i33_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53482_4_lut (.I0(n356[17]), .I1(n71281), .I2(n382[17]), .I3(n69071), 
            .O(n69657));
    defparam i53482_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i37_rep_137_2_lut (.I0(n356[18]), .I1(n382[18]), 
            .I2(GND_net), .I3(GND_net), .O(n71246));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i37_rep_137_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53666_4_lut (.I0(n356[19]), .I1(n71246), .I2(n382[19]), .I3(n69657), 
            .O(n69841));
    defparam i53666_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_21_i41_rep_134_2_lut (.I0(n356[20]), .I1(n382[20]), 
            .I2(GND_net), .I3(GND_net), .O(n71243));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i41_rep_134_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n356[5]), .I1(n356[9]), .I2(n19), 
            .I3(GND_net), .O(n10_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52619_4_lut (.I0(n11_c), .I1(n9), .I2(deadband[3]), .I3(n356[3]), 
            .O(n68794));
    defparam i52619_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52948_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n68794), 
            .O(n69123));
    defparam i52948_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52946_4_lut (.I0(n23), .I1(n21), .I2(n19), .I3(n69123), 
            .O(n69121));
    defparam i52946_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51782_4_lut (.I0(n29), .I1(n27), .I2(n25), .I3(n69121), 
            .O(n67956));
    defparam i51782_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51126_4_lut (.I0(deadband[1]), .I1(n356[0]), .I2(n379), .I3(deadband[0]), 
            .O(n66952));   // verilog/motorControl.v(51[12:29])
    defparam i51126_4_lut.LUT_INIT = 16'h50d4;
    SB_LUT4 LessThan_19_i6_3_lut (.I0(n66952), .I1(n356[2]), .I2(deadband[2]), 
            .I3(GND_net), .O(n6_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53151_3_lut (.I0(n6_c), .I1(n356[14]), .I2(n29), .I3(GND_net), 
            .O(n69326));   // verilog/motorControl.v(51[12:29])
    defparam i53151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i14_3_lut (.I0(n356[8]), .I1(n356[17]), .I2(n35), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n356[6]), .I1(n356[7]), .I2(n15), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i32_3_lut (.I0(n14), .I1(n356[18]), .I2(n37_c), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4561));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51747_4_lut (.I0(n29), .I1(n17), .I2(n15), .I3(n13), .O(n67921));
    defparam i51747_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53152_3_lut (.I0(n69326), .I1(n356[15]), .I2(n31), .I3(GND_net), 
            .O(n69327));   // verilog/motorControl.v(51[12:29])
    defparam i53152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51725_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n67921), 
            .O(n67899));
    defparam i51725_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53406_4_lut (.I0(n32), .I1(n12), .I2(n37_c), .I3(n67877), 
            .O(n69581));   // verilog/motorControl.v(51[12:29])
    defparam i53406_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52008_3_lut (.I0(n69327), .I1(n356[16]), .I2(n33), .I3(GND_net), 
            .O(n68182));   // verilog/motorControl.v(51[12:29])
    defparam i52008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n382[2]), .I1(n382[3]), .I2(n356[3]), 
            .I3(GND_net), .O(n6_adj_4562));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53147_3_lut (.I0(n6_adj_4562), .I1(n382[10]), .I2(n356[10]), 
            .I3(GND_net), .O(n69322));   // verilog/motorControl.v(51[33:53])
    defparam i53147_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53148_3_lut (.I0(n69322), .I1(n382[11]), .I2(n356[11]), .I3(GND_net), 
            .O(n69323));   // verilog/motorControl.v(51[33:53])
    defparam i53148_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53145_3_lut (.I0(n4), .I1(n382[13]), .I2(n356[13]), .I3(GND_net), 
            .O(n69320));   // verilog/motorControl.v(51[33:53])
    defparam i53145_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53146_3_lut (.I0(n69320), .I1(n382[14]), .I2(n356[14]), .I3(GND_net), 
            .O(n69321));   // verilog/motorControl.v(51[33:53])
    defparam i53146_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51643_4_lut (.I0(n356[16]), .I1(n71251), .I2(n382[16]), .I3(n68690), 
            .O(n67817));
    defparam i51643_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i35_rep_168_2_lut (.I0(n356[17]), .I1(n382[17]), 
            .I2(GND_net), .I3(GND_net), .O(n71277));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i35_rep_168_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53408_4_lut (.I0(n30), .I1(n10_adj_4563), .I2(n71277), .I3(n67815), 
            .O(n69583));   // verilog/motorControl.v(51[33:53])
    defparam i53408_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52018_3_lut (.I0(n69321), .I1(n382[15]), .I2(n356[15]), .I3(GND_net), 
            .O(n68192));   // verilog/motorControl.v(51[33:53])
    defparam i52018_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53632_4_lut (.I0(n68192), .I1(n69583), .I2(n71277), .I3(n67817), 
            .O(n69807));   // verilog/motorControl.v(51[33:53])
    defparam i53632_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53633_3_lut (.I0(n69807), .I1(n382[18]), .I2(n356[18]), .I3(GND_net), 
            .O(n69808));   // verilog/motorControl.v(51[33:53])
    defparam i53633_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53621_3_lut (.I0(n69808), .I1(n382[19]), .I2(n356[19]), .I3(GND_net), 
            .O(n69796));   // verilog/motorControl.v(51[33:53])
    defparam i53621_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51627_4_lut (.I0(n356[21]), .I1(n71265), .I2(n382[21]), .I3(n68698), 
            .O(n67801));
    defparam i51627_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i53000_4_lut (.I0(n24), .I1(n8), .I2(n71241), .I3(n67799), 
            .O(n69175));   // verilog/motorControl.v(51[33:53])
    defparam i53000_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52016_3_lut (.I0(n69323), .I1(n382[12]), .I2(n356[12]), .I3(GND_net), 
            .O(n68190));   // verilog/motorControl.v(51[33:53])
    defparam i52016_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51633_4_lut (.I0(n356[21]), .I1(n71243), .I2(n382[21]), .I3(n69841), 
            .O(n67807));
    defparam i51633_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i45_rep_132_2_lut (.I0(n356[22]), .I1(n382[22]), 
            .I2(GND_net), .I3(GND_net), .O(n71241));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i45_rep_132_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4564));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53309_4_lut (.I0(n68190), .I1(n69175), .I2(n71241), .I3(n67801), 
            .O(n69484));   // verilog/motorControl.v(51[33:53])
    defparam i53309_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52024_3_lut (.I0(n69796), .I1(n382[20]), .I2(n356[20]), .I3(GND_net), 
            .O(n68198));   // verilog/motorControl.v(51[33:53])
    defparam i52024_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n356[3]), .I1(n356[4]), .I2(n9), 
            .I3(GND_net), .O(n8_adj_4565));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53153_3_lut (.I0(n8_adj_4565), .I1(n356[11]), .I2(n23), .I3(GND_net), 
            .O(n69328));   // verilog/motorControl.v(51[12:29])
    defparam i53153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53154_3_lut (.I0(n69328), .I1(n356[12]), .I2(n25), .I3(GND_net), 
            .O(n69329));   // verilog/motorControl.v(51[12:29])
    defparam i53154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52589_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n68013), 
            .O(n68764));
    defparam i52589_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52996_3_lut (.I0(n10_c), .I1(n356[10]), .I2(n21), .I3(GND_net), 
            .O(n69171));   // verilog/motorControl.v(51[12:29])
    defparam i52996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52006_3_lut (.I0(n69329), .I1(n356[13]), .I2(n27), .I3(GND_net), 
            .O(n68180));   // verilog/motorControl.v(51[12:29])
    defparam i52006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53261_4_lut (.I0(n35), .I1(n33), .I2(n31), .I3(n67956), 
            .O(n69436));
    defparam i53261_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53630_4_lut (.I0(n68182), .I1(n69581), .I2(n37_c), .I3(n67899), 
            .O(n69805));   // verilog/motorControl.v(51[12:29])
    defparam i53630_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53245_4_lut (.I0(n68180), .I1(n69171), .I2(n27), .I3(n68764), 
            .O(n69420));   // verilog/motorControl.v(51[12:29])
    defparam i53245_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53710_4_lut (.I0(n69420), .I1(n69805), .I2(n37_c), .I3(n69436), 
            .O(n69885));   // verilog/motorControl.v(51[12:29])
    defparam i53710_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53711_3_lut (.I0(n69885), .I1(n356[19]), .I2(deadband[19]), 
            .I3(GND_net), .O(n69886));   // verilog/motorControl.v(51[12:29])
    defparam i53711_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53544_3_lut (.I0(n69886), .I1(n356[20]), .I2(deadband[20]), 
            .I3(GND_net), .O(n69719));   // verilog/motorControl.v(51[12:29])
    defparam i53544_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53454_3_lut (.I0(n69719), .I1(n356[21]), .I2(deadband[21]), 
            .I3(GND_net), .O(n69629));   // verilog/motorControl.v(51[12:29])
    defparam i53454_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53455_3_lut (.I0(n69629), .I1(n356[22]), .I2(deadband[22]), 
            .I3(GND_net), .O(n69630));   // verilog/motorControl.v(51[12:29])
    defparam i53455_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53520_4_lut (.I0(n68198), .I1(n69484), .I2(n71241), .I3(n67807), 
            .O(n69695));   // verilog/motorControl.v(51[33:53])
    defparam i53520_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut (.I0(n69630), .I1(control_update), .I2(deadband[23]), 
            .I3(n356[23]), .O(n63914));
    defparam i1_4_lut.LUT_INIT = 16'h4c04;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n63914), .I1(n69695), .I2(n356[23]), 
            .I3(n47), .O(n62203));
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h0a22;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[15] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4566));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4567));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3843));   // verilog/motorControl.v(23[10] 30[6])
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4568));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4569));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[2]), 
            .I3(n51539), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4571));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n51539), .I0(GND_net), .I1(n1_adj_5099[2]), 
            .CO(n51540));
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[1]), 
            .I3(n51538), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4573));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4574));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4575));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4576));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n51538), .I0(GND_net), .I1(n1_adj_5099[1]), 
            .CO(n51539));
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4577));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5099[0]), 
            .CO(n51538));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n1[13]), .I3(n51458), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n51458), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n1[13]), .CO(n51459));
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4579));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4580));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n1[12]), .I3(n51457), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6242_20_lut (.I0(GND_net), .I1(n16118[17]), .I2(GND_net), 
            .I3(n51912), .O(n15358[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13909_3_lut (.I0(n379), .I1(n436[1]), .I2(n12030), .I3(GND_net), 
            .O(n28308));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4582));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30174_4_lut (.I0(PWMLimit[1]), .I1(n62203), .I2(n28308), 
            .I3(n12028), .O(n49[1]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30174_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6242_19_lut (.I0(GND_net), .I1(n16118[16]), .I2(GND_net), 
            .I3(n51911), .O(n15358[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4583));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13904_3_lut (.I0(n356[2]), .I1(n436[2]), .I2(n12030), .I3(GND_net), 
            .O(n28303));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30173_4_lut (.I0(PWMLimit[2]), .I1(n62203), .I2(n28303), 
            .I3(n12028), .O(n49[2]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30173_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6242_19 (.CI(n51911), .I0(n16118[16]), .I1(GND_net), 
            .CO(n51912));
    SB_LUT4 i13899_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n12030), .I3(GND_net), 
            .O(n28298));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30172_4_lut (.I0(PWMLimit[3]), .I1(n62203), .I2(n28298), 
            .I3(n12028), .O(n49[3]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30172_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6242_18_lut (.I0(GND_net), .I1(n16118[15]), .I2(GND_net), 
            .I3(n51910), .O(n15358[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13894_3_lut (.I0(n356[4]), .I1(n436[4]), .I2(n12030), .I3(GND_net), 
            .O(n28293));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13894_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_9_14 (.CI(n51457), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n1[12]), .CO(n51458));
    SB_LUT4 i30171_4_lut (.I0(PWMLimit[4]), .I1(n62203), .I2(n28293), 
            .I3(n12028), .O(n49[4]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30171_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n1[11]), .I3(n51456), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4585));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13889_3_lut (.I0(n356[5]), .I1(n436[5]), .I2(n12030), .I3(GND_net), 
            .O(n28288));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n49[0]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4586));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30170_4_lut (.I0(PWMLimit[5]), .I1(n62203), .I2(n28288), 
            .I3(n12028), .O(n49[5]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30170_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4587));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13884_3_lut (.I0(n356[6]), .I1(n436[6]), .I2(n12030), .I3(GND_net), 
            .O(n28283));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30169_4_lut (.I0(PWMLimit[6]), .I1(n62203), .I2(n28283), 
            .I3(n12028), .O(n49[6]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30169_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13879_3_lut (.I0(n356[7]), .I1(n436[7]), .I2(n12030), .I3(GND_net), 
            .O(n28278));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4589));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30168_4_lut (.I0(PWMLimit[7]), .I1(n62203), .I2(n28278), 
            .I3(n12028), .O(n49[7]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30168_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13874_3_lut (.I0(n356[8]), .I1(n436[8]), .I2(n12030), .I3(GND_net), 
            .O(n28273));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30167_4_lut (.I0(PWMLimit[8]), .I1(n62203), .I2(n28273), 
            .I3(n12028), .O(n49[8]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30167_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6242_18 (.CI(n51910), .I0(n16118[15]), .I1(GND_net), 
            .CO(n51911));
    SB_CARRY add_9_13 (.CI(n51456), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n1[11]), .CO(n51457));
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13869_3_lut (.I0(n356[9]), .I1(n436[9]), .I2(n12030), .I3(GND_net), 
            .O(n28268));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30166_4_lut (.I0(PWMLimit[9]), .I1(n62203), .I2(n28268), 
            .I3(n12028), .O(n49[9]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30166_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_6242_17_lut (.I0(GND_net), .I1(n16118[14]), .I2(GND_net), 
            .I3(n51909), .O(n15358[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4591));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6242_17 (.CI(n51909), .I0(n16118[14]), .I1(GND_net), 
            .CO(n51910));
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n1[10]), .I3(n51455), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13864_3_lut (.I0(n356[10]), .I1(n436[10]), .I2(n12030), .I3(GND_net), 
            .O(n28263));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4592));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6242_16_lut (.I0(GND_net), .I1(n16118[13]), .I2(n1108), 
            .I3(n51908), .O(n15358[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30165_4_lut (.I0(PWMLimit[10]), .I1(n62203), .I2(n28263), 
            .I3(n12028), .O(n49[10]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30165_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13859_3_lut (.I0(n356[11]), .I1(n436[11]), .I2(n12030), .I3(GND_net), 
            .O(n28258));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4593));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30164_4_lut (.I0(PWMLimit[11]), .I1(n62203), .I2(n28258), 
            .I3(n12028), .O(n49[11]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30164_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13854_3_lut (.I0(n356[12]), .I1(n436[12]), .I2(n12030), .I3(GND_net), 
            .O(n28253));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30163_4_lut (.I0(PWMLimit[12]), .I1(n62203), .I2(n28253), 
            .I3(n12028), .O(n49[12]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30163_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4595));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4596));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4597));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13849_3_lut (.I0(n356[13]), .I1(n436[13]), .I2(n12030), .I3(GND_net), 
            .O(n28248));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30162_4_lut (.I0(PWMLimit[13]), .I1(n62203), .I2(n28248), 
            .I3(n12028), .O(n49[13]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30162_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13844_3_lut (.I0(n356[14]), .I1(n436[14]), .I2(n12030), .I3(GND_net), 
            .O(n28243));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30161_4_lut (.I0(PWMLimit[14]), .I1(n62203), .I2(n28243), 
            .I3(n12028), .O(n49[14]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30161_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4598));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13839_3_lut (.I0(n356[15]), .I1(n436[15]), .I2(n12030), .I3(GND_net), 
            .O(n28238));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13839_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6242_16 (.CI(n51908), .I0(n16118[13]), .I1(n1108), .CO(n51909));
    SB_LUT4 add_6242_15_lut (.I0(GND_net), .I1(n16118[12]), .I2(n1035), 
            .I3(n51907), .O(n15358[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30160_4_lut (.I0(PWMLimit[15]), .I1(n62203), .I2(n28238), 
            .I3(n12028), .O(n49[15]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30160_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6242_15 (.CI(n51907), .I0(n16118[12]), .I1(n1035), .CO(n51908));
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4599));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4600));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4601));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13834_3_lut (.I0(n356[16]), .I1(n436[16]), .I2(n12030), .I3(GND_net), 
            .O(n28233));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30159_4_lut (.I0(PWMLimit[16]), .I1(n62203), .I2(n28233), 
            .I3(n12028), .O(n49[16]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30159_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13829_3_lut (.I0(n356[17]), .I1(n436[17]), .I2(n12030), .I3(GND_net), 
            .O(n28228));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6242_14_lut (.I0(GND_net), .I1(n16118[11]), .I2(n962), 
            .I3(n51906), .O(n15358[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_14 (.CI(n51906), .I0(n16118[11]), .I1(n962), .CO(n51907));
    SB_LUT4 add_6242_13_lut (.I0(GND_net), .I1(n16118[10]), .I2(n889), 
            .I3(n51905), .O(n15358[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_13 (.CI(n51905), .I0(n16118[10]), .I1(n889), .CO(n51906));
    SB_CARRY add_9_12 (.CI(n51455), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n1[10]), .CO(n51456));
    SB_LUT4 add_6242_12_lut (.I0(GND_net), .I1(n16118[9]), .I2(n816_adj_4602), 
            .I3(n51904), .O(n15358[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_12 (.CI(n51904), .I0(n16118[9]), .I1(n816_adj_4602), 
            .CO(n51905));
    SB_LUT4 add_6242_11_lut (.I0(GND_net), .I1(n16118[8]), .I2(n743_adj_4603), 
            .I3(n51903), .O(n15358[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n1[9]), .I3(n51454), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_11 (.CI(n51903), .I0(n16118[8]), .I1(n743_adj_4603), 
            .CO(n51904));
    SB_CARRY add_9_11 (.CI(n51454), .I0(\PID_CONTROLLER.integral [9]), .I1(n1[9]), 
            .CO(n51455));
    SB_LUT4 add_6242_10_lut (.I0(GND_net), .I1(n16118[7]), .I2(n670_adj_4605), 
            .I3(n51902), .O(n15358[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n1[8]), .I3(n51453), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30158_4_lut (.I0(PWMLimit[17]), .I1(n62203), .I2(n28228), 
            .I3(n12028), .O(n49[17]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30158_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6242_10 (.CI(n51902), .I0(n16118[7]), .I1(n670_adj_4605), 
            .CO(n51903));
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4606));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_10 (.CI(n51453), .I0(\PID_CONTROLLER.integral [8]), .I1(n1[8]), 
            .CO(n51454));
    SB_LUT4 add_6242_9_lut (.I0(GND_net), .I1(n16118[6]), .I2(n597_adj_4607), 
            .I3(n51901), .O(n15358[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_9 (.CI(n51901), .I0(n16118[6]), .I1(n597_adj_4607), 
            .CO(n51902));
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4608));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n1[7]), .I3(n51452), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_9 (.CI(n51452), .I0(\PID_CONTROLLER.integral [7]), .I1(n1[7]), 
            .CO(n51453));
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n1[6]), .I3(n51451), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_8 (.CI(n51451), .I0(\PID_CONTROLLER.integral [6]), .I1(n1[6]), 
            .CO(n51452));
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4610));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13824_3_lut (.I0(n356[18]), .I1(n436[18]), .I2(n12030), .I3(GND_net), 
            .O(n28223));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30157_4_lut (.I0(PWMLimit[18]), .I1(n62203), .I2(n28223), 
            .I3(n12028), .O(n49[18]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30157_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6242_8_lut (.I0(GND_net), .I1(n16118[5]), .I2(n524_adj_4611), 
            .I3(n51900), .O(n15358[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_8 (.CI(n51900), .I0(n16118[5]), .I1(n524_adj_4611), 
            .CO(n51901));
    SB_LUT4 add_6242_7_lut (.I0(GND_net), .I1(n16118[4]), .I2(n451_adj_4612), 
            .I3(n51899), .O(n15358[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n1[5]), .I3(n51450), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n136), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4613));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6242_7 (.CI(n51899), .I0(n16118[4]), .I1(n451_adj_4612), 
            .CO(n51900));
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4614));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6242_6_lut (.I0(GND_net), .I1(n16118[3]), .I2(n378_adj_4616), 
            .I3(n51898), .O(n15358[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_6 (.CI(n51898), .I0(n16118[3]), .I1(n378_adj_4616), 
            .CO(n51899));
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4617));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n356[20]), .I1(n436[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4618));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13819_3_lut (.I0(n356[19]), .I1(n436[19]), .I2(n12030), .I3(GND_net), 
            .O(n28218));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6242_5_lut (.I0(GND_net), .I1(n16118[2]), .I2(n305_adj_4619), 
            .I3(n51897), .O(n15358[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_5 (.CI(n51897), .I0(n16118[2]), .I1(n305_adj_4619), 
            .CO(n51898));
    SB_LUT4 add_6242_4_lut (.I0(GND_net), .I1(n16118[1]), .I2(n232_adj_4620), 
            .I3(n51896), .O(n15358[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n356[19]), .I1(n436[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4621));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n356[22]), .I1(n436[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4622));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n356[21]), .I1(n436[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4624));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4625));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n356[18]), .I1(n436[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4626));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30156_4_lut (.I0(PWMLimit[19]), .I1(n62203), .I2(n28218), 
            .I3(n12028), .O(n49[19]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30156_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4627));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n356[14]), .I1(n436[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4628));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_9_7 (.CI(n51450), .I0(\PID_CONTROLLER.integral [5]), .I1(n1[5]), 
            .CO(n51451));
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4629));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4630));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n356[15]), .I1(n436[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4631));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4632));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6242_4 (.CI(n51896), .I0(n16118[1]), .I1(n232_adj_4620), 
            .CO(n51897));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n1[4]), .I3(n51449), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13814_3_lut (.I0(n356[20]), .I1(n436[20]), .I2(n12030), .I3(GND_net), 
            .O(n28213));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4634));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4635));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n356[11]), .I1(n436[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4636));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30155_4_lut (.I0(PWMLimit[20]), .I1(n62203), .I2(n28213), 
            .I3(n12028), .O(n49[20]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30155_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n356[12]), .I1(n436[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4638));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6242_3_lut (.I0(GND_net), .I1(n16118[0]), .I2(n159_adj_4639), 
            .I3(n51895), .O(n15358[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6242_3 (.CI(n51895), .I0(n16118[0]), .I1(n159_adj_4639), 
            .CO(n51896));
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4640));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4641));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_6 (.CI(n51449), .I0(\PID_CONTROLLER.integral [4]), .I1(n1[4]), 
            .CO(n51450));
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n1[3]), .I3(n51448), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_5 (.CI(n51448), .I0(\PID_CONTROLLER.integral [3]), .I1(n1[3]), 
            .CO(n51449));
    SB_LUT4 i13809_3_lut (.I0(n356[21]), .I1(n436[21]), .I2(n12030), .I3(GND_net), 
            .O(n28208));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6242_2_lut (.I0(GND_net), .I1(n17_adj_4642), .I2(n86_adj_4643), 
            .I3(GND_net), .O(n15358[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6242_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30154_4_lut (.I0(PWMLimit[21]), .I1(n62203), .I2(n28208), 
            .I3(n12028), .O(n49[21]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30154_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4645));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n356[17]), .I1(n436[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4646));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4647));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4648));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36752_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[21] ), .I3(\Ki[1] ), 
            .O(n20670[0]));   // verilog/motorControl.v(50[27:38])
    defparam i36752_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4649));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13804_3_lut (.I0(n356[22]), .I1(n436[22]), .I2(n12030), .I3(GND_net), 
            .O(n28203));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4650));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n1[2]), .I3(n51447), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30153_4_lut (.I0(PWMLimit[22]), .I1(n62203), .I2(n28203), 
            .I3(n12028), .O(n49[22]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30153_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6242_2 (.CI(GND_net), .I0(n17_adj_4642), .I1(n86_adj_4643), 
            .CO(n51895));
    SB_LUT4 i36754_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[21] ), .I3(\Ki[1] ), 
            .O(n51027));   // verilog/motorControl.v(50[27:38])
    defparam i36754_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4651));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4652));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51361_4_lut (.I0(n21_adj_4647), .I1(n19_adj_4645), .I2(n17_adj_4640), 
            .I3(n9_adj_4635), .O(n67535));
    defparam i51361_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51346_4_lut (.I0(n27_adj_4652), .I1(n15_adj_4651), .I2(n13_adj_4648), 
            .I3(n11), .O(n67520));
    defparam i51346_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_4630), 
            .I3(GND_net), .O(n12_adj_4654));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6482_12_lut (.I0(GND_net), .I1(n19798[9]), .I2(n840), 
            .I3(n51675), .O(n19534[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n149), .I1(n130[6]), .I2(n13_adj_4648), 
            .I3(GND_net), .O(n10_adj_4655));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_4654), .I1(n130[17]), .I2(n35_adj_4629), 
            .I3(GND_net), .O(n30_adj_4656));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n356[16]), .I1(n436[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4657));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n356[5]), .I1(n436[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4658));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n356[6]), .I1(n436[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4659));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n356[7]), .I1(n436[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4660));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n356[13]), .I1(n436[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4661));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52298_4_lut (.I0(n13_adj_4648), .I1(n11), .I2(n9_adj_4635), 
            .I3(n67578), .O(n68472));
    defparam i52298_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n356[4]), .I1(n436[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4662));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52284_4_lut (.I0(n19_adj_4645), .I1(n17_adj_4640), .I2(n15_adj_4651), 
            .I3(n68472), .O(n68458));
    defparam i52284_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6482_11_lut (.I0(GND_net), .I1(n19798[8]), .I2(n767), 
            .I3(n51674), .O(n19534[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53396_4_lut (.I0(n25_adj_4617), .I1(n23_adj_4614), .I2(n21_adj_4647), 
            .I3(n68458), .O(n69571));
    defparam i53396_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n356[8]), .I1(n436[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4663));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4664));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13799_3_lut (.I0(n356[23]), .I1(n436[23]), .I2(n12030), .I3(GND_net), 
            .O(n28198));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30152_4_lut (.I0(PWMLimit[23]), .I1(n62203), .I2(n28198), 
            .I3(n12028), .O(n49[23]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i30152_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52776_4_lut (.I0(n31_adj_4627), .I1(n29_adj_4625), .I2(n27_adj_4652), 
            .I3(n69571), .O(n68951));
    defparam i52776_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n356[9]), .I1(n436[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4666));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6482_11 (.CI(n51674), .I0(n19798[8]), .I1(n767), .CO(n51675));
    SB_CARRY add_9_4 (.CI(n51447), .I0(\PID_CONTROLLER.integral [2]), .I1(n1[2]), 
            .CO(n51448));
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n1[1]), .I3(n51446), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4667));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4668));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36908_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[20] ), .I3(\Ki[1] ), 
            .O(n20653[0]));   // verilog/motorControl.v(50[27:38])
    defparam i36908_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36910_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[20] ), .I3(\Ki[1] ), 
            .O(n51191));   // verilog/motorControl.v(50[27:38])
    defparam i36910_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i53530_4_lut (.I0(n37_adj_4613), .I1(n35_adj_4629), .I2(n33_adj_4630), 
            .I3(n68951), .O(n69705));
    defparam i53530_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52790_3_lut (.I0(n6_adj_4669), .I1(n130[10]), .I2(n21_adj_4647), 
            .I3(GND_net), .O(n68965));   // verilog/motorControl.v(45[12:34])
    defparam i52790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4670));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_3 (.CI(n51446), .I0(\PID_CONTROLLER.integral [1]), .I1(n1[1]), 
            .CO(n51447));
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4671));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n356[10]), .I1(n436[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4672));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n1[0]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6482_10_lut (.I0(GND_net), .I1(n19798[7]), .I2(n694), 
            .I3(n51673), .O(n19534[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n1[0]), 
            .CO(n51446));
    SB_LUT4 i51539_4_lut (.I0(n21_adj_4672), .I1(n19_adj_4666), .I2(n17_adj_4663), 
            .I3(n9_adj_4662), .O(n67713));
    defparam i51539_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52791_3_lut (.I0(n68965), .I1(n130[11]), .I2(n23_adj_4614), 
            .I3(GND_net), .O(n68966));   // verilog/motorControl.v(45[12:34])
    defparam i52791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n51445), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_10 (.CI(n51673), .I0(n19798[7]), .I1(n694), .CO(n51674));
    SB_LUT4 add_6482_9_lut (.I0(GND_net), .I1(n19798[6]), .I2(n621), .I3(n51672), 
            .O(n19534[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_24_lut (.I0(n1[23]), .I1(n12570[21]), .I2(GND_net), 
            .I3(n52069), .O(n12063[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6482_9 (.CI(n51672), .I0(n19798[6]), .I1(n621), .CO(n51673));
    SB_LUT4 mult_16_add_1225_23_lut (.I0(GND_net), .I1(n12570[20]), .I2(GND_net), 
            .I3(n52068), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51533_4_lut (.I0(n27_adj_4661), .I1(n15_adj_4660), .I2(n13_adj_4659), 
            .I3(n11_adj_4658), .O(n67707));
    defparam i51533_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n436[7]), .I1(n436[16]), .I2(n33_adj_4657), 
            .I3(GND_net), .O(n12_adj_4673));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_4640), 
            .I3(GND_net), .O(n8_adj_4674));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16), .I1(n130[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4675));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n436[5]), .I1(n436[6]), .I2(n13_adj_4659), 
            .I3(GND_net), .O(n10_adj_4676));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12_adj_4673), .I1(n436[17]), .I2(n35_adj_4646), 
            .I3(GND_net), .O(n30_adj_4677));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4678));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51304_4_lut (.I0(n43), .I1(n25_adj_4617), .I2(n23_adj_4614), 
            .I3(n67535), .O(n67478));
    defparam i51304_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52986_4_lut (.I0(n24_adj_4675), .I1(n8_adj_4674), .I2(n45), 
            .I3(n67443), .O(n69161));   // verilog/motorControl.v(45[12:34])
    defparam i52986_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51994_3_lut (.I0(n68966), .I1(n130[12]), .I2(n25_adj_4617), 
            .I3(GND_net), .O(n68168));   // verilog/motorControl.v(45[12:34])
    defparam i51994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(n1_adj_5099[0]), .O(n4_adj_4679));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h8e0c;
    SB_LUT4 i52788_3_lut (.I0(n4_adj_4679), .I1(n130[13]), .I2(n27_adj_4652), 
            .I3(GND_net), .O(n68963));   // verilog/motorControl.v(45[12:34])
    defparam i52788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52789_3_lut (.I0(n68963), .I1(n130[14]), .I2(n29_adj_4625), 
            .I3(GND_net), .O(n68964));   // verilog/motorControl.v(45[12:34])
    defparam i52789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51329_4_lut (.I0(n33_adj_4630), .I1(n31_adj_4627), .I2(n29_adj_4625), 
            .I3(n67520), .O(n67503));
    defparam i51329_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52434_4_lut (.I0(n13_adj_4659), .I1(n11_adj_4658), .I2(n9_adj_4662), 
            .I3(n67729), .O(n68608));
    defparam i52434_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53195_4_lut (.I0(n30_adj_4656), .I1(n10_adj_4655), .I2(n35_adj_4629), 
            .I3(n67499), .O(n69370));   // verilog/motorControl.v(45[12:34])
    defparam i53195_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52428_4_lut (.I0(n19_adj_4666), .I1(n17_adj_4663), .I2(n15_adj_4660), 
            .I3(n68608), .O(n68602));
    defparam i52428_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53466_4_lut (.I0(n25_adj_4638), .I1(n23_adj_4636), .I2(n21_adj_4672), 
            .I3(n68602), .O(n69641));
    defparam i53466_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(n4_adj_4680), .I3(n20653[1]), .O(n20622[2]));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i52846_4_lut (.I0(n31_adj_4631), .I1(n29_adj_4628), .I2(n27_adj_4661), 
            .I3(n69641), .O(n69021));
    defparam i52846_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36959_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(n4_adj_4680), .I3(n20653[1]), .O(n6_adj_4681));   // verilog/motorControl.v(50[27:38])
    defparam i36959_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53567_4_lut (.I0(n37_adj_4626), .I1(n35_adj_4646), .I2(n33_adj_4657), 
            .I3(n69021), .O(n69742));
    defparam i53567_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36951_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(n51223), .I3(n20653[0]), .O(n4_adj_4680));   // verilog/motorControl.v(50[27:38])
    defparam i36951_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i51996_3_lut (.I0(n68964), .I1(n130[15]), .I2(n31_adj_4627), 
            .I3(GND_net), .O(n68170));   // verilog/motorControl.v(45[12:34])
    defparam i51996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53624_4_lut (.I0(n68170), .I1(n69370), .I2(n35_adj_4629), 
            .I3(n67503), .O(n69799));   // verilog/motorControl.v(45[12:34])
    defparam i53624_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53625_3_lut (.I0(n69799), .I1(n136), .I2(n37_adj_4613), .I3(GND_net), 
            .O(n69800));   // verilog/motorControl.v(45[12:34])
    defparam i53625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53540_3_lut (.I0(n69800), .I1(n130[19]), .I2(n39), .I3(GND_net), 
            .O(n69715));   // verilog/motorControl.v(45[12:34])
    defparam i53540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53074_3_lut (.I0(n6_adj_4682), .I1(n436[10]), .I2(n21_adj_4672), 
            .I3(GND_net), .O(n69249));   // verilog/motorControl.v(54[23:39])
    defparam i53074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51306_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69705), 
            .O(n67480));
    defparam i51306_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n436[9]), .I1(n436[21]), .I2(n43_adj_4624), 
            .I3(GND_net), .O(n16_adj_4683));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53303_4_lut (.I0(n68168), .I1(n69161), .I2(n45), .I3(n67478), 
            .O(n69478));   // verilog/motorControl.v(45[12:34])
    defparam i53303_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52002_3_lut (.I0(n69715), .I1(n130[20]), .I2(n41), .I3(GND_net), 
            .O(n68176));   // verilog/motorControl.v(45[12:34])
    defparam i52002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53514_4_lut (.I0(n68176), .I1(n69478), .I2(n45), .I3(n67480), 
            .O(n69689));   // verilog/motorControl.v(45[12:34])
    defparam i53514_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6482_8_lut (.I0(GND_net), .I1(n19798[5]), .I2(n548), .I3(n51671), 
            .O(n19534[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53515_3_lut (.I0(n69689), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(45[12:34])
    defparam i53515_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4684));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4685));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4686));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4687));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[3]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4688));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4689));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n436[4]), .I1(n436[8]), .I2(n17_adj_4663), 
            .I3(GND_net), .O(n8_adj_4690));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4691));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4693));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4694));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_4683), .I1(n436[22]), .I2(n45_adj_4622), 
            .I3(GND_net), .O(n24_adj_4695));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4697));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4698));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n149), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4699));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4700));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[4]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4702));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53075_3_lut (.I0(n69249), .I1(n436[11]), .I2(n23_adj_4636), 
            .I3(GND_net), .O(n69250));   // verilog/motorControl.v(54[23:39])
    defparam i53075_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_16_add_1225_23 (.CI(n52068), .I0(n12570[20]), .I1(GND_net), 
            .CO(n52069));
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4703));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_add_1225_22_lut (.I0(GND_net), .I1(n12570[19]), .I2(GND_net), 
            .I3(n52067), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51504_4_lut (.I0(n43_adj_4624), .I1(n25_adj_4638), .I2(n23_adj_4636), 
            .I3(n67713), .O(n67678));
    defparam i51504_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4704));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4705));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53004_4_lut (.I0(n24_adj_4695), .I1(n8_adj_4690), .I2(n45_adj_4622), 
            .I3(n67676), .O(n69179));   // verilog/motorControl.v(54[23:39])
    defparam i53004_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY mult_16_add_1225_22 (.CI(n52067), .I0(n12570[19]), .I1(GND_net), 
            .CO(n52068));
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[5]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52036_3_lut (.I0(n69250), .I1(n436[12]), .I2(n25_adj_4638), 
            .I3(GND_net), .O(n68210));   // verilog/motorControl.v(54[23:39])
    defparam i52036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[6]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[7]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[8]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[9]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6482_8 (.CI(n51671), .I0(n19798[5]), .I1(n548), .CO(n51672));
    SB_LUT4 add_6482_7_lut (.I0(GND_net), .I1(n19798[4]), .I2(n475), .I3(n51670), 
            .O(n19534[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n20622[2]), .I1(n6), .I2(n37023), .I3(\Ki[4] ), 
            .O(n20573[3]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h9666;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4711));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4713));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4714));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4715));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51226_4_lut (.I0(n21_adj_4715), .I1(n19_adj_4714), .I2(n17_adj_4713), 
            .I3(n9_adj_4705), .O(n67400));
    defparam i51226_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51195_4_lut (.I0(n27_adj_4704), .I1(n15_adj_4703), .I2(n13_adj_4702), 
            .I3(n11_adj_4699), .O(n67369));
    defparam i51195_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_25_i4_4_lut (.I0(n436[0]), .I1(n436[1]), .I2(n379), 
            .I3(n356[0]), .O(n4_adj_4717));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_16_add_1225_21_lut (.I0(GND_net), .I1(n12570[18]), .I2(GND_net), 
            .I3(n52066), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_4698), 
            .I3(GND_net), .O(n12_adj_4718));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_4702), 
            .I3(GND_net), .O(n10_adj_4719));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_16_add_1225_21 (.CI(n52066), .I0(n12570[18]), .I1(GND_net), 
            .CO(n52067));
    SB_LUT4 i53072_3_lut (.I0(n4_adj_4717), .I1(n436[13]), .I2(n27_adj_4661), 
            .I3(GND_net), .O(n69247));   // verilog/motorControl.v(54[23:39])
    defparam i53072_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6482_7 (.CI(n51670), .I0(n19798[4]), .I1(n475), .CO(n51671));
    SB_LUT4 i1_4_lut_adj_950 (.I0(n20670[0]), .I1(n51191), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3844[20] ), .O(n20653[1]));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_4718), .I1(n182[17]), .I2(n35_adj_4697), 
            .I3(GND_net), .O(n30_adj_4720));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n51444), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53073_3_lut (.I0(n69247), .I1(n436[14]), .I2(n29_adj_4628), 
            .I3(GND_net), .O(n69248));   // verilog/motorControl.v(54[23:39])
    defparam i53073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52131_4_lut (.I0(n13_adj_4702), .I1(n11_adj_4699), .I2(n9_adj_4705), 
            .I3(n67435), .O(n68305));
    defparam i52131_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_6482_6_lut (.I0(GND_net), .I1(n19798[3]), .I2(n402), .I3(n51669), 
            .O(n19534[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51524_4_lut (.I0(n33_adj_4657), .I1(n31_adj_4631), .I2(n29_adj_4628), 
            .I3(n67707), .O(n67698));
    defparam i51524_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4721));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_951 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3844[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3844[23] ), .O(n63894));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_952 (.I0(n37023), .I1(\Ki[4] ), .I2(\Ki[5] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3844[19] ), .O(n63898));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_953 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3844[20] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3844[21] ), .O(n63896));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h6ca0;
    SB_LUT4 i52117_4_lut (.I0(n19_adj_4714), .I1(n17_adj_4713), .I2(n15_adj_4703), 
            .I3(n68305), .O(n68291));
    defparam i52117_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4722));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4723));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_24 (.CI(n51444), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n51445));
    SB_LUT4 i1_3_lut_4_lut_adj_954 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(n51223), .I3(n20653[0]), .O(n20625));   // verilog/motorControl.v(50[27:38])
    defparam i1_3_lut_4_lut_adj_954.LUT_INIT = 16'h8778;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n63896), .I1(n51027), .I2(n63898), .I3(n63894), 
            .O(n63904));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i36921_4_lut (.I0(n20670[0]), .I1(\Ki[2] ), .I2(n51191), .I3(\PID_CONTROLLER.integral_23__N_3844[20] ), 
            .O(n4_adj_4724));   // verilog/motorControl.v(50[27:38])
    defparam i36921_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i37013_4_lut (.I0(n20622[2]), .I1(n37023), .I2(n6), .I3(\Ki[4] ), 
            .O(n8_adj_4725));   // verilog/motorControl.v(50[27:38])
    defparam i37013_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i53337_4_lut (.I0(n25_adj_4686), .I1(n23_adj_4688), .I2(n21_adj_4715), 
            .I3(n68291), .O(n69512));
    defparam i53337_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_956 (.I0(n6_adj_4681), .I1(n8_adj_4725), .I2(n4_adj_4724), 
            .I3(n63904), .O(n61143));   // verilog/motorControl.v(50[27:38])
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i52699_4_lut (.I0(n31_adj_4694), .I1(n29_adj_4693), .I2(n27_adj_4704), 
            .I3(n69512), .O(n68874));
    defparam i52699_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53506_4_lut (.I0(n37), .I1(n35_adj_4697), .I2(n33_adj_4698), 
            .I3(n68874), .O(n69681));
    defparam i53506_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_4689), 
            .I3(GND_net), .O(n16_adj_4727));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4728));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36938_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[20] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[19] ), .I3(\Ki[1] ), 
            .O(n20626));   // verilog/motorControl.v(50[27:38])
    defparam i36938_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36940_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[20] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3844[19] ), .I3(\Ki[1] ), 
            .O(n51223));   // verilog/motorControl.v(50[27:38])
    defparam i36940_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i52782_3_lut (.I0(n6_adj_4729), .I1(n182[10]), .I2(n21_adj_4715), 
            .I3(GND_net), .O(n68957));   // verilog/motorControl.v(47[21:44])
    defparam i52782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53436_4_lut (.I0(n30_adj_4677), .I1(n10_adj_4676), .I2(n35_adj_4646), 
            .I3(n67696), .O(n69611));   // verilog/motorControl.v(54[23:39])
    defparam i53436_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n51443), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52038_3_lut (.I0(n69248), .I1(n436[15]), .I2(n31_adj_4631), 
            .I3(GND_net), .O(n68212));   // verilog/motorControl.v(54[23:39])
    defparam i52038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[10]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[11]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4732));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52783_3_lut (.I0(n68957), .I1(n182[11]), .I2(n23_adj_4688), 
            .I3(GND_net), .O(n68958));   // verilog/motorControl.v(47[21:44])
    defparam i52783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4733));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4734));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[12]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_4713), 
            .I3(GND_net), .O(n8_adj_4736));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[13]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_4727), .I1(n182[22]), .I2(n45_adj_4687), 
            .I3(GND_net), .O(n24_adj_4738));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53642_4_lut (.I0(n68212), .I1(n69611), .I2(n35_adj_4646), 
            .I3(n67698), .O(n69817));   // verilog/motorControl.v(54[23:39])
    defparam i53642_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53643_3_lut (.I0(n69817), .I1(n436[18]), .I2(n37_adj_4626), 
            .I3(GND_net), .O(n69818));   // verilog/motorControl.v(54[23:39])
    defparam i53643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4739));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[14]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6482_6 (.CI(n51669), .I0(n19798[3]), .I1(n402), .CO(n51670));
    SB_LUT4 mult_16_add_1225_20_lut (.I0(GND_net), .I1(n12570[17]), .I2(GND_net), 
            .I3(n52065), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53606_3_lut (.I0(n69818), .I1(n436[19]), .I2(n39_adj_4621), 
            .I3(GND_net), .O(n69781));   // verilog/motorControl.v(54[23:39])
    defparam i53606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[15]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[16]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4743));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[17]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_8_add_2_23 (.CI(n51443), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n51444));
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51863_4_lut (.I0(n43_adj_4689), .I1(n25_adj_4686), .I2(n23_adj_4688), 
            .I3(n67400), .O(n68037));
    defparam i51863_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[18]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52992_4_lut (.I0(n24_adj_4738), .I1(n8_adj_4736), .I2(n45_adj_4687), 
            .I3(n68033), .O(n69167));   // verilog/motorControl.v(47[21:44])
    defparam i52992_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52004_3_lut (.I0(n68958), .I1(n182[12]), .I2(n25_adj_4686), 
            .I3(GND_net), .O(n68178));   // verilog/motorControl.v(47[21:44])
    defparam i52004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_4745));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51508_4_lut (.I0(n43_adj_4624), .I1(n41_adj_4618), .I2(n39_adj_4621), 
            .I3(n69742), .O(n67682));
    defparam i51508_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[19]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53313_4_lut (.I0(n68210), .I1(n69179), .I2(n45_adj_4622), 
            .I3(n67678), .O(n69488));   // verilog/motorControl.v(54[23:39])
    defparam i53313_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52044_3_lut (.I0(n69781), .I1(n436[20]), .I2(n41_adj_4618), 
            .I3(GND_net), .O(n68218));   // verilog/motorControl.v(54[23:39])
    defparam i52044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[20]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[21]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53249_3_lut (.I0(n4_adj_4745), .I1(n182[13]), .I2(n27_adj_4704), 
            .I3(GND_net), .O(n69424));   // verilog/motorControl.v(47[21:44])
    defparam i53249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4749));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[22]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53250_3_lut (.I0(n69424), .I1(n182[14]), .I2(n29_adj_4693), 
            .I3(GND_net), .O(n69425));   // verilog/motorControl.v(47[21:44])
    defparam i53250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51067_4_lut (.I0(n33_adj_4698), .I1(n31_adj_4694), .I2(n29_adj_4693), 
            .I3(n67369), .O(n67241));
    defparam i51067_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4750));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4751));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[23]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4752));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53542_4_lut (.I0(n30_adj_4720), .I1(n10_adj_4719), .I2(n35_adj_4697), 
            .I3(n67232), .O(n69717));   // verilog/motorControl.v(47[21:44])
    defparam i53542_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52989_3_lut (.I0(n69425), .I1(n182[15]), .I2(n31_adj_4694), 
            .I3(GND_net), .O(n69164));   // verilog/motorControl.v(47[21:44])
    defparam i52989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23001_1_lut (.I0(n356[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37361));   // verilog/motorControl.v(50[18:38])
    defparam i23001_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53688_4_lut (.I0(n69164), .I1(n69717), .I2(n35_adj_4697), 
            .I3(n67241), .O(n69863));   // verilog/motorControl.v(47[21:44])
    defparam i53688_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53689_3_lut (.I0(n69863), .I1(n188), .I2(n37), .I3(GND_net), 
            .O(n69864));   // verilog/motorControl.v(47[21:44])
    defparam i53689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53649_3_lut (.I0(n69864), .I1(n182[19]), .I2(n39_adj_4684), 
            .I3(GND_net), .O(n69824));   // verilog/motorControl.v(47[21:44])
    defparam i53649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[0]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4754));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53524_4_lut (.I0(n68218), .I1(n69488), .I2(n45_adj_4622), 
            .I3(n67682), .O(n69699));   // verilog/motorControl.v(54[23:39])
    defparam i53524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53525_3_lut (.I0(n69699), .I1(n356[23]), .I2(n436[23]), .I3(GND_net), 
            .O(n69700));   // verilog/motorControl.v(54[23:39])
    defparam i53525_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i6036_3_lut (.I0(control_update), .I1(n409), .I2(n69700), 
            .I3(GND_net), .O(n12030));   // verilog/motorControl.v(20[7:21])
    defparam i6036_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i51867_4_lut (.I0(n43_adj_4689), .I1(n41_adj_4685), .I2(n39_adj_4684), 
            .I3(n69681), .O(n68041));
    defparam i51867_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53516_4_lut (.I0(n68178), .I1(n69167), .I2(n45_adj_4687), 
            .I3(n68037), .O(n69691));   // verilog/motorControl.v(47[21:44])
    defparam i53516_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13754_3_lut (.I0(n356[0]), .I1(n436[0]), .I2(n12030), .I3(GND_net), 
            .O(n28153));   // verilog/motorControl.v(41[14] 61[8])
    defparam i13754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4755));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53598_3_lut (.I0(n69824), .I1(n182[20]), .I2(n41_adj_4685), 
            .I3(GND_net), .O(n40_adj_4756));   // verilog/motorControl.v(47[21:44])
    defparam i53598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n405_c));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53518_4_lut (.I0(n40_adj_4756), .I1(n69691), .I2(n45_adj_4687), 
            .I3(n68041), .O(n69693));   // verilog/motorControl.v(47[21:44])
    defparam i53518_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29682_4_lut (.I0(PWMLimit[0]), .I1(n62203), .I2(n28153), 
            .I3(n12028), .O(n49[0]));   // verilog/motorControl.v(41[14] 61[8])
    defparam i29682_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4757));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53519_3_lut (.I0(n69693), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(47[21:44])
    defparam i53519_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4759));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[14] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4760));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4762));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4763));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4764));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n51442), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4765));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4766));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4767));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4768));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4769));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4770));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[1]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4772));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4773));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4774));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4775));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4776));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4777));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4778));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4779));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4780));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4781));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[2]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4783));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4784));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4785));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_22 (.CI(n51442), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n51443));
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4786));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6482_5_lut (.I0(GND_net), .I1(n19798[2]), .I2(n329_adj_4787), 
            .I3(n51668), .O(n19534[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_5 (.CI(n51668), .I0(n19798[2]), .I1(n329_adj_4787), 
            .CO(n51669));
    SB_CARRY mult_16_add_1225_20 (.CI(n52065), .I0(n12570[17]), .I1(GND_net), 
            .CO(n52066));
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4788));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4789));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6482_4_lut (.I0(GND_net), .I1(n19798[1]), .I2(n256_adj_4790), 
            .I3(n51667), .O(n19534[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4791));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4792));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4793));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4794));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4795));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_19_lut (.I0(GND_net), .I1(n12570[16]), .I2(GND_net), 
            .I3(n52064), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6279_19_lut (.I0(GND_net), .I1(n16802[16]), .I2(GND_net), 
            .I3(n51880), .O(n16118[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4796));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n51441), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_19 (.CI(n52064), .I0(n12570[16]), .I1(GND_net), 
            .CO(n52065));
    SB_CARRY sub_8_add_2_21 (.CI(n51441), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n51442));
    SB_LUT4 mult_16_add_1225_18_lut (.I0(GND_net), .I1(n12570[15]), .I2(GND_net), 
            .I3(n52063), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[3]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6482_4 (.CI(n51667), .I0(n19798[1]), .I1(n256_adj_4790), 
            .CO(n51668));
    SB_CARRY mult_16_add_1225_18 (.CI(n52063), .I0(n12570[15]), .I1(GND_net), 
            .CO(n52064));
    SB_LUT4 add_6482_3_lut (.I0(GND_net), .I1(n19798[0]), .I2(n183_adj_4798), 
            .I3(n51666), .O(n19534[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4799));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6279_18_lut (.I0(GND_net), .I1(n16802[15]), .I2(GND_net), 
            .I3(n51879), .O(n16118[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4800));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6279_18 (.CI(n51879), .I0(n16802[15]), .I1(GND_net), 
            .CO(n51880));
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n51440), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[4]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[5]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4803));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6482_3 (.CI(n51666), .I0(n19798[0]), .I1(n183_adj_4798), 
            .CO(n51667));
    SB_LUT4 add_6482_2_lut (.I0(GND_net), .I1(n41_adj_4804), .I2(n110_adj_4805), 
            .I3(GND_net), .O(n19534[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6482_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6279_17_lut (.I0(GND_net), .I1(n16802[14]), .I2(GND_net), 
            .I3(n51878), .O(n16118[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6482_2 (.CI(GND_net), .I0(n41_adj_4804), .I1(n110_adj_4805), 
            .CO(n51666));
    SB_CARRY sub_8_add_2_20 (.CI(n51440), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n51441));
    SB_LUT4 mult_16_add_1225_17_lut (.I0(GND_net), .I1(n12570[14]), .I2(GND_net), 
            .I3(n52062), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[6]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n51439), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_17 (.CI(n52062), .I0(n12570[14]), .I1(GND_net), 
            .CO(n52063));
    SB_CARRY add_6279_17 (.CI(n51878), .I0(n16802[14]), .I1(GND_net), 
            .CO(n51879));
    SB_LUT4 mult_16_add_1225_16_lut (.I0(GND_net), .I1(n12570[13]), .I2(n1096_adj_4807), 
            .I3(n52061), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6279_16_lut (.I0(GND_net), .I1(n16802[13]), .I2(n1111_adj_4808), 
            .I3(n51877), .O(n16118[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6279_16 (.CI(n51877), .I0(n16802[13]), .I1(n1111_adj_4808), 
            .CO(n51878));
    SB_LUT4 add_6279_15_lut (.I0(GND_net), .I1(n16802[12]), .I2(n1038_adj_4809), 
            .I3(n51876), .O(n16118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_16 (.CI(n52061), .I0(n12570[13]), .I1(n1096_adj_4807), 
            .CO(n52062));
    SB_CARRY add_6279_15 (.CI(n51876), .I0(n16802[12]), .I1(n1038_adj_4809), 
            .CO(n51877));
    SB_CARRY sub_8_add_2_19 (.CI(n51439), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n51440));
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[7]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[8]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6279_14_lut (.I0(GND_net), .I1(n16802[11]), .I2(n965_adj_4812), 
            .I3(n51875), .O(n16118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[9]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_15_lut (.I0(GND_net), .I1(n12570[12]), .I2(n1023_adj_4814), 
            .I3(n52060), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[10]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6279_14 (.CI(n51875), .I0(n16802[11]), .I1(n965_adj_4812), 
            .CO(n51876));
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4816));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6279_13_lut (.I0(GND_net), .I1(n16802[10]), .I2(n892_adj_4817), 
            .I3(n51874), .O(n16118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6279_13 (.CI(n51874), .I0(n16802[10]), .I1(n892_adj_4817), 
            .CO(n51875));
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[11]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4819));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n51438), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4820));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_15 (.CI(n52060), .I0(n12570[12]), .I1(n1023_adj_4814), 
            .CO(n52061));
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[12]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6279_12_lut (.I0(GND_net), .I1(n16802[9]), .I2(n819_adj_4822), 
            .I3(n51873), .O(n16118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4823));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4824));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[13]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6279_12 (.CI(n51873), .I0(n16802[9]), .I1(n819_adj_4822), 
            .CO(n51874));
    SB_LUT4 add_6279_11_lut (.I0(GND_net), .I1(n16802[8]), .I2(n746_adj_4826), 
            .I3(n51872), .O(n16118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4827));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[14]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6279_11 (.CI(n51872), .I0(n16802[8]), .I1(n746_adj_4826), 
            .CO(n51873));
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_18 (.CI(n51438), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n51439));
    SB_LUT4 mult_16_add_1225_14_lut (.I0(GND_net), .I1(n12570[11]), .I2(n950_adj_4829), 
            .I3(n52059), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_14 (.CI(n52059), .I0(n12570[11]), .I1(n950_adj_4829), 
            .CO(n52060));
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[15]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4831));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[16]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_13_lut (.I0(GND_net), .I1(n12570[10]), .I2(n877_adj_4834), 
            .I3(n52058), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6279_10_lut (.I0(GND_net), .I1(n16802[7]), .I2(n673_adj_4835), 
            .I3(n51871), .O(n16118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4836));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6279_10 (.CI(n51871), .I0(n16802[7]), .I1(n673_adj_4835), 
            .CO(n51872));
    SB_CARRY mult_16_add_1225_13 (.CI(n52058), .I0(n12570[10]), .I1(n877_adj_4834), 
            .CO(n52059));
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n51437), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_17 (.CI(n51437), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n51438));
    SB_LUT4 mult_16_add_1225_12_lut (.I0(GND_net), .I1(n12570[9]), .I2(n804_adj_4837), 
            .I3(n52057), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_12 (.CI(n52057), .I0(n12570[9]), .I1(n804_adj_4837), 
            .CO(n52058));
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n51436), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_11_lut (.I0(GND_net), .I1(n12570[8]), .I2(n731_adj_4838), 
            .I3(n52056), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_16 (.CI(n51436), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n51437));
    SB_LUT4 add_6279_9_lut (.I0(GND_net), .I1(n16802[6]), .I2(n600_adj_4839), 
            .I3(n51870), .O(n16118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_11 (.CI(n52056), .I0(n12570[8]), .I1(n731_adj_4838), 
            .CO(n52057));
    SB_CARRY add_6279_9 (.CI(n51870), .I0(n16802[6]), .I1(n600_adj_4839), 
            .CO(n51871));
    SB_LUT4 add_6279_8_lut (.I0(GND_net), .I1(n16802[5]), .I2(n527_adj_4840), 
            .I3(n51869), .O(n16118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36984_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(\Ki[1] ), .I3(n37023), .O(n20573[0]));   // verilog/motorControl.v(50[27:38])
    defparam i36984_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4841));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4842));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1225_10_lut (.I0(GND_net), .I1(n12570[7]), .I2(n658_adj_4844), 
            .I3(n52055), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[17]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[18]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(n10), 
            .I3(n51435), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_15 (.CI(n51435), .I0(setpoint[13]), .I1(n10), 
            .CO(n51436));
    SB_CARRY add_6279_8 (.CI(n51869), .I0(n16802[5]), .I1(n527_adj_4840), 
            .CO(n51870));
    SB_LUT4 add_6279_7_lut (.I0(GND_net), .I1(n16802[4]), .I2(n454_adj_4848), 
            .I3(n51868), .O(n16118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4849));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_10 (.CI(n52055), .I0(n12570[7]), .I1(n658_adj_4844), 
            .CO(n52056));
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n51434), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6279_7 (.CI(n51868), .I0(n16802[4]), .I1(n454_adj_4848), 
            .CO(n51869));
    SB_LUT4 add_6279_6_lut (.I0(GND_net), .I1(n16802[3]), .I2(n381_adj_4850), 
            .I3(n51867), .O(n16118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6279_6 (.CI(n51867), .I0(n16802[3]), .I1(n381_adj_4850), 
            .CO(n51868));
    SB_LUT4 i36986_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[19] ), 
            .I2(\Ki[1] ), .I3(n37023), .O(n51273));   // verilog/motorControl.v(50[27:38])
    defparam i36986_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6279_5_lut (.I0(GND_net), .I1(n16802[2]), .I2(n308_adj_4851), 
            .I3(n51866), .O(n16118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4852));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4853));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6279_5 (.CI(n51866), .I0(n16802[2]), .I1(n308_adj_4851), 
            .CO(n51867));
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[19]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_14 (.CI(n51434), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n51435));
    SB_LUT4 mult_16_add_1225_9_lut (.I0(GND_net), .I1(n12570[6]), .I2(n585_adj_4855), 
            .I3(n52054), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[20]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n51433), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_13 (.CI(n51433), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n51434));
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4857));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_9 (.CI(n52054), .I0(n12570[6]), .I1(n585_adj_4855), 
            .CO(n52055));
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n51432), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_8_lut (.I0(GND_net), .I1(n12570[5]), .I2(n512_adj_4858), 
            .I3(n52053), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_8 (.CI(n52053), .I0(n12570[5]), .I1(n512_adj_4858), 
            .CO(n52054));
    SB_LUT4 mult_16_add_1225_7_lut (.I0(GND_net), .I1(n12570[4]), .I2(n439_adj_4859), 
            .I3(n52052), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[21]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6279_4_lut (.I0(GND_net), .I1(n16802[1]), .I2(n235_adj_4861), 
            .I3(n51865), .O(n16118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_7 (.CI(n52052), .I0(n12570[4]), .I1(n439_adj_4859), 
            .CO(n52053));
    SB_CARRY add_6279_4 (.CI(n51865), .I0(n16802[1]), .I1(n235_adj_4861), 
            .CO(n51866));
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[22]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5100[23]));   // verilog/motorControl.v(51[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_6_lut (.I0(GND_net), .I1(n12570[3]), .I2(n366_adj_4783), 
            .I3(n52051), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6279_3_lut (.I0(GND_net), .I1(n16802[0]), .I2(n162_adj_4774), 
            .I3(n51864), .O(n16118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6279_3 (.CI(n51864), .I0(n16802[0]), .I1(n162_adj_4774), 
            .CO(n51865));
    SB_LUT4 add_6279_2_lut (.I0(GND_net), .I1(n20_adj_4773), .I2(n89_adj_4772), 
            .I3(GND_net), .O(n16118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6279_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6279_2 (.CI(GND_net), .I0(n20_adj_4773), .I1(n89_adj_4772), 
            .CO(n51864));
    SB_CARRY sub_8_add_2_12 (.CI(n51432), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n51433));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n51431), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_10_lut (.I0(GND_net), .I1(n20278[7]), .I2(n700_adj_4760), 
            .I3(n51863), .O(n20117[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4864));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6531_9_lut (.I0(GND_net), .I1(n20278[6]), .I2(n627_adj_4608), 
            .I3(n51862), .O(n20117[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_9 (.CI(n51862), .I0(n20278[6]), .I1(n627_adj_4608), 
            .CO(n51863));
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[0]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6531_8_lut (.I0(GND_net), .I1(n20278[5]), .I2(n554_adj_4606), 
            .I3(n51861), .O(n20117[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_11 (.CI(n51431), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n51432));
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n51430), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_10 (.CI(n51430), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n51431));
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_6 (.CI(n52051), .I0(n12570[3]), .I1(n366_adj_4783), 
            .CO(n52052));
    SB_LUT4 i51261_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n67435));   // verilog/motorControl.v(47[21:44])
    defparam i51261_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6531_8 (.CI(n51861), .I0(n20278[5]), .I1(n554_adj_4606), 
            .CO(n51862));
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n51429), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_9 (.CI(n51429), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n51430));
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n51428), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_adj_4729));   // verilog/motorControl.v(47[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_add_1225_5_lut (.I0(GND_net), .I1(n12570[2]), .I2(n293_adj_4600), 
            .I3(n52050), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_5 (.CI(n52050), .I0(n12570[2]), .I1(n293_adj_4600), 
            .CO(n52051));
    SB_LUT4 add_6531_7_lut (.I0(GND_net), .I1(n20278[4]), .I2(n481_adj_4599), 
            .I3(n51860), .O(n20117[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1225_4_lut (.I0(GND_net), .I1(n12570[1]), .I2(n220_adj_4597), 
            .I3(n52049), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4867));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_8 (.CI(n51428), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n51429));
    SB_CARRY add_6531_7 (.CI(n51860), .I0(n20278[4]), .I1(n481_adj_4599), 
            .CO(n51861));
    SB_LUT4 add_6531_6_lut (.I0(GND_net), .I1(n20278[3]), .I2(n408_adj_4595), 
            .I3(n51859), .O(n20117[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[1]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[2]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[3]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n306[0]));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1225_4 (.CI(n52049), .I0(n12570[1]), .I1(n220_adj_4597), 
            .CO(n52050));
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6531_6 (.CI(n51859), .I0(n20278[3]), .I1(n408_adj_4595), 
            .CO(n51860));
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[4]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_add_1225_3_lut (.I0(GND_net), .I1(n12570[0]), .I2(n147_adj_4593), 
            .I3(n52048), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1225_3 (.CI(n52048), .I0(n12570[0]), .I1(n147_adj_4593), 
            .CO(n52049));
    SB_LUT4 add_6531_5_lut (.I0(GND_net), .I1(n20278[2]), .I2(n335_adj_4592), 
            .I3(n51858), .O(n20117[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[5]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[6]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6531_5 (.CI(n51858), .I0(n20278[2]), .I1(n335_adj_4592), 
            .CO(n51859));
    SB_LUT4 add_6531_4_lut (.I0(GND_net), .I1(n20278[1]), .I2(n262_adj_4591), 
            .I3(n51857), .O(n20117[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[7]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[8]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4877));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n20598[2]), .I1(n6_adj_4878), .I2(\Kp[4] ), 
            .I3(n1[18]), .O(n20538[3]));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_957.LUT_INIT = 16'h9666;
    SB_CARRY add_6531_4 (.CI(n51857), .I0(n20278[1]), .I1(n262_adj_4591), 
            .CO(n51858));
    SB_LUT4 mult_16_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4571), .I2(n74_adj_4569), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n51427), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4879));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4880));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204_adj_4881));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36969_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n20662[0]));   // verilog/motorControl.v(50[18:24])
    defparam i36969_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_4882));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4883));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4861));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4884));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_958 (.I0(\Kp[4] ), .I1(\Kp[5] ), .I2(n1[19]), 
            .I3(n1[18]), .O(n63928));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_3_lut (.I0(\Kp[3] ), .I1(n63928), .I2(n1[20]), .I3(GND_net), 
            .O(n63930));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i142_2_lut (.I0(\Kp[2] ), .I1(n1[21]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_959 (.I0(\Kp[1] ), .I1(n210), .I2(n1[22]), .I3(n63930), 
            .O(n63934));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h936c;
    SB_LUT4 i36971_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n51257));   // verilog/motorControl.v(50[18:24])
    defparam i36971_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_960 (.I0(n51257), .I1(\Kp[0] ), .I2(n63934), 
            .I3(n1[23]), .O(n63938));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_960.LUT_INIT = 16'h695a;
    SB_LUT4 i36891_4_lut (.I0(n20598[2]), .I1(\Kp[4] ), .I2(n6_adj_4878), 
            .I3(n1[18]), .O(n8_adj_4885));   // verilog/motorControl.v(50[18:24])
    defparam i36891_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_961 (.I0(n6_adj_4886), .I1(n8_adj_4885), .I2(n4_adj_4887), 
            .I3(n63938), .O(n61880));   // verilog/motorControl.v(50[18:24])
    defparam i1_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 add_6531_3_lut (.I0(GND_net), .I1(n20278[0]), .I2(n189), .I3(n51856), 
            .O(n20117[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n51427), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n51428));
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4888));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4889));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6531_3 (.CI(n51856), .I0(n20278[0]), .I1(n189), .CO(n51857));
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4859));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n51426), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_2_lut (.I0(GND_net), .I1(n47_adj_4566), .I2(n116), 
            .I3(GND_net), .O(n20117[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[9]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4891));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4892));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4893));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[10]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4895));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[11]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4897));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[12]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4858));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_6 (.CI(n51426), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n51427));
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4899));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[13]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_16_add_1225_2 (.CI(GND_net), .I0(n5_adj_4571), .I1(n74_adj_4569), 
            .CO(n52048));
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4901));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[14]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4903));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4904));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[15]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4906));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4907));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4908));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[16]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[17]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6531_2 (.CI(GND_net), .I0(n47_adj_4566), .I1(n116), .CO(n51856));
    SB_LUT4 sub_8_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(\motor_state[3] ), 
            .I3(n51425), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4911));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[18]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[19]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[20]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_8_add_2_5 (.CI(n51425), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n51426));
    SB_LUT4 sub_8_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(\motor_state[2] ), 
            .I3(n51424), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[21]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4916));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[22]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_4 (.CI(n51424), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n51425));
    SB_LUT4 sub_8_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(\motor_state[1] ), 
            .I3(n51423), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4855));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4851));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4850));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5101[23]));   // verilog/motorControl.v(55[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20591_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n34987));   // verilog/motorControl.v(41[14] 61[8])
    defparam i20591_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4919));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(GND_net), .O(n6_adj_4682));   // verilog/motorControl.v(54[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY sub_8_add_2_3 (.CI(n51423), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n51424));
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4848));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51555_3_lut_4_lut (.I0(n356[3]), .I1(n436[3]), .I2(n436[2]), 
            .I3(n356[2]), .O(n67729));   // verilog/motorControl.v(54[23:39])
    defparam i51555_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4920));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(\motor_state[0] ), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4921));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4844));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4922));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4923));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4924));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4925));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4840));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4926));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4927));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4928));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4929));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4839));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4930));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4838));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4931));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4837));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4932));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4933));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4934));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4935));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4936));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4937));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4938));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4939));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n51423));
    SB_LUT4 add_6314_18_lut (.I0(GND_net), .I1(n17414[15]), .I2(GND_net), 
            .I3(n51842), .O(n16802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6314_17_lut (.I0(GND_net), .I1(n17414[14]), .I2(GND_net), 
            .I3(n51841), .O(n16802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_17 (.CI(n51841), .I0(n17414[14]), .I1(GND_net), 
            .CO(n51842));
    SB_LUT4 add_6314_16_lut (.I0(GND_net), .I1(n17414[13]), .I2(n1114_adj_4940), 
            .I3(n51840), .O(n16802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4941));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4942));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4943));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4944));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4945));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4946));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4947));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4948));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4949));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4950));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4951));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4952));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4953));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4954));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4835));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4834));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_16 (.CI(n51840), .I0(n17414[13]), .I1(n1114_adj_4940), 
            .CO(n51841));
    SB_LUT4 add_6314_15_lut (.I0(GND_net), .I1(n17414[12]), .I2(n1041_adj_4955), 
            .I3(n51839), .O(n16802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_15 (.CI(n51839), .I0(n17414[12]), .I1(n1041_adj_4955), 
            .CO(n51840));
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4956));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4957));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4829));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6314_14_lut (.I0(GND_net), .I1(n17414[11]), .I2(n968_adj_4958), 
            .I3(n51838), .O(n16802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4959));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4826));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4960));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4822));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_14 (.CI(n51838), .I0(n17414[11]), .I1(n968_adj_4958), 
            .CO(n51839));
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4961));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6314_13_lut (.I0(GND_net), .I1(n17414[10]), .I2(n895_adj_4962), 
            .I3(n51837), .O(n16802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_13 (.CI(n51837), .I0(n17414[10]), .I1(n895_adj_4962), 
            .CO(n51838));
    SB_LUT4 add_6314_12_lut (.I0(GND_net), .I1(n17414[9]), .I2(n822_adj_4963), 
            .I3(n51836), .O(n16802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4964));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51404_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n67578));   // verilog/motorControl.v(45[12:34])
    defparam i51404_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4965));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4966));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4967));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4968));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4969));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4970));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4971));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4972));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_12 (.CI(n51836), .I0(n17414[9]), .I1(n822_adj_4963), 
            .CO(n51837));
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4973));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4974));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6314_11_lut (.I0(GND_net), .I1(n17414[8]), .I2(n749_adj_4975), 
            .I3(n51835), .O(n16802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_11 (.CI(n51835), .I0(n17414[8]), .I1(n749_adj_4975), 
            .CO(n51836));
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4976));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4977));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4978));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4979));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4980));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4981));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_4669));   // verilog/motorControl.v(45[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_6314_10_lut (.I0(GND_net), .I1(n17414[7]), .I2(n676_adj_4982), 
            .I3(n51834), .O(n16802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_10 (.CI(n51834), .I0(n17414[7]), .I1(n676_adj_4982), 
            .CO(n51835));
    SB_LUT4 add_6314_9_lut (.I0(GND_net), .I1(n17414[6]), .I2(n603_adj_4983), 
            .I3(n51833), .O(n16802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_9 (.CI(n51833), .I0(n17414[6]), .I1(n603_adj_4983), 
            .CO(n51834));
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4817));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4814));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6314_8_lut (.I0(GND_net), .I1(n17414[5]), .I2(n530_adj_4984), 
            .I3(n51832), .O(n16802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_8 (.CI(n51832), .I0(n17414[5]), .I1(n530_adj_4984), 
            .CO(n51833));
    SB_LUT4 add_6314_7_lut (.I0(GND_net), .I1(n17414[4]), .I2(n457_adj_4985), 
            .I3(n51831), .O(n16802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4812));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4809));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4808));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_7 (.CI(n51831), .I0(n17414[4]), .I1(n457_adj_4985), 
            .CO(n51832));
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4807));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6314_6_lut (.I0(GND_net), .I1(n17414[3]), .I2(n384_adj_4986), 
            .I3(n51830), .O(n16802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4805));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4804));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4798));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4790));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4787));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_6 (.CI(n51830), .I0(n17414[3]), .I1(n384_adj_4986), 
            .CO(n51831));
    SB_LUT4 add_6314_5_lut (.I0(GND_net), .I1(n17414[2]), .I2(n311_adj_4987), 
            .I3(n51829), .O(n16802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n30012), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_5 (.CI(n51829), .I0(n17414[2]), .I1(n311_adj_4987), 
            .CO(n51830));
    SB_LUT4 add_6314_4_lut (.I0(GND_net), .I1(n17414[1]), .I2(n238_adj_4988), 
            .I3(n51828), .O(n16802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_4 (.CI(n51828), .I0(n17414[1]), .I1(n238_adj_4988), 
            .CO(n51829));
    SB_DFFSR counter_2053__i0 (.Q(counter[0]), .C(clk16MHz), .D(n51[0]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i31 (.Q(counter[31]), .C(clk16MHz), .D(n51[31]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i30 (.Q(counter[30]), .C(clk16MHz), .D(n51[30]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i29 (.Q(counter[29]), .C(clk16MHz), .D(n51[29]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i28 (.Q(counter[28]), .C(clk16MHz), .D(n51[28]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i27 (.Q(counter[27]), .C(clk16MHz), .D(n51[27]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i26 (.Q(counter[26]), .C(clk16MHz), .D(n51[26]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i25 (.Q(counter[25]), .C(clk16MHz), .D(n51[25]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i24 (.Q(counter[24]), .C(clk16MHz), .D(n51[24]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i23 (.Q(counter[23]), .C(clk16MHz), .D(n51[23]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i22 (.Q(counter[22]), .C(clk16MHz), .D(n51[22]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i21 (.Q(counter[21]), .C(clk16MHz), .D(n51[21]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i20 (.Q(counter[20]), .C(clk16MHz), .D(n51[20]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i19 (.Q(counter[19]), .C(clk16MHz), .D(n51[19]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i18 (.Q(counter[18]), .C(clk16MHz), .D(n51[18]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i17 (.Q(counter[17]), .C(clk16MHz), .D(n51[17]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i16 (.Q(counter[16]), .C(clk16MHz), .D(n51[16]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i15 (.Q(counter[15]), .C(clk16MHz), .D(n51[15]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i14 (.Q(counter[14]), .C(clk16MHz), .D(n51[14]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i13 (.Q(counter[13]), .C(clk16MHz), .D(n51[13]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i12 (.Q(counter[12]), .C(clk16MHz), .D(n51[12]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i11 (.Q(counter[11]), .C(clk16MHz), .D(n51[11]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i10 (.Q(counter[10]), .C(clk16MHz), .D(n51[10]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i9 (.Q(counter[9]), .C(clk16MHz), .D(n51[9]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i8 (.Q(counter[8]), .C(clk16MHz), .D(n51[8]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i7 (.Q(counter[7]), .C(clk16MHz), .D(n51[7]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i6 (.Q(counter[6]), .C(clk16MHz), .D(n51[6]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i5 (.Q(counter[5]), .C(clk16MHz), .D(n51[5]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i4 (.Q(counter[4]), .C(clk16MHz), .D(n51[4]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i3 (.Q(counter[3]), .C(clk16MHz), .D(n51[3]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i2 (.Q(counter[2]), .C(clk16MHz), .D(n51[2]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_2053__i1 (.Q(counter[1]), .C(clk16MHz), .D(n51[1]), 
            .R(counter_31__N_3843));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 add_6314_3_lut (.I0(GND_net), .I1(n17414[0]), .I2(n165_adj_5015), 
            .I3(n51827), .O(n16802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6314_3 (.CI(n51827), .I0(n17414[0]), .I1(n165_adj_5015), 
            .CO(n51828));
    SB_LUT4 add_6113_23_lut (.I0(GND_net), .I1(n13590[20]), .I2(GND_net), 
            .I3(n52029), .O(n12570[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6314_2_lut (.I0(GND_net), .I1(n23_adj_5016), .I2(n92_adj_5017), 
            .I3(GND_net), .O(n16802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6314_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6314_2 (.CI(GND_net), .I0(n23_adj_5016), .I1(n92_adj_5017), 
            .CO(n51827));
    SB_LUT4 add_6113_22_lut (.I0(GND_net), .I1(n13590[19]), .I2(GND_net), 
            .I3(n52028), .O(n12570[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_22 (.CI(n52028), .I0(n13590[19]), .I1(GND_net), 
            .CO(n52029));
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4643));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6113_21_lut (.I0(GND_net), .I1(n13590[18]), .I2(GND_net), 
            .I3(n52027), .O(n12570[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_21 (.CI(n52027), .I0(n13590[18]), .I1(GND_net), 
            .CO(n52028));
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30827), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30826), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30825), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30824), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30823), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30822), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30821), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30820), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30819), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30818), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30817), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30816), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30815), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30814), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30813), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4642));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30812), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30811), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30810), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30809), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30808), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30807), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30806), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30805), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4639));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6113_20_lut (.I0(GND_net), .I1(n13590[17]), .I2(GND_net), 
            .I3(n52026), .O(n12570[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_20 (.CI(n52026), .I0(n13590[17]), .I1(GND_net), 
            .CO(n52027));
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_5018));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6113_19_lut (.I0(GND_net), .I1(n13590[16]), .I2(GND_net), 
            .I3(n52025), .O(n12570[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n49[23]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n49[22]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4620));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n49[21]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n49[20]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n49[19]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n49[18]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n49[17]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n49[16]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n49[15]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n49[14]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n49[13]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n49[12]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n49[11]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n49[10]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n49[9]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n49[8]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n49[7]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n49[6]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n49[5]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n49[4]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n49[3]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n49[2]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n49[1]), .R(reset));   // verilog/motorControl.v(41[14] 61[8])
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4619));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4616));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4612));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4611));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4607));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4605));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4603));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4602));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3844[23] ), 
            .I1(n13105[21]), .I2(GND_net), .I3(n53109), .O(n12598[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n13105[20]), .I2(GND_net), 
            .I3(n53108), .O(n306[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_23 (.CI(n53108), .I0(n13105[20]), .I1(GND_net), 
            .CO(n53109));
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n13105[19]), .I2(GND_net), 
            .I3(n53107), .O(n306[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n53107), .I0(n13105[19]), .I1(GND_net), 
            .CO(n53108));
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n13105[18]), .I2(GND_net), 
            .I3(n53106), .O(n306[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n53106), .I0(n13105[18]), .I1(GND_net), 
            .CO(n53107));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n13105[17]), .I2(GND_net), 
            .I3(n53105), .O(n306[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n53105), .I0(n13105[17]), .I1(GND_net), 
            .CO(n53106));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n13105[16]), .I2(GND_net), 
            .I3(n53104), .O(n306[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n53104), .I0(n13105[16]), .I1(GND_net), 
            .CO(n53105));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n13105[15]), .I2(GND_net), 
            .I3(n53103), .O(n306[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n53103), .I0(n13105[15]), .I1(GND_net), 
            .CO(n53104));
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n13105[14]), .I2(GND_net), 
            .I3(n53102), .O(n306[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_17 (.CI(n53102), .I0(n13105[14]), .I1(GND_net), 
            .CO(n53103));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n13105[13]), .I2(n1096), 
            .I3(n53101), .O(n306[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n53101), .I0(n13105[13]), .I1(n1096), 
            .CO(n53102));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n13105[12]), .I2(n1023), 
            .I3(n53100), .O(n306[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_15 (.CI(n53100), .I0(n13105[12]), .I1(n1023), 
            .CO(n53101));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n13105[11]), .I2(n950), 
            .I3(n53099), .O(n306[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_14 (.CI(n53099), .I0(n13105[11]), .I1(n950), 
            .CO(n53100));
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n13105[10]), .I2(n877), 
            .I3(n53098), .O(n306[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_13 (.CI(n53098), .I0(n13105[10]), .I1(n877), 
            .CO(n53099));
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n13105[9]), .I2(n804), 
            .I3(n53097), .O(n306[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_12 (.CI(n53097), .I0(n13105[9]), .I1(n804), 
            .CO(n53098));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n13105[8]), .I2(n731), 
            .I3(n53096), .O(n306[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_11 (.CI(n53096), .I0(n13105[8]), .I1(n731), 
            .CO(n53097));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n13105[7]), .I2(n658), 
            .I3(n53095), .O(n306[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_10 (.CI(n53095), .I0(n13105[7]), .I1(n658), 
            .CO(n53096));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n13105[6]), .I2(n585), 
            .I3(n53094), .O(n306[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_9 (.CI(n53094), .I0(n13105[6]), .I1(n585), 
            .CO(n53095));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n13105[5]), .I2(n512), 
            .I3(n53093), .O(n306[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_8 (.CI(n53093), .I0(n13105[5]), .I1(n512), 
            .CO(n53094));
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n13105[4]), .I2(n439), 
            .I3(n53092), .O(n306[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_7 (.CI(n53092), .I0(n13105[4]), .I1(n439), 
            .CO(n53093));
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n13105[3]), .I2(n366_adj_4560), 
            .I3(n53091), .O(n306[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n53091), .I0(n13105[3]), .I1(n366_adj_4560), 
            .CO(n53092));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n13105[2]), .I2(n293), 
            .I3(n53090), .O(n306[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n53090), .I0(n13105[2]), .I1(n293), 
            .CO(n53091));
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n13105[1]), .I2(n220), 
            .I3(n53089), .O(n306[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_4 (.CI(n53089), .I0(n13105[1]), .I1(n220), 
            .CO(n53090));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n13105[0]), .I2(n147), 
            .I3(n53088), .O(n306[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_3 (.CI(n53088), .I0(n13105[0]), .I1(n147), 
            .CO(n53089));
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n306[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n53088));
    SB_LUT4 add_6139_23_lut (.I0(GND_net), .I1(n14074[20]), .I2(GND_net), 
            .I3(n53087), .O(n13105[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6139_22_lut (.I0(GND_net), .I1(n14074[19]), .I2(GND_net), 
            .I3(n53086), .O(n13105[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_22 (.CI(n53086), .I0(n14074[19]), .I1(GND_net), 
            .CO(n53087));
    SB_LUT4 add_6139_21_lut (.I0(GND_net), .I1(n14074[18]), .I2(GND_net), 
            .I3(n53085), .O(n13105[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_21 (.CI(n53085), .I0(n14074[18]), .I1(GND_net), 
            .CO(n53086));
    SB_LUT4 add_6139_20_lut (.I0(GND_net), .I1(n14074[17]), .I2(GND_net), 
            .I3(n53084), .O(n13105[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_20 (.CI(n53084), .I0(n14074[17]), .I1(GND_net), 
            .CO(n53085));
    SB_LUT4 add_6139_19_lut (.I0(GND_net), .I1(n14074[16]), .I2(GND_net), 
            .I3(n53083), .O(n13105[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_19 (.CI(n53083), .I0(n14074[16]), .I1(GND_net), 
            .CO(n53084));
    SB_LUT4 add_6139_18_lut (.I0(GND_net), .I1(n14074[15]), .I2(GND_net), 
            .I3(n53082), .O(n13105[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_18 (.CI(n53082), .I0(n14074[15]), .I1(GND_net), 
            .CO(n53083));
    SB_LUT4 add_6139_17_lut (.I0(GND_net), .I1(n14074[14]), .I2(GND_net), 
            .I3(n53081), .O(n13105[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_17 (.CI(n53081), .I0(n14074[14]), .I1(GND_net), 
            .CO(n53082));
    SB_LUT4 add_6139_16_lut (.I0(GND_net), .I1(n14074[13]), .I2(n1099), 
            .I3(n53080), .O(n13105[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_16 (.CI(n53080), .I0(n14074[13]), .I1(n1099), .CO(n53081));
    SB_LUT4 add_6139_15_lut (.I0(GND_net), .I1(n14074[12]), .I2(n1026), 
            .I3(n53079), .O(n13105[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_15 (.CI(n53079), .I0(n14074[12]), .I1(n1026), .CO(n53080));
    SB_LUT4 add_6139_14_lut (.I0(GND_net), .I1(n14074[11]), .I2(n953_adj_5024), 
            .I3(n53078), .O(n13105[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_14 (.CI(n53078), .I0(n14074[11]), .I1(n953_adj_5024), 
            .CO(n53079));
    SB_LUT4 add_6139_13_lut (.I0(GND_net), .I1(n14074[10]), .I2(n880_adj_5025), 
            .I3(n53077), .O(n13105[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_13 (.CI(n53077), .I0(n14074[10]), .I1(n880_adj_5025), 
            .CO(n53078));
    SB_LUT4 add_6139_12_lut (.I0(GND_net), .I1(n14074[9]), .I2(n807_adj_5026), 
            .I3(n53076), .O(n13105[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[0]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6139_12 (.CI(n53076), .I0(n14074[9]), .I1(n807_adj_5026), 
            .CO(n53077));
    SB_LUT4 add_6139_11_lut (.I0(GND_net), .I1(n14074[8]), .I2(n734_adj_5027), 
            .I3(n53075), .O(n13105[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_11 (.CI(n53075), .I0(n14074[8]), .I1(n734_adj_5027), 
            .CO(n53076));
    SB_LUT4 add_6139_10_lut (.I0(GND_net), .I1(n14074[7]), .I2(n661_adj_5028), 
            .I3(n53074), .O(n13105[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_10 (.CI(n53074), .I0(n14074[7]), .I1(n661_adj_5028), 
            .CO(n53075));
    SB_LUT4 add_6139_9_lut (.I0(GND_net), .I1(n14074[6]), .I2(n588_adj_5029), 
            .I3(n53073), .O(n13105[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_9 (.CI(n53073), .I0(n14074[6]), .I1(n588_adj_5029), 
            .CO(n53074));
    SB_CARRY add_6113_19 (.CI(n52025), .I0(n13590[16]), .I1(GND_net), 
            .CO(n52026));
    SB_LUT4 add_6139_8_lut (.I0(GND_net), .I1(n14074[5]), .I2(n515_adj_5030), 
            .I3(n53072), .O(n13105[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_8 (.CI(n53072), .I0(n14074[5]), .I1(n515_adj_5030), 
            .CO(n53073));
    SB_LUT4 add_6139_7_lut (.I0(GND_net), .I1(n14074[4]), .I2(n442_adj_5031), 
            .I3(n53071), .O(n13105[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_7 (.CI(n53071), .I0(n14074[4]), .I1(n442_adj_5031), 
            .CO(n53072));
    SB_LUT4 add_6139_6_lut (.I0(GND_net), .I1(n14074[3]), .I2(n369_adj_5032), 
            .I3(n53070), .O(n13105[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_6 (.CI(n53070), .I0(n14074[3]), .I1(n369_adj_5032), 
            .CO(n53071));
    SB_LUT4 add_6139_5_lut (.I0(GND_net), .I1(n14074[2]), .I2(n296_adj_5033), 
            .I3(n53069), .O(n13105[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_5 (.CI(n53069), .I0(n14074[2]), .I1(n296_adj_5033), 
            .CO(n53070));
    SB_LUT4 add_6139_4_lut (.I0(GND_net), .I1(n14074[1]), .I2(n223_adj_5034), 
            .I3(n53068), .O(n13105[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_4 (.CI(n53068), .I0(n14074[1]), .I1(n223_adj_5034), 
            .CO(n53069));
    SB_LUT4 add_6139_3_lut (.I0(GND_net), .I1(n14074[0]), .I2(n150_adj_5035), 
            .I3(n53067), .O(n13105[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[1]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5099[2]));   // verilog/motorControl.v(48[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6139_3 (.CI(n53067), .I0(n14074[0]), .I1(n150_adj_5035), 
            .CO(n53068));
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_5036));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_6139_2_lut (.I0(GND_net), .I1(n8_adj_5037), .I2(n77_adj_5038), 
            .I3(GND_net), .O(n13105[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_3_lut (.I0(counter[5]), .I1(counter[2]), .I2(counter[0]), 
            .I3(GND_net), .O(n11_adj_5039));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(counter[19]), .I1(counter[28]), .I2(counter[27]), 
            .I3(GND_net), .O(n62077));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2825_4_lut (.I0(n11_adj_5039), .I1(counter[8]), .I2(counter[7]), 
            .I3(n12_adj_5036), .O(n18_adj_5040));
    defparam i2825_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_5041));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_4_lut (.I0(counter[24]), .I1(counter[30]), .I2(counter[29]), 
            .I3(n62077), .O(n16_adj_5042));
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_962 (.I0(counter[23]), .I1(counter[12]), .I2(n10_adj_5041), 
            .I3(n18_adj_5040), .O(n15_adj_5043));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'heaaa;
    SB_LUT4 i10_4_lut (.I0(counter[21]), .I1(counter[18]), .I2(counter[22]), 
            .I3(counter[26]), .O(n24_adj_5044));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(counter[17]), .I1(counter[20]), .I2(counter[16]), 
            .I3(counter[14]), .O(n23_adj_5045));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_6139_2 (.CI(GND_net), .I0(n8_adj_5037), .I1(n77_adj_5038), 
            .CO(n53067));
    SB_LUT4 add_6182_22_lut (.I0(GND_net), .I1(n14958[19]), .I2(GND_net), 
            .I3(n53066), .O(n14074[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6182_21_lut (.I0(GND_net), .I1(n14958[18]), .I2(GND_net), 
            .I3(n53065), .O(n14074[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut (.I0(counter[15]), .I1(n15_adj_5043), .I2(counter[25]), 
            .I3(n16_adj_5042), .O(n25_adj_5046));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29752_4_lut (.I0(n25_adj_5046), .I1(counter[31]), .I2(n23_adj_5045), 
            .I3(n24_adj_5044), .O(counter_31__N_3843));   // verilog/motorControl.v(26[8:41])
    defparam i29752_4_lut.LUT_INIT = 16'h3332;
    SB_CARRY add_6182_21 (.CI(n53065), .I0(n14958[18]), .I1(GND_net), 
            .CO(n53066));
    SB_LUT4 add_6182_20_lut (.I0(GND_net), .I1(n14958[17]), .I2(GND_net), 
            .I3(n53064), .O(n14074[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_20 (.CI(n53064), .I0(n14958[17]), .I1(GND_net), 
            .CO(n53065));
    SB_LUT4 add_6182_19_lut (.I0(GND_net), .I1(n14958[16]), .I2(GND_net), 
            .I3(n53063), .O(n14074[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_19 (.CI(n53063), .I0(n14958[16]), .I1(GND_net), 
            .CO(n53064));
    SB_LUT4 add_6182_18_lut (.I0(GND_net), .I1(n14958[15]), .I2(GND_net), 
            .I3(n53062), .O(n14074[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_18 (.CI(n53062), .I0(n14958[15]), .I1(GND_net), 
            .CO(n53063));
    SB_LUT4 add_6182_17_lut (.I0(GND_net), .I1(n14958[14]), .I2(GND_net), 
            .I3(n53061), .O(n14074[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_17 (.CI(n53061), .I0(n14958[14]), .I1(GND_net), 
            .CO(n53062));
    SB_LUT4 add_6113_18_lut (.I0(GND_net), .I1(n13590[15]), .I2(GND_net), 
            .I3(n52024), .O(n12570[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_18 (.CI(n52024), .I0(n13590[15]), .I1(GND_net), 
            .CO(n52025));
    SB_LUT4 add_6182_16_lut (.I0(GND_net), .I1(n14958[13]), .I2(n1102_adj_5047), 
            .I3(n53060), .O(n14074[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_16 (.CI(n53060), .I0(n14958[13]), .I1(n1102_adj_5047), 
            .CO(n53061));
    SB_LUT4 add_6182_15_lut (.I0(GND_net), .I1(n14958[12]), .I2(n1029_adj_5048), 
            .I3(n53059), .O(n14074[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[23] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6182_15 (.CI(n53059), .I0(n14958[12]), .I1(n1029_adj_5048), 
            .CO(n53060));
    SB_LUT4 add_6182_14_lut (.I0(GND_net), .I1(n14958[11]), .I2(n956_adj_5049), 
            .I3(n53058), .O(n14074[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_14 (.CI(n53058), .I0(n14958[11]), .I1(n956_adj_5049), 
            .CO(n53059));
    SB_LUT4 add_6182_13_lut (.I0(GND_net), .I1(n14958[10]), .I2(n883_adj_5050), 
            .I3(n53057), .O(n14074[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_13 (.CI(n53057), .I0(n14958[10]), .I1(n883_adj_5050), 
            .CO(n53058));
    SB_LUT4 add_6182_12_lut (.I0(GND_net), .I1(n14958[9]), .I2(n810_adj_5051), 
            .I3(n53056), .O(n14074[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_12 (.CI(n53056), .I0(n14958[9]), .I1(n810_adj_5051), 
            .CO(n53057));
    SB_LUT4 add_6182_11_lut (.I0(GND_net), .I1(n14958[8]), .I2(n737_adj_5052), 
            .I3(n53055), .O(n14074[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n12063[0]), .I2(n12598[0]), 
            .I3(n51491), .O(n356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_11 (.CI(n53055), .I0(n14958[8]), .I1(n737_adj_5052), 
            .CO(n53056));
    SB_LUT4 add_6182_10_lut (.I0(GND_net), .I1(n14958[7]), .I2(n664_adj_5053), 
            .I3(n53054), .O(n14074[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6182_10 (.CI(n53054), .I0(n14958[7]), .I1(n664_adj_5053), 
            .CO(n53055));
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6182_9_lut (.I0(GND_net), .I1(n14958[6]), .I2(n591_adj_5054), 
            .I3(n53053), .O(n14074[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_9 (.CI(n53053), .I0(n14958[6]), .I1(n591_adj_5054), 
            .CO(n53054));
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[22] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[21] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6182_8_lut (.I0(GND_net), .I1(n14958[5]), .I2(n518_adj_5056), 
            .I3(n53052), .O(n14074[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_8 (.CI(n53052), .I0(n14958[5]), .I1(n518_adj_5056), 
            .CO(n53053));
    SB_LUT4 add_6182_7_lut (.I0(GND_net), .I1(n14958[4]), .I2(n445_adj_5018), 
            .I3(n53051), .O(n14074[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_7 (.CI(n53051), .I0(n14958[4]), .I1(n445_adj_5018), 
            .CO(n53052));
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[20] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2053_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n52733), .O(n51[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n52732), .O(n51[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_32 (.CI(n52732), .I0(GND_net), .I1(counter[30]), 
            .CO(n52733));
    SB_LUT4 counter_2053_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n52731), .O(n51[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_31 (.CI(n52731), .I0(GND_net), .I1(counter[29]), 
            .CO(n52732));
    SB_LUT4 counter_2053_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n52730), .O(n51[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6182_6_lut (.I0(GND_net), .I1(n14958[3]), .I2(n372_adj_4981), 
            .I3(n53050), .O(n14074[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_6 (.CI(n53050), .I0(n14958[3]), .I1(n372_adj_4981), 
            .CO(n53051));
    SB_CARRY counter_2053_add_4_30 (.CI(n52730), .I0(GND_net), .I1(counter[28]), 
            .CO(n52731));
    SB_LUT4 counter_2053_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n52729), .O(n51[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_17_lut (.I0(GND_net), .I1(n13590[14]), .I2(GND_net), 
            .I3(n52023), .O(n12570[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_17 (.CI(n52023), .I0(n13590[14]), .I1(GND_net), 
            .CO(n52024));
    SB_LUT4 add_6113_16_lut (.I0(GND_net), .I1(n13590[13]), .I2(n1099_adj_4921), 
            .I3(n52022), .O(n12570[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_29 (.CI(n52729), .I0(GND_net), .I1(counter[27]), 
            .CO(n52730));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n306[22]), 
            .I3(n51490), .O(n356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_24 (.CI(n51490), .I0(n257[22]), .I1(n306[22]), .CO(n51491));
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n207[19]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6182_5_lut (.I0(GND_net), .I1(n14958[2]), .I2(n299_adj_4919), 
            .I3(n53049), .O(n14074[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n52728), .O(n51[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_28 (.CI(n52728), .I0(GND_net), .I1(counter[26]), 
            .CO(n52729));
    SB_LUT4 mux_15_i20_3_lut (.I0(n207[19]), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[19] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6182_5 (.CI(n53049), .I0(n14958[2]), .I1(n299_adj_4919), 
            .CO(n53050));
    SB_LUT4 add_6182_4_lut (.I0(GND_net), .I1(n14958[1]), .I2(n226), .I3(n53048), 
            .O(n14074[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_4 (.CI(n53048), .I0(n14958[1]), .I1(n226), .CO(n53049));
    SB_LUT4 add_6182_3_lut (.I0(GND_net), .I1(n14958[0]), .I2(n153_adj_4824), 
            .I3(n53047), .O(n14074[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_16 (.CI(n52022), .I0(n13590[13]), .I1(n1099_adj_4921), 
            .CO(n52023));
    SB_CARRY add_6182_3 (.CI(n53047), .I0(n14958[0]), .I1(n153_adj_4824), 
            .CO(n53048));
    SB_LUT4 counter_2053_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n52727), .O(n51[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6182_2_lut (.I0(GND_net), .I1(n11_adj_4819), .I2(n80), 
            .I3(GND_net), .O(n14074[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6182_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n306[21]), 
            .I3(n51489), .O(n356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6182_2 (.CI(GND_net), .I0(n11_adj_4819), .I1(n80), .CO(n53047));
    SB_LUT4 add_6503_11_lut (.I0(GND_net), .I1(n20018[8]), .I2(n770_adj_4796), 
            .I3(n53046), .O(n19798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6503_10_lut (.I0(GND_net), .I1(n20018[7]), .I2(n697_adj_4786), 
            .I3(n53045), .O(n19798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_23 (.CI(n51489), .I0(n257[21]), .I1(n306[21]), .CO(n51490));
    SB_CARRY add_6503_10 (.CI(n53045), .I0(n20018[7]), .I1(n697_adj_4786), 
            .CO(n53046));
    SB_LUT4 add_6503_9_lut (.I0(GND_net), .I1(n20018[6]), .I2(n624_adj_4784), 
            .I3(n53044), .O(n19798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_9 (.CI(n53044), .I0(n20018[6]), .I1(n624_adj_4784), 
            .CO(n53045));
    SB_LUT4 add_6113_15_lut (.I0(GND_net), .I1(n13590[12]), .I2(n1026_adj_4776), 
            .I3(n52021), .O(n12570[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_27 (.CI(n52727), .I0(GND_net), .I1(counter[25]), 
            .CO(n52728));
    SB_LUT4 counter_2053_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n52726), .O(n51[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6503_8_lut (.I0(GND_net), .I1(n20018[5]), .I2(n551_adj_4764), 
            .I3(n53043), .O(n19798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_15 (.CI(n52021), .I0(n13590[12]), .I1(n1026_adj_4776), 
            .CO(n52022));
    SB_CARRY add_6503_8 (.CI(n53043), .I0(n20018[5]), .I1(n551_adj_4764), 
            .CO(n53044));
    SB_LUT4 add_6503_7_lut (.I0(GND_net), .I1(n20018[4]), .I2(n478_adj_4761), 
            .I3(n53042), .O(n19798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_7 (.CI(n53042), .I0(n20018[4]), .I1(n478_adj_4761), 
            .CO(n53043));
    SB_LUT4 add_6503_6_lut (.I0(GND_net), .I1(n20018[3]), .I2(n405_adj_4757), 
            .I3(n53041), .O(n19798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_6 (.CI(n53041), .I0(n20018[3]), .I1(n405_adj_4757), 
            .CO(n53042));
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n306[20]), 
            .I3(n51488), .O(n356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_14_lut (.I0(GND_net), .I1(n13590[11]), .I2(n953), 
            .I3(n52020), .O(n12570[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_14 (.CI(n52020), .I0(n13590[11]), .I1(n953), .CO(n52021));
    SB_LUT4 add_6503_5_lut (.I0(GND_net), .I1(n20018[2]), .I2(n332), .I3(n53040), 
            .O(n19798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_17_lut (.I0(GND_net), .I1(n17958[14]), .I2(GND_net), 
            .I3(n51814), .O(n17414[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_5 (.CI(n53040), .I0(n20018[2]), .I1(n332), .CO(n53041));
    SB_CARRY add_18_22 (.CI(n51488), .I0(n257[20]), .I1(n306[20]), .CO(n51489));
    SB_LUT4 add_6347_16_lut (.I0(GND_net), .I1(n17958[13]), .I2(n1117_adj_4739), 
            .I3(n51813), .O(n17414[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n306[19]), 
            .I3(n51487), .O(n356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_16 (.CI(n51813), .I0(n17958[13]), .I1(n1117_adj_4739), 
            .CO(n51814));
    SB_LUT4 add_6347_15_lut (.I0(GND_net), .I1(n17958[12]), .I2(n1044_adj_4732), 
            .I3(n51812), .O(n17414[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6503_4_lut (.I0(GND_net), .I1(n20018[1]), .I2(n259), .I3(n53039), 
            .O(n19798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_4 (.CI(n53039), .I0(n20018[1]), .I1(n259), .CO(n53040));
    SB_LUT4 add_6503_3_lut (.I0(GND_net), .I1(n20018[0]), .I2(n186_adj_4728), 
            .I3(n53038), .O(n19798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_3 (.CI(n53038), .I0(n20018[0]), .I1(n186_adj_4728), 
            .CO(n53039));
    SB_LUT4 add_6503_2_lut (.I0(GND_net), .I1(n44_adj_4723), .I2(n113_adj_4722), 
            .I3(GND_net), .O(n19798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_13_lut (.I0(GND_net), .I1(n13590[10]), .I2(n880), 
            .I3(n52019), .O(n12570[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6503_2 (.CI(GND_net), .I0(n44_adj_4723), .I1(n113_adj_4722), 
            .CO(n53038));
    SB_LUT4 add_6223_21_lut (.I0(GND_net), .I1(n15757[18]), .I2(GND_net), 
            .I3(n53037), .O(n14958[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6223_20_lut (.I0(GND_net), .I1(n15757[17]), .I2(GND_net), 
            .I3(n53036), .O(n14958[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_13 (.CI(n52019), .I0(n13590[10]), .I1(n880), .CO(n52020));
    SB_CARRY add_6223_20 (.CI(n53036), .I0(n15757[17]), .I1(GND_net), 
            .CO(n53037));
    SB_LUT4 add_6223_19_lut (.I0(GND_net), .I1(n15757[16]), .I2(GND_net), 
            .I3(n53035), .O(n14958[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_15 (.CI(n51812), .I0(n17958[12]), .I1(n1044_adj_4732), 
            .CO(n51813));
    SB_CARRY add_6223_19 (.CI(n53035), .I0(n15757[16]), .I1(GND_net), 
            .CO(n53036));
    SB_LUT4 add_6347_14_lut (.I0(GND_net), .I1(n17958[11]), .I2(n971_adj_4721), 
            .I3(n51811), .O(n17414[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6223_18_lut (.I0(GND_net), .I1(n15757[15]), .I2(GND_net), 
            .I3(n53034), .O(n14958[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_18 (.CI(n53034), .I0(n15757[15]), .I1(GND_net), 
            .CO(n53035));
    SB_LUT4 add_6223_17_lut (.I0(GND_net), .I1(n15757[14]), .I2(GND_net), 
            .I3(n53033), .O(n14958[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_17 (.CI(n53033), .I0(n15757[14]), .I1(GND_net), 
            .CO(n53034));
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n207[17]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6113_12_lut (.I0(GND_net), .I1(n13590[9]), .I2(n807), 
            .I3(n52018), .O(n12570[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_14 (.CI(n51811), .I0(n17958[11]), .I1(n971_adj_4721), 
            .CO(n51812));
    SB_LUT4 add_6223_16_lut (.I0(GND_net), .I1(n15757[13]), .I2(n1105), 
            .I3(n53032), .O(n14958[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_16 (.CI(n53032), .I0(n15757[13]), .I1(n1105), .CO(n53033));
    SB_LUT4 mux_15_i18_3_lut (.I0(n207[17]), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[17] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6347_13_lut (.I0(GND_net), .I1(n17958[10]), .I2(n898_adj_4691), 
            .I3(n51810), .O(n17414[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6223_15_lut (.I0(GND_net), .I1(n15757[12]), .I2(n1032), 
            .I3(n53031), .O(n14958[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_26 (.CI(n52726), .I0(GND_net), .I1(counter[24]), 
            .CO(n52727));
    SB_LUT4 counter_2053_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n52725), .O(n51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_15 (.CI(n53031), .I0(n15757[12]), .I1(n1032), .CO(n53032));
    SB_LUT4 add_6223_14_lut (.I0(GND_net), .I1(n15757[11]), .I2(n959), 
            .I3(n53030), .O(n14958[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6223_14 (.CI(n53030), .I0(n15757[11]), .I1(n959), .CO(n53031));
    SB_CARRY add_6347_13 (.CI(n51810), .I0(n17958[10]), .I1(n898_adj_4691), 
            .CO(n51811));
    SB_LUT4 add_6223_13_lut (.I0(GND_net), .I1(n15757[10]), .I2(n886), 
            .I3(n53029), .O(n14958[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_25 (.CI(n52725), .I0(GND_net), .I1(counter[23]), 
            .CO(n52726));
    SB_CARRY add_6223_13 (.CI(n53029), .I0(n15757[10]), .I1(n886), .CO(n53030));
    SB_LUT4 add_6223_12_lut (.I0(GND_net), .I1(n15757[9]), .I2(n813), 
            .I3(n53028), .O(n14958[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_12 (.CI(n53028), .I0(n15757[9]), .I1(n813), .CO(n53029));
    SB_LUT4 add_6223_11_lut (.I0(GND_net), .I1(n15757[8]), .I2(n740), 
            .I3(n53027), .O(n14958[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[16] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6113_12 (.CI(n52018), .I0(n13590[9]), .I1(n807), .CO(n52019));
    SB_LUT4 add_6113_11_lut (.I0(GND_net), .I1(n13590[8]), .I2(n734), 
            .I3(n52017), .O(n12570[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_12_lut (.I0(GND_net), .I1(n17958[9]), .I2(n825_adj_4678), 
            .I3(n51809), .O(n17414[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_11 (.CI(n53027), .I0(n15757[8]), .I1(n740), .CO(n53028));
    SB_LUT4 add_6223_10_lut (.I0(GND_net), .I1(n15757[7]), .I2(n667), 
            .I3(n53026), .O(n14958[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_10 (.CI(n53026), .I0(n15757[7]), .I1(n667), .CO(n53027));
    SB_LUT4 counter_2053_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n52724), .O(n51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6223_9_lut (.I0(GND_net), .I1(n15757[6]), .I2(n594), .I3(n53025), 
            .O(n14958[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_9 (.CI(n53025), .I0(n15757[6]), .I1(n594), .CO(n53026));
    SB_LUT4 add_6223_8_lut (.I0(GND_net), .I1(n15757[5]), .I2(n521), .I3(n53024), 
            .O(n14958[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_12 (.CI(n51809), .I0(n17958[9]), .I1(n825_adj_4678), 
            .CO(n51810));
    SB_CARRY add_6113_11 (.CI(n52017), .I0(n13590[8]), .I1(n734), .CO(n52018));
    SB_CARRY add_6223_8 (.CI(n53024), .I0(n15757[5]), .I1(n521), .CO(n53025));
    SB_CARRY add_18_21 (.CI(n51487), .I0(n257[19]), .I1(n306[19]), .CO(n51488));
    SB_LUT4 add_6223_7_lut (.I0(GND_net), .I1(n15757[4]), .I2(n448_adj_4671), 
            .I3(n53023), .O(n14958[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_7 (.CI(n53023), .I0(n15757[4]), .I1(n448_adj_4671), 
            .CO(n53024));
    SB_LUT4 add_6223_6_lut (.I0(GND_net), .I1(n15757[3]), .I2(n375_adj_4670), 
            .I3(n53022), .O(n14958[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_6 (.CI(n53022), .I0(n15757[3]), .I1(n375_adj_4670), 
            .CO(n53023));
    SB_LUT4 add_6113_10_lut (.I0(GND_net), .I1(n13590[7]), .I2(n661), 
            .I3(n52016), .O(n12570[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6223_5_lut (.I0(GND_net), .I1(n15757[2]), .I2(n302), .I3(n53021), 
            .O(n14958[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_24 (.CI(n52724), .I0(GND_net), .I1(counter[22]), 
            .CO(n52725));
    SB_CARRY add_6223_5 (.CI(n53021), .I0(n15757[2]), .I1(n302), .CO(n53022));
    SB_LUT4 add_6223_4_lut (.I0(GND_net), .I1(n15757[1]), .I2(n229), .I3(n53020), 
            .O(n14958[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n52723), .O(n51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_4 (.CI(n53020), .I0(n15757[1]), .I1(n229), .CO(n53021));
    SB_LUT4 add_6223_3_lut (.I0(GND_net), .I1(n15757[0]), .I2(n156), .I3(n53019), 
            .O(n14958[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_10 (.CI(n52016), .I0(n13590[7]), .I1(n661), .CO(n52017));
    SB_LUT4 add_6347_11_lut (.I0(GND_net), .I1(n17958[8]), .I2(n752_adj_4668), 
            .I3(n51808), .O(n17414[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_3 (.CI(n53019), .I0(n15757[0]), .I1(n156), .CO(n53020));
    SB_LUT4 add_6223_2_lut (.I0(GND_net), .I1(n14_adj_4667), .I2(n83), 
            .I3(GND_net), .O(n14958[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6223_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6223_2 (.CI(GND_net), .I0(n14_adj_4667), .I1(n83), .CO(n53019));
    SB_LUT4 add_6261_20_lut (.I0(GND_net), .I1(n16478[17]), .I2(GND_net), 
            .I3(n53018), .O(n15757[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_23 (.CI(n52723), .I0(GND_net), .I1(counter[21]), 
            .CO(n52724));
    SB_LUT4 counter_2053_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n52722), .O(n51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6261_19_lut (.I0(GND_net), .I1(n16478[16]), .I2(GND_net), 
            .I3(n53017), .O(n15757[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_19 (.CI(n53017), .I0(n16478[16]), .I1(GND_net), 
            .CO(n53018));
    SB_LUT4 add_6261_18_lut (.I0(GND_net), .I1(n16478[15]), .I2(GND_net), 
            .I3(n53016), .O(n15757[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_18 (.CI(n53016), .I0(n16478[15]), .I1(GND_net), 
            .CO(n53017));
    SB_CARRY add_6347_11 (.CI(n51808), .I0(n17958[8]), .I1(n752_adj_4668), 
            .CO(n51809));
    SB_LUT4 add_6347_10_lut (.I0(GND_net), .I1(n17958[7]), .I2(n679_adj_4664), 
            .I3(n51807), .O(n17414[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6261_17_lut (.I0(GND_net), .I1(n16478[14]), .I2(GND_net), 
            .I3(n53015), .O(n15757[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_22 (.CI(n52722), .I0(GND_net), .I1(counter[20]), 
            .CO(n52723));
    SB_LUT4 add_6113_9_lut (.I0(GND_net), .I1(n13590[6]), .I2(n588), .I3(n52015), 
            .O(n12570[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n52721), .O(n51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_9 (.CI(n52015), .I0(n13590[6]), .I1(n588), .CO(n52016));
    SB_CARRY add_6261_17 (.CI(n53015), .I0(n16478[14]), .I1(GND_net), 
            .CO(n53016));
    SB_LUT4 add_6261_16_lut (.I0(GND_net), .I1(n16478[13]), .I2(n1108_adj_4650), 
            .I3(n53014), .O(n15757[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_8_lut (.I0(GND_net), .I1(n13590[5]), .I2(n515), .I3(n52014), 
            .O(n12570[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_8 (.CI(n52014), .I0(n13590[5]), .I1(n515), .CO(n52015));
    SB_CARRY counter_2053_add_4_21 (.CI(n52721), .I0(GND_net), .I1(counter[19]), 
            .CO(n52722));
    SB_LUT4 add_6113_7_lut (.I0(GND_net), .I1(n13590[4]), .I2(n442_adj_4649), 
            .I3(n52013), .O(n12570[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_16 (.CI(n53014), .I0(n16478[13]), .I1(n1108_adj_4650), 
            .CO(n53015));
    SB_LUT4 add_6261_15_lut (.I0(GND_net), .I1(n16478[12]), .I2(n1035_adj_4641), 
            .I3(n53013), .O(n15757[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_7 (.CI(n52013), .I0(n13590[4]), .I1(n442_adj_4649), 
            .CO(n52014));
    SB_CARRY add_6261_15 (.CI(n53013), .I0(n16478[12]), .I1(n1035_adj_4641), 
            .CO(n53014));
    SB_CARRY add_6347_10 (.CI(n51807), .I0(n17958[7]), .I1(n679_adj_4664), 
            .CO(n51808));
    SB_LUT4 counter_2053_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n52720), .O(n51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6261_14_lut (.I0(GND_net), .I1(n16478[11]), .I2(n962_adj_4634), 
            .I3(n53012), .O(n15757[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_9_lut (.I0(GND_net), .I1(n17958[6]), .I2(n606_adj_4632), 
            .I3(n51806), .O(n17414[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_6_lut (.I0(GND_net), .I1(n13590[3]), .I2(n369_adj_4615), 
            .I3(n52012), .O(n12570[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_20 (.CI(n52720), .I0(GND_net), .I1(counter[18]), 
            .CO(n52721));
    SB_CARRY add_6261_14 (.CI(n53012), .I0(n16478[11]), .I1(n962_adj_4634), 
            .CO(n53013));
    SB_LUT4 add_6261_13_lut (.I0(GND_net), .I1(n16478[10]), .I2(n889_adj_4610), 
            .I3(n53011), .O(n15757[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_9 (.CI(n51806), .I0(n17958[6]), .I1(n606_adj_4632), 
            .CO(n51807));
    SB_LUT4 counter_2053_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n52719), .O(n51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_19 (.CI(n52719), .I0(GND_net), .I1(counter[17]), 
            .CO(n52720));
    SB_CARRY add_6261_13 (.CI(n53011), .I0(n16478[10]), .I1(n889_adj_4610), 
            .CO(n53012));
    SB_LUT4 add_6261_12_lut (.I0(GND_net), .I1(n16478[9]), .I2(n816), 
            .I3(n53010), .O(n15757[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n306[18]), 
            .I3(n51486), .O(n356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_8_lut (.I0(GND_net), .I1(n17958[5]), .I2(n533_adj_4601), 
            .I3(n51805), .O(n17414[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_6 (.CI(n52012), .I0(n13590[3]), .I1(n369_adj_4615), 
            .CO(n52013));
    SB_LUT4 counter_2053_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n52718), .O(n51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_12 (.CI(n53010), .I0(n16478[9]), .I1(n816), .CO(n53011));
    SB_LUT4 add_6261_11_lut (.I0(GND_net), .I1(n16478[8]), .I2(n743), 
            .I3(n53009), .O(n15757[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_8 (.CI(n51805), .I0(n17958[5]), .I1(n533_adj_4601), 
            .CO(n51806));
    SB_CARRY counter_2053_add_4_18 (.CI(n52718), .I0(GND_net), .I1(counter[16]), 
            .CO(n52719));
    SB_LUT4 add_6347_7_lut (.I0(GND_net), .I1(n17958[4]), .I2(n460_adj_4598), 
            .I3(n51804), .O(n17414[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_5_lut (.I0(GND_net), .I1(n13590[2]), .I2(n296), .I3(n52011), 
            .O(n12570[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_20 (.CI(n51486), .I0(n257[18]), .I1(n306[18]), .CO(n51487));
    SB_CARRY add_6347_7 (.CI(n51804), .I0(n17958[4]), .I1(n460_adj_4598), 
            .CO(n51805));
    SB_CARRY add_6113_5 (.CI(n52011), .I0(n13590[2]), .I1(n296), .CO(n52012));
    SB_CARRY add_6261_11 (.CI(n53009), .I0(n16478[8]), .I1(n743), .CO(n53010));
    SB_LUT4 add_6261_10_lut (.I0(GND_net), .I1(n16478[7]), .I2(n670), 
            .I3(n53008), .O(n15757[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_10 (.CI(n53008), .I0(n16478[7]), .I1(n670), .CO(n53009));
    SB_LUT4 add_6261_9_lut (.I0(GND_net), .I1(n16478[6]), .I2(n597), .I3(n53007), 
            .O(n15757[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_6_lut (.I0(GND_net), .I1(n17958[3]), .I2(n387_adj_4596), 
            .I3(n51803), .O(n17414[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n52717), .O(n51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_9 (.CI(n53007), .I0(n16478[6]), .I1(n597), .CO(n53008));
    SB_LUT4 add_6261_8_lut (.I0(GND_net), .I1(n16478[5]), .I2(n524), .I3(n53006), 
            .O(n15757[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n306[17]), 
            .I3(n51485), .O(n356[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_6 (.CI(n51803), .I0(n17958[3]), .I1(n387_adj_4596), 
            .CO(n51804));
    SB_LUT4 add_6347_5_lut (.I0(GND_net), .I1(n17958[2]), .I2(n314), .I3(n51802), 
            .O(n17414[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n51485), .I0(n257[17]), .I1(n306[17]), .CO(n51486));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n306[16]), 
            .I3(n51484), .O(n356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_5 (.CI(n51802), .I0(n17958[2]), .I1(n314), .CO(n51803));
    SB_CARRY add_18_18 (.CI(n51484), .I0(n257[16]), .I1(n306[16]), .CO(n51485));
    SB_LUT4 add_6347_4_lut (.I0(GND_net), .I1(n17958[1]), .I2(n241), .I3(n51801), 
            .O(n17414[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_17 (.CI(n52717), .I0(GND_net), .I1(counter[15]), 
            .CO(n52718));
    SB_LUT4 add_6113_4_lut (.I0(GND_net), .I1(n13590[1]), .I2(n223), .I3(n52010), 
            .O(n12570[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_4 (.CI(n51801), .I0(n17958[1]), .I1(n241), .CO(n51802));
    SB_LUT4 add_6347_3_lut (.I0(GND_net), .I1(n17958[0]), .I2(n168), .I3(n51800), 
            .O(n17414[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_4 (.CI(n52010), .I0(n13590[1]), .I1(n223), .CO(n52011));
    SB_CARRY add_6347_3 (.CI(n51800), .I0(n17958[0]), .I1(n168), .CO(n51801));
    SB_LUT4 counter_2053_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n52716), .O(n51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6347_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17414[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6347_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_8 (.CI(n53006), .I0(n16478[5]), .I1(n524), .CO(n53007));
    SB_LUT4 add_6261_7_lut (.I0(GND_net), .I1(n16478[4]), .I2(n451), .I3(n53005), 
            .O(n15757[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n306[15]), 
            .I3(n51483), .O(n356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6347_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n51800));
    SB_LUT4 add_6547_9_lut (.I0(GND_net), .I1(n20405[6]), .I2(n630_adj_4589), 
            .I3(n51799), .O(n20278[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6113_3_lut (.I0(GND_net), .I1(n13590[0]), .I2(n150), .I3(n52009), 
            .O(n12570[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_3 (.CI(n52009), .I0(n13590[0]), .I1(n150), .CO(n52010));
    SB_LUT4 add_6547_8_lut (.I0(GND_net), .I1(n20405[5]), .I2(n557_adj_4587), 
            .I3(n51798), .O(n20278[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_7 (.CI(n53005), .I0(n16478[4]), .I1(n451), .CO(n53006));
    SB_LUT4 add_6113_2_lut (.I0(GND_net), .I1(n8_adj_4586), .I2(n77), 
            .I3(GND_net), .O(n12570[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6113_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6261_6_lut (.I0(GND_net), .I1(n16478[3]), .I2(n378_adj_4585), 
            .I3(n53004), .O(n15757[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_6 (.CI(n53004), .I0(n16478[3]), .I1(n378_adj_4585), 
            .CO(n53005));
    SB_CARRY add_18_17 (.CI(n51483), .I0(n257[15]), .I1(n306[15]), .CO(n51484));
    SB_CARRY counter_2053_add_4_16 (.CI(n52716), .I0(GND_net), .I1(counter[14]), 
            .CO(n52717));
    SB_LUT4 add_6261_5_lut (.I0(GND_net), .I1(n16478[2]), .I2(n305), .I3(n53003), 
            .O(n15757[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6547_8 (.CI(n51798), .I0(n20405[5]), .I1(n557_adj_4587), 
            .CO(n51799));
    SB_CARRY add_6261_5 (.CI(n53003), .I0(n16478[2]), .I1(n305), .CO(n53004));
    SB_LUT4 add_6261_4_lut (.I0(GND_net), .I1(n16478[1]), .I2(n232), .I3(n53002), 
            .O(n15757[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6113_2 (.CI(GND_net), .I0(n8_adj_4586), .I1(n77), .CO(n52009));
    SB_CARRY add_6261_4 (.CI(n53002), .I0(n16478[1]), .I1(n232), .CO(n53003));
    SB_LUT4 counter_2053_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n52715), .O(n51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6261_3_lut (.I0(GND_net), .I1(n16478[0]), .I2(n159), .I3(n53001), 
            .O(n15757[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6547_7_lut (.I0(GND_net), .I1(n20405[4]), .I2(n484_adj_4583), 
            .I3(n51797), .O(n20278[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_3 (.CI(n53001), .I0(n16478[0]), .I1(n159), .CO(n53002));
    SB_CARRY counter_2053_add_4_15 (.CI(n52715), .I0(GND_net), .I1(counter[13]), 
            .CO(n52716));
    SB_LUT4 add_6261_2_lut (.I0(GND_net), .I1(n17_adj_4582), .I2(n86), 
            .I3(GND_net), .O(n15757[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6261_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n52714), .O(n51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6261_2 (.CI(GND_net), .I0(n17_adj_4582), .I1(n86), .CO(n53001));
    SB_LUT4 add_6522_10_lut (.I0(GND_net), .I1(n20198[7]), .I2(n700), 
            .I3(n53000), .O(n20018[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_14 (.CI(n52714), .I0(GND_net), .I1(counter[12]), 
            .CO(n52715));
    SB_CARRY add_6547_7 (.CI(n51797), .I0(n20405[4]), .I1(n484_adj_4583), 
            .CO(n51798));
    SB_LUT4 add_6522_9_lut (.I0(GND_net), .I1(n20198[6]), .I2(n627), .I3(n52999), 
            .O(n20018[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6547_6_lut (.I0(GND_net), .I1(n20405[3]), .I2(n411_adj_4580), 
            .I3(n51796), .O(n20278[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_9 (.CI(n52999), .I0(n20198[6]), .I1(n627), .CO(n53000));
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[13] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2053_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n52713), .O(n51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6522_8_lut (.I0(GND_net), .I1(n20198[5]), .I2(n554), .I3(n52998), 
            .O(n20018[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6547_6 (.CI(n51796), .I0(n20405[3]), .I1(n411_adj_4580), 
            .CO(n51797));
    SB_CARRY add_6522_8 (.CI(n52998), .I0(n20198[5]), .I1(n554), .CO(n52999));
    SB_LUT4 add_6547_5_lut (.I0(GND_net), .I1(n20405[2]), .I2(n338_adj_4579), 
            .I3(n51795), .O(n20278[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6547_5 (.CI(n51795), .I0(n20405[2]), .I1(n338_adj_4579), 
            .CO(n51796));
    SB_CARRY counter_2053_add_4_13 (.CI(n52713), .I0(GND_net), .I1(counter[11]), 
            .CO(n52714));
    SB_LUT4 add_6522_7_lut (.I0(GND_net), .I1(n20198[4]), .I2(n481), .I3(n52997), 
            .O(n20018[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_7 (.CI(n52997), .I0(n20198[4]), .I1(n481), .CO(n52998));
    SB_LUT4 add_6522_6_lut (.I0(GND_net), .I1(n20198[3]), .I2(n408), .I3(n52996), 
            .O(n20018[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_6 (.CI(n52996), .I0(n20198[3]), .I1(n408), .CO(n52997));
    SB_LUT4 add_6522_5_lut (.I0(GND_net), .I1(n20198[2]), .I2(n335), .I3(n52995), 
            .O(n20018[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_5 (.CI(n52995), .I0(n20198[2]), .I1(n335), .CO(n52996));
    SB_LUT4 add_6547_4_lut (.I0(GND_net), .I1(n20405[1]), .I2(n265_adj_4577), 
            .I3(n51794), .O(n20278[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6522_4_lut (.I0(GND_net), .I1(n20198[1]), .I2(n262), .I3(n52994), 
            .O(n20018[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_4 (.CI(n52994), .I0(n20198[1]), .I1(n262), .CO(n52995));
    SB_LUT4 add_6522_3_lut (.I0(GND_net), .I1(n20198[0]), .I2(n189_adj_4576), 
            .I3(n52993), .O(n20018[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n52712), .O(n51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6547_4 (.CI(n51794), .I0(n20405[1]), .I1(n265_adj_4577), 
            .CO(n51795));
    SB_CARRY add_6522_3 (.CI(n52993), .I0(n20198[0]), .I1(n189_adj_4576), 
            .CO(n52994));
    SB_LUT4 add_6522_2_lut (.I0(GND_net), .I1(n47_adj_4575), .I2(n116_adj_4574), 
            .I3(GND_net), .O(n20018[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6522_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6522_2 (.CI(GND_net), .I0(n47_adj_4575), .I1(n116_adj_4574), 
            .CO(n52993));
    SB_LUT4 add_6297_19_lut (.I0(GND_net), .I1(n17125[16]), .I2(GND_net), 
            .I3(n52992), .O(n16478[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6297_18_lut (.I0(GND_net), .I1(n17125[15]), .I2(GND_net), 
            .I3(n52991), .O(n16478[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n306[14]), 
            .I3(n51482), .O(n356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6547_3_lut (.I0(GND_net), .I1(n20405[0]), .I2(n192_adj_4573), 
            .I3(n51793), .O(n20278[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_18 (.CI(n52991), .I0(n17125[15]), .I1(GND_net), 
            .CO(n52992));
    SB_LUT4 add_6297_17_lut (.I0(GND_net), .I1(n17125[14]), .I2(GND_net), 
            .I3(n52990), .O(n16478[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_17 (.CI(n52990), .I0(n17125[14]), .I1(GND_net), 
            .CO(n52991));
    SB_LUT4 add_6297_16_lut (.I0(GND_net), .I1(n17125[13]), .I2(n1111), 
            .I3(n52989), .O(n16478[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_12 (.CI(n52712), .I0(GND_net), .I1(counter[10]), 
            .CO(n52713));
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n219));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6297_16 (.CI(n52989), .I0(n17125[13]), .I1(n1111), .CO(n52990));
    SB_LUT4 add_6297_15_lut (.I0(GND_net), .I1(n17125[12]), .I2(n1038), 
            .I3(n52988), .O(n16478[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6547_3 (.CI(n51793), .I0(n20405[0]), .I1(n192_adj_4573), 
            .CO(n51794));
    SB_CARRY add_6297_15 (.CI(n52988), .I0(n17125[12]), .I1(n1038), .CO(n52989));
    SB_LUT4 counter_2053_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n52711), .O(n51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_16 (.CI(n51482), .I0(n257[14]), .I1(n306[14]), .CO(n51483));
    SB_LUT4 add_6547_2_lut (.I0(GND_net), .I1(n50_adj_4568), .I2(n119_adj_4567), 
            .I3(GND_net), .O(n20278[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6547_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6297_14_lut (.I0(GND_net), .I1(n17125[11]), .I2(n965), 
            .I3(n52987), .O(n16478[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_14 (.CI(n52987), .I0(n17125[11]), .I1(n965), .CO(n52988));
    SB_CARRY add_6547_2 (.CI(GND_net), .I0(n50_adj_4568), .I1(n119_adj_4567), 
            .CO(n51793));
    SB_LUT4 add_6297_13_lut (.I0(GND_net), .I1(n17125[10]), .I2(n892), 
            .I3(n52986), .O(n16478[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_13 (.CI(n52986), .I0(n17125[10]), .I1(n892), .CO(n52987));
    SB_LUT4 add_6297_12_lut (.I0(GND_net), .I1(n17125[9]), .I2(n819), 
            .I3(n52985), .O(n16478[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_11 (.CI(n52711), .I0(GND_net), .I1(counter[9]), 
            .CO(n52712));
    SB_LUT4 counter_2053_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n52710), .O(n51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_12 (.CI(n52985), .I0(n17125[9]), .I1(n819), .CO(n52986));
    SB_LUT4 add_6297_11_lut (.I0(GND_net), .I1(n17125[8]), .I2(n746), 
            .I3(n52984), .O(n16478[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_10 (.CI(n52710), .I0(GND_net), .I1(counter[8]), 
            .CO(n52711));
    SB_CARRY add_6297_11 (.CI(n52984), .I0(n17125[8]), .I1(n746), .CO(n52985));
    SB_LUT4 add_6297_10_lut (.I0(GND_net), .I1(n17125[7]), .I2(n673), 
            .I3(n52983), .O(n16478[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n52709), .O(n51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_10 (.CI(n52983), .I0(n17125[7]), .I1(n673), .CO(n52984));
    SB_CARRY counter_2053_add_4_9 (.CI(n52709), .I0(GND_net), .I1(counter[7]), 
            .CO(n52710));
    SB_LUT4 add_6297_9_lut (.I0(GND_net), .I1(n17125[6]), .I2(n600), .I3(n52982), 
            .O(n16478[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 counter_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n52708), .O(n51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_9 (.CI(n52982), .I0(n17125[6]), .I1(n600), .CO(n52983));
    SB_LUT4 add_6297_8_lut (.I0(GND_net), .I1(n17125[5]), .I2(n527), .I3(n52981), 
            .O(n16478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_8 (.CI(n52981), .I0(n17125[5]), .I1(n527), .CO(n52982));
    SB_CARRY counter_2053_add_4_8 (.CI(n52708), .I0(GND_net), .I1(counter[6]), 
            .CO(n52709));
    SB_LUT4 add_6297_7_lut (.I0(GND_net), .I1(n17125[4]), .I2(n454), .I3(n52980), 
            .O(n16478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_7 (.CI(n52980), .I0(n17125[4]), .I1(n454), .CO(n52981));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n306[13]), 
            .I3(n51481), .O(n356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6297_6_lut (.I0(GND_net), .I1(n17125[3]), .I2(n381), .I3(n52979), 
            .O(n16478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_6 (.CI(n52979), .I0(n17125[3]), .I1(n381), .CO(n52980));
    SB_LUT4 counter_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n52707), .O(n51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_7 (.CI(n52707), .I0(GND_net), .I1(counter[5]), 
            .CO(n52708));
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6297_5_lut (.I0(GND_net), .I1(n17125[2]), .I2(n308), .I3(n52978), 
            .O(n16478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_15 (.CI(n51481), .I0(n257[13]), .I1(n306[13]), .CO(n51482));
    SB_CARRY add_6297_5 (.CI(n52978), .I0(n17125[2]), .I1(n308), .CO(n52979));
    SB_LUT4 counter_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n52706), .O(n51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6297_4_lut (.I0(GND_net), .I1(n17125[1]), .I2(n235), .I3(n52977), 
            .O(n16478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_6 (.CI(n52706), .I0(GND_net), .I1(counter[4]), 
            .CO(n52707));
    SB_CARRY add_6297_4 (.CI(n52977), .I0(n17125[1]), .I1(n235), .CO(n52978));
    SB_LUT4 counter_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n52705), .O(n51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_5 (.CI(n52705), .I0(GND_net), .I1(counter[3]), 
            .CO(n52706));
    SB_LUT4 counter_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n52704), .O(n51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY counter_2053_add_4_4 (.CI(n52704), .I0(GND_net), .I1(counter[2]), 
            .CO(n52705));
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6297_3_lut (.I0(GND_net), .I1(n17125[0]), .I2(n162), .I3(n52976), 
            .O(n16478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n52703), .O(n51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_3 (.CI(n52703), .I0(GND_net), .I1(counter[1]), 
            .CO(n52704));
    SB_CARRY add_6297_3 (.CI(n52976), .I0(n17125[0]), .I1(n162), .CO(n52977));
    SB_LUT4 add_6297_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n16478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6297_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6297_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n52976));
    SB_LUT4 counter_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6331_18_lut (.I0(GND_net), .I1(n17702[15]), .I2(GND_net), 
            .I3(n52975), .O(n17125[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n52703));
    SB_LUT4 add_6331_17_lut (.I0(GND_net), .I1(n17702[14]), .I2(GND_net), 
            .I3(n52974), .O(n17125[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_17 (.CI(n52974), .I0(n17702[14]), .I1(GND_net), 
            .CO(n52975));
    SB_LUT4 add_6331_16_lut (.I0(GND_net), .I1(n17702[13]), .I2(n1114), 
            .I3(n52973), .O(n17125[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_16 (.CI(n52973), .I0(n17702[13]), .I1(n1114), .CO(n52974));
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[11] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6331_15_lut (.I0(GND_net), .I1(n17702[12]), .I2(n1041), 
            .I3(n52972), .O(n17125[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_15 (.CI(n52972), .I0(n17702[12]), .I1(n1041), .CO(n52973));
    SB_LUT4 add_6331_14_lut (.I0(GND_net), .I1(n17702[11]), .I2(n968), 
            .I3(n52971), .O(n17125[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_14 (.CI(n52971), .I0(n17702[11]), .I1(n968), .CO(n52972));
    SB_LUT4 add_6331_13_lut (.I0(GND_net), .I1(n17702[10]), .I2(n895), 
            .I3(n52970), .O(n17125[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_13 (.CI(n52970), .I0(n17702[10]), .I1(n895), .CO(n52971));
    SB_LUT4 add_6331_12_lut (.I0(GND_net), .I1(n17702[9]), .I2(n822), 
            .I3(n52969), .O(n17125[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_12 (.CI(n52969), .I0(n17702[9]), .I1(n822), .CO(n52970));
    SB_LUT4 add_6331_11_lut (.I0(GND_net), .I1(n17702[8]), .I2(n749), 
            .I3(n52968), .O(n17125[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_11 (.CI(n52968), .I0(n17702[8]), .I1(n749), .CO(n52969));
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6331_10_lut (.I0(GND_net), .I1(n17702[7]), .I2(n676), 
            .I3(n52967), .O(n17125[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_10 (.CI(n52967), .I0(n17702[7]), .I1(n676), .CO(n52968));
    SB_LUT4 add_6331_9_lut (.I0(GND_net), .I1(n17702[6]), .I2(n603), .I3(n52966), 
            .O(n17125[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_9 (.CI(n52966), .I0(n17702[6]), .I1(n603), .CO(n52967));
    SB_LUT4 add_6331_8_lut (.I0(GND_net), .I1(n17702[5]), .I2(n530), .I3(n52965), 
            .O(n17125[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_8 (.CI(n52965), .I0(n17702[5]), .I1(n530), .CO(n52966));
    SB_LUT4 add_6331_7_lut (.I0(GND_net), .I1(n17702[4]), .I2(n457), .I3(n52964), 
            .O(n17125[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_7 (.CI(n52964), .I0(n17702[4]), .I1(n457), .CO(n52965));
    SB_LUT4 add_6331_6_lut (.I0(GND_net), .I1(n17702[3]), .I2(n384_adj_4564), 
            .I3(n52963), .O(n17125[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_6 (.CI(n52963), .I0(n17702[3]), .I1(n384_adj_4564), 
            .CO(n52964));
    SB_LUT4 add_6331_5_lut (.I0(GND_net), .I1(n17702[2]), .I2(n311), .I3(n52962), 
            .O(n17125[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_5 (.CI(n52962), .I0(n17702[2]), .I1(n311), .CO(n52963));
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6331_4_lut (.I0(GND_net), .I1(n17702[1]), .I2(n238), .I3(n52961), 
            .O(n17125[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_4 (.CI(n52961), .I0(n17702[1]), .I1(n238), .CO(n52962));
    SB_LUT4 add_6331_3_lut (.I0(GND_net), .I1(n17702[0]), .I2(n165), .I3(n52960), 
            .O(n17125[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_3 (.CI(n52960), .I0(n17702[0]), .I1(n165), .CO(n52961));
    SB_LUT4 add_6331_2_lut (.I0(GND_net), .I1(n23_adj_4561), .I2(n92), 
            .I3(GND_net), .O(n17125[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6331_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6331_2 (.CI(GND_net), .I0(n23_adj_4561), .I1(n92), .CO(n52960));
    SB_LUT4 add_6539_9_lut (.I0(GND_net), .I1(n20342[6]), .I2(n630), .I3(n52959), 
            .O(n20198[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6539_8_lut (.I0(GND_net), .I1(n20342[5]), .I2(n557), .I3(n52958), 
            .O(n20198[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_8 (.CI(n52958), .I0(n20342[5]), .I1(n557), .CO(n52959));
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6539_7_lut (.I0(GND_net), .I1(n20342[4]), .I2(n484), .I3(n52957), 
            .O(n20198[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_7 (.CI(n52957), .I0(n20342[4]), .I1(n484), .CO(n52958));
    SB_LUT4 add_6539_6_lut (.I0(GND_net), .I1(n20342[3]), .I2(n411), .I3(n52956), 
            .O(n20198[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_6 (.CI(n52956), .I0(n20342[3]), .I1(n411), .CO(n52957));
    SB_LUT4 add_6539_5_lut (.I0(GND_net), .I1(n20342[2]), .I2(n338), .I3(n52955), 
            .O(n20198[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_5 (.CI(n52955), .I0(n20342[2]), .I1(n338), .CO(n52956));
    SB_LUT4 add_6539_4_lut (.I0(GND_net), .I1(n20342[1]), .I2(n265), .I3(n52954), 
            .O(n20198[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_4 (.CI(n52954), .I0(n20342[1]), .I1(n265), .CO(n52955));
    SB_LUT4 add_6539_3_lut (.I0(GND_net), .I1(n20342[0]), .I2(n192), .I3(n52953), 
            .O(n20198[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6378_16_lut (.I0(GND_net), .I1(n18438[13]), .I2(n1120), 
            .I3(n51781), .O(n17958[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6378_15_lut (.I0(GND_net), .I1(n18438[12]), .I2(n1047), 
            .I3(n51780), .O(n17958[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_3 (.CI(n52953), .I0(n20342[0]), .I1(n192), .CO(n52954));
    SB_LUT4 add_6539_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20198[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6539_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6539_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n52953));
    SB_LUT4 add_6363_17_lut (.I0(GND_net), .I1(n18213[14]), .I2(GND_net), 
            .I3(n52952), .O(n17702[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n306[12]), 
            .I3(n51480), .O(n356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_15 (.CI(n51780), .I0(n18438[12]), .I1(n1047), .CO(n51781));
    SB_CARRY add_18_14 (.CI(n51480), .I0(n257[12]), .I1(n306[12]), .CO(n51481));
    SB_LUT4 add_6363_16_lut (.I0(GND_net), .I1(n18213[13]), .I2(n1117), 
            .I3(n52951), .O(n17702[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_16 (.CI(n52951), .I0(n18213[13]), .I1(n1117), .CO(n52952));
    SB_LUT4 add_6378_14_lut (.I0(GND_net), .I1(n18438[11]), .I2(n974), 
            .I3(n51779), .O(n17958[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_14 (.CI(n51779), .I0(n18438[11]), .I1(n974), .CO(n51780));
    SB_LUT4 add_6378_13_lut (.I0(GND_net), .I1(n18438[10]), .I2(n901), 
            .I3(n51778), .O(n17958[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6363_15_lut (.I0(GND_net), .I1(n18213[12]), .I2(n1044), 
            .I3(n52950), .O(n17702[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_15 (.CI(n52950), .I0(n18213[12]), .I1(n1044), .CO(n52951));
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n306[11]), 
            .I3(n51479), .O(n356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6363_14_lut (.I0(GND_net), .I1(n18213[11]), .I2(n971), 
            .I3(n52949), .O(n17702[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_14 (.CI(n52949), .I0(n18213[11]), .I1(n971), .CO(n52950));
    SB_LUT4 add_6363_13_lut (.I0(GND_net), .I1(n18213[10]), .I2(n898), 
            .I3(n52948), .O(n17702[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_13 (.CI(n52948), .I0(n18213[10]), .I1(n898), .CO(n52949));
    SB_LUT4 add_6363_12_lut (.I0(GND_net), .I1(n18213[9]), .I2(n825), 
            .I3(n52947), .O(n17702[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_13 (.CI(n51778), .I0(n18438[10]), .I1(n901), .CO(n51779));
    SB_CARRY add_6363_12 (.CI(n52947), .I0(n18213[9]), .I1(n825), .CO(n52948));
    SB_LUT4 add_6363_11_lut (.I0(GND_net), .I1(n18213[8]), .I2(n752), 
            .I3(n52946), .O(n17702[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_11 (.CI(n52946), .I0(n18213[8]), .I1(n752), .CO(n52947));
    SB_LUT4 add_6378_12_lut (.I0(GND_net), .I1(n18438[9]), .I2(n828), 
            .I3(n51777), .O(n17958[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_12 (.CI(n51777), .I0(n18438[9]), .I1(n828), .CO(n51778));
    SB_LUT4 add_6363_10_lut (.I0(GND_net), .I1(n18213[7]), .I2(n679), 
            .I3(n52945), .O(n17702[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_10 (.CI(n52945), .I0(n18213[7]), .I1(n679), .CO(n52946));
    SB_CARRY add_18_13 (.CI(n51479), .I0(n257[11]), .I1(n306[11]), .CO(n51480));
    SB_LUT4 add_6363_9_lut (.I0(GND_net), .I1(n18213[6]), .I2(n606), .I3(n52944), 
            .O(n17702[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_9 (.CI(n52944), .I0(n18213[6]), .I1(n606), .CO(n52945));
    SB_LUT4 add_6363_8_lut (.I0(GND_net), .I1(n18213[5]), .I2(n533), .I3(n52943), 
            .O(n17702[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_8 (.CI(n52943), .I0(n18213[5]), .I1(n533), .CO(n52944));
    SB_LUT4 add_6363_7_lut (.I0(GND_net), .I1(n18213[4]), .I2(n460), .I3(n52942), 
            .O(n17702[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_7 (.CI(n52942), .I0(n18213[4]), .I1(n460), .CO(n52943));
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[10] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6363_6_lut (.I0(GND_net), .I1(n18213[3]), .I2(n387_adj_4980), 
            .I3(n52941), .O(n17702[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_6 (.CI(n52941), .I0(n18213[3]), .I1(n387_adj_4980), 
            .CO(n52942));
    SB_LUT4 add_6378_11_lut (.I0(GND_net), .I1(n18438[8]), .I2(n755_adj_4979), 
            .I3(n51776), .O(n17958[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_11 (.CI(n51776), .I0(n18438[8]), .I1(n755_adj_4979), 
            .CO(n51777));
    SB_LUT4 add_6363_5_lut (.I0(GND_net), .I1(n18213[2]), .I2(n314_adj_4978), 
            .I3(n52940), .O(n17702[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_5 (.CI(n52940), .I0(n18213[2]), .I1(n314_adj_4978), 
            .CO(n52941));
    SB_LUT4 add_6378_10_lut (.I0(GND_net), .I1(n18438[7]), .I2(n682_adj_4977), 
            .I3(n51775), .O(n17958[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6363_4_lut (.I0(GND_net), .I1(n18213[1]), .I2(n241_adj_4976), 
            .I3(n52939), .O(n17702[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_4 (.CI(n52939), .I0(n18213[1]), .I1(n241_adj_4976), 
            .CO(n52940));
    SB_LUT4 add_6363_3_lut (.I0(GND_net), .I1(n18213[0]), .I2(n168_adj_4974), 
            .I3(n52938), .O(n17702[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_3 (.CI(n52938), .I0(n18213[0]), .I1(n168_adj_4974), 
            .CO(n52939));
    SB_LUT4 add_6363_2_lut (.I0(GND_net), .I1(n26_adj_4973), .I2(n95_adj_4972), 
            .I3(GND_net), .O(n17702[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6363_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6363_2 (.CI(GND_net), .I0(n26_adj_4973), .I1(n95_adj_4972), 
            .CO(n52938));
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n306[10]), 
            .I3(n51478), .O(n356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6393_16_lut (.I0(GND_net), .I1(n18662[13]), .I2(n1120_adj_4971), 
            .I3(n52937), .O(n18213[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_10 (.CI(n51775), .I0(n18438[7]), .I1(n682_adj_4977), 
            .CO(n51776));
    SB_LUT4 add_6378_9_lut (.I0(GND_net), .I1(n18438[6]), .I2(n609_adj_4970), 
            .I3(n51774), .O(n17958[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6393_15_lut (.I0(GND_net), .I1(n18662[12]), .I2(n1047_adj_4969), 
            .I3(n52936), .O(n18213[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_15 (.CI(n52936), .I0(n18662[12]), .I1(n1047_adj_4969), 
            .CO(n52937));
    SB_CARRY add_18_12 (.CI(n51478), .I0(n257[10]), .I1(n306[10]), .CO(n51479));
    SB_CARRY add_6378_9 (.CI(n51774), .I0(n18438[6]), .I1(n609_adj_4970), 
            .CO(n51775));
    SB_LUT4 add_6393_14_lut (.I0(GND_net), .I1(n18662[11]), .I2(n974_adj_4968), 
            .I3(n52935), .O(n18213[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_14 (.CI(n52935), .I0(n18662[11]), .I1(n974_adj_4968), 
            .CO(n52936));
    SB_LUT4 add_6393_13_lut (.I0(GND_net), .I1(n18662[10]), .I2(n901_adj_4967), 
            .I3(n52934), .O(n18213[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_13 (.CI(n52934), .I0(n18662[10]), .I1(n901_adj_4967), 
            .CO(n52935));
    SB_LUT4 add_6393_12_lut (.I0(GND_net), .I1(n18662[9]), .I2(n828_adj_4966), 
            .I3(n52933), .O(n18213[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6378_8_lut (.I0(GND_net), .I1(n18438[5]), .I2(n536_adj_4965), 
            .I3(n51773), .O(n17958[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_12 (.CI(n52933), .I0(n18662[9]), .I1(n828_adj_4966), 
            .CO(n52934));
    SB_LUT4 add_6393_11_lut (.I0(GND_net), .I1(n18662[8]), .I2(n755), 
            .I3(n52932), .O(n18213[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_11 (.CI(n52932), .I0(n18662[8]), .I1(n755), .CO(n52933));
    SB_LUT4 add_6393_10_lut (.I0(GND_net), .I1(n18662[7]), .I2(n682), 
            .I3(n52931), .O(n18213[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[9] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6378_8 (.CI(n51773), .I0(n18438[5]), .I1(n536_adj_4965), 
            .CO(n51774));
    SB_CARRY add_6393_10 (.CI(n52931), .I0(n18662[7]), .I1(n682), .CO(n52932));
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n306[9]), .I3(n51477), 
            .O(n356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6378_7_lut (.I0(GND_net), .I1(n18438[4]), .I2(n463_adj_4964), 
            .I3(n51772), .O(n17958[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6393_9_lut (.I0(GND_net), .I1(n18662[6]), .I2(n609), .I3(n52930), 
            .O(n18213[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6378_7 (.CI(n51772), .I0(n18438[4]), .I1(n463_adj_4964), 
            .CO(n51773));
    SB_LUT4 add_6378_6_lut (.I0(GND_net), .I1(n18438[3]), .I2(n390_adj_4961), 
            .I3(n51771), .O(n17958[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_6 (.CI(n51771), .I0(n18438[3]), .I1(n390_adj_4961), 
            .CO(n51772));
    SB_CARRY add_6393_9 (.CI(n52930), .I0(n18662[6]), .I1(n609), .CO(n52931));
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_18_11 (.CI(n51477), .I0(n257[9]), .I1(n306[9]), .CO(n51478));
    SB_LUT4 add_6160_22_lut (.I0(GND_net), .I1(n14518[19]), .I2(GND_net), 
            .I3(n51991), .O(n13590[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6378_5_lut (.I0(GND_net), .I1(n18438[2]), .I2(n317_adj_4960), 
            .I3(n51770), .O(n17958[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6393_8_lut (.I0(GND_net), .I1(n18662[5]), .I2(n536), .I3(n52929), 
            .O(n18213[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_5 (.CI(n51770), .I0(n18438[2]), .I1(n317_adj_4960), 
            .CO(n51771));
    SB_LUT4 add_6378_4_lut (.I0(GND_net), .I1(n18438[1]), .I2(n244_adj_4959), 
            .I3(n51769), .O(n17958[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_8 (.CI(n52929), .I0(n18662[5]), .I1(n536), .CO(n52930));
    SB_LUT4 add_6160_21_lut (.I0(GND_net), .I1(n14518[18]), .I2(GND_net), 
            .I3(n51990), .O(n13590[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[8] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6393_7_lut (.I0(GND_net), .I1(n18662[4]), .I2(n463), .I3(n52928), 
            .O(n18213[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_7 (.CI(n52928), .I0(n18662[4]), .I1(n463), .CO(n52929));
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n306[8]), .I3(n51476), 
            .O(n356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_21 (.CI(n51990), .I0(n14518[18]), .I1(GND_net), 
            .CO(n51991));
    SB_LUT4 add_6393_6_lut (.I0(GND_net), .I1(n18662[3]), .I2(n390_adj_4957), 
            .I3(n52927), .O(n18213[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_6 (.CI(n52927), .I0(n18662[3]), .I1(n390_adj_4957), 
            .CO(n52928));
    SB_LUT4 add_6393_5_lut (.I0(GND_net), .I1(n18662[2]), .I2(n317), .I3(n52926), 
            .O(n18213[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_5 (.CI(n52926), .I0(n18662[2]), .I1(n317), .CO(n52927));
    SB_CARRY add_6378_4 (.CI(n51769), .I0(n18438[1]), .I1(n244_adj_4959), 
            .CO(n51770));
    SB_LUT4 add_6378_3_lut (.I0(GND_net), .I1(n18438[0]), .I2(n171_adj_4956), 
            .I3(n51768), .O(n17958[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6393_4_lut (.I0(GND_net), .I1(n18662[1]), .I2(n244), .I3(n52925), 
            .O(n18213[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[7] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6160_20_lut (.I0(GND_net), .I1(n14518[17]), .I2(GND_net), 
            .I3(n51989), .O(n13590[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6393_4 (.CI(n52925), .I0(n18662[1]), .I1(n244), .CO(n52926));
    SB_LUT4 add_6393_3_lut (.I0(GND_net), .I1(n18662[0]), .I2(n171), .I3(n52924), 
            .O(n18213[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_3 (.CI(n52924), .I0(n18662[0]), .I1(n171), .CO(n52925));
    SB_LUT4 add_6393_2_lut (.I0(GND_net), .I1(n29_adj_4954), .I2(n98_adj_4953), 
            .I3(GND_net), .O(n18213[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6393_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6393_2 (.CI(GND_net), .I0(n29_adj_4954), .I1(n98_adj_4953), 
            .CO(n52924));
    SB_LUT4 add_6554_8_lut (.I0(GND_net), .I1(n20454[5]), .I2(n560_adj_4952), 
            .I3(n52923), .O(n20342[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6554_7_lut (.I0(GND_net), .I1(n20454[4]), .I2(n487_adj_4951), 
            .I3(n52922), .O(n20342[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6554_7 (.CI(n52922), .I0(n20454[4]), .I1(n487_adj_4951), 
            .CO(n52923));
    SB_LUT4 add_6554_6_lut (.I0(GND_net), .I1(n20454[3]), .I2(n414_adj_4950), 
            .I3(n52921), .O(n20342[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6554_6 (.CI(n52921), .I0(n20454[3]), .I1(n414_adj_4950), 
            .CO(n52922));
    SB_LUT4 add_6554_5_lut (.I0(GND_net), .I1(n20454[2]), .I2(n341_adj_4949), 
            .I3(n52920), .O(n20342[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6554_5 (.CI(n52920), .I0(n20454[2]), .I1(n341_adj_4949), 
            .CO(n52921));
    SB_LUT4 add_6554_4_lut (.I0(GND_net), .I1(n20454[1]), .I2(n268_adj_4948), 
            .I3(n52919), .O(n20342[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[6] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_c));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(51[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n356[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5059));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n356[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5060));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i45_2_lut (.I0(PWMLimit[22]), .I1(n356[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5061));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6554_4 (.CI(n52919), .I0(n20454[1]), .I1(n268_adj_4948), 
            .CO(n52920));
    SB_LUT4 add_6554_3_lut (.I0(GND_net), .I1(n20454[0]), .I2(n195_adj_4947), 
            .I3(n52918), .O(n20342[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5062));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6554_3 (.CI(n52918), .I0(n20454[0]), .I1(n195_adj_4947), 
            .CO(n52919));
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n356[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5063));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6554_2_lut (.I0(GND_net), .I1(n53_adj_4946), .I2(n122_adj_4945), 
            .I3(GND_net), .O(n20342[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6554_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i6_3_lut (.I0(n149), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_18_10 (.CI(n51476), .I0(n257[8]), .I1(n306[8]), .CO(n51477));
    SB_CARRY add_6554_2 (.CI(GND_net), .I0(n53_adj_4946), .I1(n122_adj_4945), 
            .CO(n52918));
    SB_LUT4 add_6421_15_lut (.I0(GND_net), .I1(n19053[12]), .I2(n1050_adj_4944), 
            .I3(n52917), .O(n18662[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_14_lut (.I0(GND_net), .I1(n19053[11]), .I2(n977_adj_4943), 
            .I3(n52916), .O(n18662[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n356[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5065));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6421_14 (.CI(n52916), .I0(n19053[11]), .I1(n977_adj_4943), 
            .CO(n52917));
    SB_LUT4 add_6421_13_lut (.I0(GND_net), .I1(n19053[10]), .I2(n904_adj_4942), 
            .I3(n52915), .O(n18662[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_13 (.CI(n52915), .I0(n19053[10]), .I1(n904_adj_4942), 
            .CO(n52916));
    SB_LUT4 add_6421_12_lut (.I0(GND_net), .I1(n19053[9]), .I2(n831_adj_4941), 
            .I3(n52914), .O(n18662[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_12 (.CI(n52914), .I0(n19053[9]), .I1(n831_adj_4941), 
            .CO(n52915));
    SB_LUT4 add_6421_11_lut (.I0(GND_net), .I1(n19053[8]), .I2(n758_adj_4939), 
            .I3(n52913), .O(n18662[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_20 (.CI(n51989), .I0(n14518[17]), .I1(GND_net), 
            .CO(n51990));
    SB_CARRY add_6421_11 (.CI(n52913), .I0(n19053[8]), .I1(n758_adj_4939), 
            .CO(n52914));
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[5] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6421_10_lut (.I0(GND_net), .I1(n19053[7]), .I2(n685_adj_4938), 
            .I3(n52912), .O(n18662[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6378_3 (.CI(n51768), .I0(n18438[0]), .I1(n171_adj_4956), 
            .CO(n51769));
    SB_CARRY add_6421_10 (.CI(n52912), .I0(n19053[7]), .I1(n685_adj_4938), 
            .CO(n52913));
    SB_LUT4 add_6421_9_lut (.I0(GND_net), .I1(n19053[6]), .I2(n612_adj_4937), 
            .I3(n52911), .O(n18662[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_9 (.CI(n52911), .I0(n19053[6]), .I1(n612_adj_4937), 
            .CO(n52912));
    SB_LUT4 add_6378_2_lut (.I0(GND_net), .I1(n29_adj_4936), .I2(n98), 
            .I3(GND_net), .O(n17958[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6378_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_8_lut (.I0(GND_net), .I1(n19053[5]), .I2(n539_adj_4935), 
            .I3(n52910), .O(n18662[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_8 (.CI(n52910), .I0(n19053[5]), .I1(n539_adj_4935), 
            .CO(n52911));
    SB_LUT4 add_6421_7_lut (.I0(GND_net), .I1(n19053[4]), .I2(n466_adj_4934), 
            .I3(n52909), .O(n18662[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_7 (.CI(n52909), .I0(n19053[4]), .I1(n466_adj_4934), 
            .CO(n52910));
    SB_LUT4 LessThan_23_i29_2_lut (.I0(PWMLimit[14]), .I1(n356[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5066));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i31_2_lut (.I0(PWMLimit[15]), .I1(n356[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5067));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n356[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5068));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i35_2_lut (.I0(PWMLimit[17]), .I1(n356[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5069));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6421_6_lut (.I0(GND_net), .I1(n19053[3]), .I2(n393_adj_4933), 
            .I3(n52908), .O(n18662[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_6 (.CI(n52908), .I0(n19053[3]), .I1(n393_adj_4933), 
            .CO(n52909));
    SB_LUT4 add_6421_5_lut (.I0(GND_net), .I1(n19053[2]), .I2(n320_adj_4932), 
            .I3(n52907), .O(n18662[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6421_5 (.CI(n52907), .I0(n19053[2]), .I1(n320_adj_4932), 
            .CO(n52908));
    SB_LUT4 add_6421_4_lut (.I0(GND_net), .I1(n19053[1]), .I2(n247_adj_4931), 
            .I3(n52906), .O(n18662[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i33_2_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5070));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n356[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5071));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6160_19_lut (.I0(GND_net), .I1(n14518[16]), .I2(GND_net), 
            .I3(n51988), .O(n13590[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_19 (.CI(n51988), .I0(n14518[16]), .I1(GND_net), 
            .CO(n51989));
    SB_CARRY add_6378_2 (.CI(GND_net), .I0(n29_adj_4936), .I1(n98), .CO(n51768));
    SB_CARRY add_6421_4 (.CI(n52906), .I0(n19053[1]), .I1(n247_adj_4931), 
            .CO(n52907));
    SB_LUT4 add_6421_3_lut (.I0(GND_net), .I1(n19053[0]), .I2(n174_adj_4930), 
            .I3(n52905), .O(n18662[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_3 (.CI(n52905), .I0(n19053[0]), .I1(n174_adj_4930), 
            .CO(n52906));
    SB_LUT4 add_6421_2_lut (.I0(GND_net), .I1(n32_adj_4929), .I2(n101_adj_4928), 
            .I3(GND_net), .O(n18662[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_2 (.CI(GND_net), .I0(n32_adj_4929), .I1(n101_adj_4928), 
            .CO(n52905));
    SB_LUT4 add_6447_14_lut (.I0(GND_net), .I1(n19390[11]), .I2(n980_adj_4927), 
            .I3(n52904), .O(n19053[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n356[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5072));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n356[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5073));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6160_18_lut (.I0(GND_net), .I1(n14518[15]), .I2(GND_net), 
            .I3(n51987), .O(n13590[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6447_13_lut (.I0(GND_net), .I1(n19390[10]), .I2(n907_adj_4926), 
            .I3(n52903), .O(n19053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_13 (.CI(n52903), .I0(n19390[10]), .I1(n907_adj_4926), 
            .CO(n52904));
    SB_LUT4 add_6447_12_lut (.I0(GND_net), .I1(n19390[9]), .I2(n834_adj_4925), 
            .I3(n52902), .O(n19053[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_12 (.CI(n52902), .I0(n19390[9]), .I1(n834_adj_4925), 
            .CO(n52903));
    SB_LUT4 add_6447_11_lut (.I0(GND_net), .I1(n19390[8]), .I2(n761_adj_4924), 
            .I3(n52901), .O(n19053[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_11 (.CI(n52901), .I0(n19390[8]), .I1(n761_adj_4924), 
            .CO(n52902));
    SB_LUT4 add_6447_10_lut (.I0(GND_net), .I1(n19390[7]), .I2(n688_adj_4923), 
            .I3(n52900), .O(n19053[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[4] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i27_2_lut (.I0(PWMLimit[13]), .I1(n356[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5074));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n356[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5075));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6447_10 (.CI(n52900), .I0(n19390[7]), .I1(n688_adj_4923), 
            .CO(n52901));
    SB_LUT4 add_6447_9_lut (.I0(GND_net), .I1(n19390[6]), .I2(n615_adj_4922), 
            .I3(n52899), .O(n19053[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_9 (.CI(n52899), .I0(n19390[6]), .I1(n615_adj_4922), 
            .CO(n52900));
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n306[7]), .I3(n51475), 
            .O(n356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[3] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6160_18 (.CI(n51987), .I0(n14518[15]), .I1(GND_net), 
            .CO(n51988));
    SB_LUT4 add_6160_17_lut (.I0(GND_net), .I1(n14518[14]), .I2(GND_net), 
            .I3(n51986), .O(n13590[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_17 (.CI(n51986), .I0(n14518[14]), .I1(GND_net), 
            .CO(n51987));
    SB_LUT4 add_6447_8_lut (.I0(GND_net), .I1(n19390[5]), .I2(n542_adj_4920), 
            .I3(n52898), .O(n19053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_8 (.CI(n52898), .I0(n19390[5]), .I1(n542_adj_4920), 
            .CO(n52899));
    SB_LUT4 add_6160_16_lut (.I0(GND_net), .I1(n14518[13]), .I2(n1102), 
            .I3(n51985), .O(n13590[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_16 (.CI(n51985), .I0(n14518[13]), .I1(n1102), .CO(n51986));
    SB_CARRY add_18_9 (.CI(n51475), .I0(n257[7]), .I1(n306[7]), .CO(n51476));
    SB_LUT4 add_6160_15_lut (.I0(GND_net), .I1(n14518[12]), .I2(n1029), 
            .I3(n51984), .O(n13590[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_15 (.CI(n51984), .I0(n14518[12]), .I1(n1029), .CO(n51985));
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n306[6]), .I3(n51474), 
            .O(n356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_14_lut (.I0(GND_net), .I1(n14518[11]), .I2(n956), 
            .I3(n51983), .O(n13590[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_14 (.CI(n51983), .I0(n14518[11]), .I1(n956), .CO(n51984));
    SB_LUT4 add_6407_15_lut (.I0(GND_net), .I1(n18858[12]), .I2(n1050), 
            .I3(n51757), .O(n18438[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_14_lut (.I0(GND_net), .I1(n18858[11]), .I2(n977), 
            .I3(n51756), .O(n18438[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_13_lut (.I0(GND_net), .I1(n14518[10]), .I2(n883), 
            .I3(n51982), .O(n13590[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[23]), 
            .I3(n51606), .O(n436[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_14 (.CI(n51756), .I0(n18858[11]), .I1(n977), .CO(n51757));
    SB_LUT4 add_6407_13_lut (.I0(GND_net), .I1(n18858[10]), .I2(n904), 
            .I3(n51755), .O(n18438[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_13 (.CI(n51982), .I0(n14518[10]), .I1(n883), .CO(n51983));
    SB_LUT4 add_6160_12_lut (.I0(GND_net), .I1(n14518[9]), .I2(n810), 
            .I3(n51981), .O(n13590[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_13 (.CI(n51755), .I0(n18858[10]), .I1(n904), .CO(n51756));
    SB_LUT4 add_6407_12_lut (.I0(GND_net), .I1(n18858[9]), .I2(n831), 
            .I3(n51754), .O(n18438[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[22]), 
            .I3(n51605), .O(n436[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_12 (.CI(n51754), .I0(n18858[9]), .I1(n831), .CO(n51755));
    SB_LUT4 add_6447_7_lut (.I0(GND_net), .I1(n19390[4]), .I2(n469_adj_4916), 
            .I3(n52897), .O(n19053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n51605), .I0(GND_net), .I1(n1_adj_5101[22]), 
            .CO(n51606));
    SB_CARRY add_6160_12 (.CI(n51981), .I0(n14518[9]), .I1(n810), .CO(n51982));
    SB_LUT4 add_6407_11_lut (.I0(GND_net), .I1(n18858[8]), .I2(n758), 
            .I3(n51753), .O(n18438[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[21]), 
            .I3(n51604), .O(n436[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_11 (.CI(n51753), .I0(n18858[8]), .I1(n758), .CO(n51754));
    SB_CARRY unary_minus_26_add_3_23 (.CI(n51604), .I0(GND_net), .I1(n1_adj_5101[21]), 
            .CO(n51605));
    SB_LUT4 add_6407_10_lut (.I0(GND_net), .I1(n18858[7]), .I2(n685), 
            .I3(n51752), .O(n18438[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_11_lut (.I0(GND_net), .I1(n14518[8]), .I2(n737), 
            .I3(n51980), .O(n13590[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_11 (.CI(n51980), .I0(n14518[8]), .I1(n737), .CO(n51981));
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[20]), 
            .I3(n51603), .O(n436[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_10_lut (.I0(GND_net), .I1(n14518[7]), .I2(n664), 
            .I3(n51979), .O(n13590[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_10 (.CI(n51752), .I0(n18858[7]), .I1(n685), .CO(n51753));
    SB_LUT4 add_6407_9_lut (.I0(GND_net), .I1(n18858[6]), .I2(n612), .I3(n51751), 
            .O(n18438[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_22 (.CI(n51603), .I0(GND_net), .I1(n1_adj_5101[20]), 
            .CO(n51604));
    SB_CARRY add_6407_9 (.CI(n51751), .I0(n18858[6]), .I1(n612), .CO(n51752));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[19]), 
            .I3(n51602), .O(n436[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_8 (.CI(n51474), .I0(n257[6]), .I1(n306[6]), .CO(n51475));
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n356[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5076));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6160_10 (.CI(n51979), .I0(n14518[7]), .I1(n664), .CO(n51980));
    SB_LUT4 add_6407_8_lut (.I0(GND_net), .I1(n18858[5]), .I2(n539), .I3(n51750), 
            .O(n18438[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_8 (.CI(n51750), .I0(n18858[5]), .I1(n539), .CO(n51751));
    SB_CARRY unary_minus_26_add_3_21 (.CI(n51602), .I0(GND_net), .I1(n1_adj_5101[19]), 
            .CO(n51603));
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[18]), 
            .I3(n51601), .O(n436[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_9_lut (.I0(GND_net), .I1(n14518[6]), .I2(n591), .I3(n51978), 
            .O(n13590[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_7_lut (.I0(GND_net), .I1(n18858[4]), .I2(n466), .I3(n51749), 
            .O(n18438[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_7 (.CI(n51749), .I0(n18858[4]), .I1(n466), .CO(n51750));
    SB_CARRY add_6160_9 (.CI(n51978), .I0(n14518[6]), .I1(n591), .CO(n51979));
    SB_LUT4 add_6407_6_lut (.I0(GND_net), .I1(n18858[3]), .I2(n393_adj_4911), 
            .I3(n51748), .O(n18438[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n306[5]), .I3(n51473), 
            .O(n356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_6 (.CI(n51748), .I0(n18858[3]), .I1(n393_adj_4911), 
            .CO(n51749));
    SB_LUT4 add_6160_8_lut (.I0(GND_net), .I1(n14518[5]), .I2(n518), .I3(n51977), 
            .O(n13590[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_5_lut (.I0(GND_net), .I1(n18858[2]), .I2(n320), .I3(n51747), 
            .O(n18438[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_7 (.CI(n51473), .I0(n257[5]), .I1(n306[5]), .CO(n51474));
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n306[4]), .I3(n51472), 
            .O(n356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_6 (.CI(n51472), .I0(n257[4]), .I1(n306[4]), .CO(n51473));
    SB_CARRY add_6407_5 (.CI(n51747), .I0(n18858[2]), .I1(n320), .CO(n51748));
    SB_CARRY unary_minus_26_add_3_20 (.CI(n51601), .I0(GND_net), .I1(n1_adj_5101[18]), 
            .CO(n51602));
    SB_CARRY add_6160_8 (.CI(n51977), .I0(n14518[5]), .I1(n518), .CO(n51978));
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[17]), 
            .I3(n51600), .O(n436[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_4_lut (.I0(GND_net), .I1(n18858[1]), .I2(n247), .I3(n51746), 
            .O(n18438[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_4 (.CI(n51746), .I0(n18858[1]), .I1(n247), .CO(n51747));
    SB_CARRY unary_minus_26_add_3_19 (.CI(n51600), .I0(GND_net), .I1(n1_adj_5101[17]), 
            .CO(n51601));
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[16]), 
            .I3(n51599), .O(n436[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_3_lut (.I0(GND_net), .I1(n18858[0]), .I2(n174), .I3(n51745), 
            .O(n18438[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_7 (.CI(n52897), .I0(n19390[4]), .I1(n469_adj_4916), 
            .CO(n52898));
    SB_LUT4 add_6447_6_lut (.I0(GND_net), .I1(n19390[3]), .I2(n396_adj_4908), 
            .I3(n52896), .O(n19053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_7_lut (.I0(GND_net), .I1(n14518[4]), .I2(n445_adj_4907), 
            .I3(n51976), .O(n13590[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_3 (.CI(n51745), .I0(n18858[0]), .I1(n174), .CO(n51746));
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n356[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5077));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6407_2_lut (.I0(GND_net), .I1(n32_adj_4906), .I2(n101), 
            .I3(GND_net), .O(n18438[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_18 (.CI(n51599), .I0(GND_net), .I1(n1_adj_5101[16]), 
            .CO(n51600));
    SB_CARRY add_6160_7 (.CI(n51976), .I0(n14518[4]), .I1(n445_adj_4907), 
            .CO(n51977));
    SB_CARRY add_6447_6 (.CI(n52896), .I0(n19390[3]), .I1(n396_adj_4908), 
            .CO(n52897));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[15]), 
            .I3(n51598), .O(n436[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_2 (.CI(GND_net), .I0(n32_adj_4906), .I1(n101), .CO(n51745));
    SB_LUT4 add_6561_8_lut (.I0(GND_net), .I1(n20502[5]), .I2(n560), .I3(n51744), 
            .O(n20405[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n51598), .I0(GND_net), .I1(n1_adj_5101[15]), 
            .CO(n51599));
    SB_LUT4 add_6561_7_lut (.I0(GND_net), .I1(n20502[4]), .I2(n487), .I3(n51743), 
            .O(n20405[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6447_5_lut (.I0(GND_net), .I1(n19390[2]), .I2(n323_adj_4904), 
            .I3(n52895), .O(n19053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6160_6_lut (.I0(GND_net), .I1(n14518[3]), .I2(n372_adj_4903), 
            .I3(n51975), .O(n13590[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n306[3]), .I3(n51471), 
            .O(n356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[14]), 
            .I3(n51597), .O(n436[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_6 (.CI(n51975), .I0(n14518[3]), .I1(n372_adj_4903), 
            .CO(n51976));
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n356[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5078));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6160_5_lut (.I0(GND_net), .I1(n14518[2]), .I2(n299_adj_4901), 
            .I3(n51974), .O(n13590[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6561_7 (.CI(n51743), .I0(n20502[4]), .I1(n487), .CO(n51744));
    SB_LUT4 add_6561_6_lut (.I0(GND_net), .I1(n20502[3]), .I2(n414), .I3(n51742), 
            .O(n20405[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_5 (.CI(n52895), .I0(n19390[2]), .I1(n323_adj_4904), 
            .CO(n52896));
    SB_CARRY unary_minus_26_add_3_16 (.CI(n51597), .I0(GND_net), .I1(n1_adj_5101[14]), 
            .CO(n51598));
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[13]), 
            .I3(n51596), .O(n436[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6561_6 (.CI(n51742), .I0(n20502[3]), .I1(n414), .CO(n51743));
    SB_LUT4 add_6561_5_lut (.I0(GND_net), .I1(n20502[2]), .I2(n341), .I3(n51741), 
            .O(n20405[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_15 (.CI(n51596), .I0(GND_net), .I1(n1_adj_5101[13]), 
            .CO(n51597));
    SB_LUT4 add_6447_4_lut (.I0(GND_net), .I1(n19390[1]), .I2(n250_adj_4899), 
            .I3(n52894), .O(n19053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[12]), 
            .I3(n51595), .O(n436[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_5 (.CI(n51974), .I0(n14518[2]), .I1(n299_adj_4901), 
            .CO(n51975));
    SB_CARRY add_6561_5 (.CI(n51741), .I0(n20502[2]), .I1(n341), .CO(n51742));
    SB_CARRY add_6447_4 (.CI(n52894), .I0(n19390[1]), .I1(n250_adj_4899), 
            .CO(n52895));
    SB_CARRY unary_minus_26_add_3_14 (.CI(n51595), .I0(GND_net), .I1(n1_adj_5101[12]), 
            .CO(n51596));
    SB_LUT4 add_6160_4_lut (.I0(GND_net), .I1(n14518[1]), .I2(n226_adj_4897), 
            .I3(n51973), .O(n13590[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[11]), 
            .I3(n51594), .O(n436[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6561_4_lut (.I0(GND_net), .I1(n20502[1]), .I2(n268), .I3(n51740), 
            .O(n20405[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6561_4 (.CI(n51740), .I0(n20502[1]), .I1(n268), .CO(n51741));
    SB_LUT4 add_6447_3_lut (.I0(GND_net), .I1(n19390[0]), .I2(n177_adj_4895), 
            .I3(n52893), .O(n19053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n51594), .I0(GND_net), .I1(n1_adj_5101[11]), 
            .CO(n51595));
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[10]), 
            .I3(n51593), .O(n436[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n51593), .I0(GND_net), .I1(n1_adj_5101[10]), 
            .CO(n51594));
    SB_LUT4 add_6561_3_lut (.I0(GND_net), .I1(n20502[0]), .I2(n195_adj_4893), 
            .I3(n51739), .O(n20405[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6160_4 (.CI(n51973), .I0(n14518[1]), .I1(n226_adj_4897), 
            .CO(n51974));
    SB_CARRY add_6561_3 (.CI(n51739), .I0(n20502[0]), .I1(n195_adj_4893), 
            .CO(n51740));
    SB_LUT4 add_6160_3_lut (.I0(GND_net), .I1(n14518[0]), .I2(n153_adj_4892), 
            .I3(n51972), .O(n13590[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6447_3 (.CI(n52893), .I0(n19390[0]), .I1(n177_adj_4895), 
            .CO(n52894));
    SB_CARRY add_6160_3 (.CI(n51972), .I0(n14518[0]), .I1(n153_adj_4892), 
            .CO(n51973));
    SB_LUT4 add_6561_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_4891), 
            .I3(GND_net), .O(n20405[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6561_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6561_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_4891), .CO(n51739));
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[9]), 
            .I3(n51592), .O(n436[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_11 (.CI(n51592), .I0(GND_net), .I1(n1_adj_5101[9]), 
            .CO(n51593));
    SB_LUT4 add_6447_2_lut (.I0(GND_net), .I1(n35_adj_4889), .I2(n104_adj_4888), 
            .I3(GND_net), .O(n19053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6447_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_5 (.CI(n51471), .I0(n257[3]), .I1(n306[3]), .CO(n51472));
    SB_CARRY add_6447_2 (.CI(GND_net), .I0(n35_adj_4889), .I1(n104_adj_4888), 
            .CO(n52893));
    SB_LUT4 add_6567_7_lut (.I0(GND_net), .I1(n61880), .I2(n490_adj_4884), 
            .I3(n52892), .O(n20454[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51598_4_lut (.I0(n21_adj_5078), .I1(n19_adj_5077), .I2(n17_adj_5076), 
            .I3(n9_adj_5075), .O(n67772));
    defparam i51598_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6160_2_lut (.I0(GND_net), .I1(n11_adj_4880), .I2(n80_adj_4879), 
            .I3(GND_net), .O(n13590[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6160_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_6_lut (.I0(GND_net), .I1(n20538[3]), .I2(n417_adj_4877), 
            .I3(n52891), .O(n20454[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n306[2]), .I3(n51470), 
            .O(n356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[8]), 
            .I3(n51591), .O(n436[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_10 (.CI(n51591), .I0(GND_net), .I1(n1_adj_5101[8]), 
            .CO(n51592));
    SB_CARRY add_6160_2 (.CI(GND_net), .I0(n11_adj_4880), .I1(n80_adj_4879), 
            .CO(n51972));
    SB_CARRY add_6567_6 (.CI(n52891), .I0(n20538[3]), .I1(n417_adj_4877), 
            .CO(n52892));
    SB_CARRY add_18_4 (.CI(n51470), .I0(n257[2]), .I1(n306[2]), .CO(n51471));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n306[1]), .I3(n51469), 
            .O(n379)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[7]), 
            .I3(n51590), .O(n436[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_9 (.CI(n51590), .I0(GND_net), .I1(n1_adj_5101[7]), 
            .CO(n51591));
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[6]), 
            .I3(n51589), .O(n436[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_8 (.CI(n51589), .I0(GND_net), .I1(n1_adj_5101[6]), 
            .CO(n51590));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[5]), 
            .I3(n51588), .O(n436[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_3 (.CI(n51469), .I0(n257[1]), .I1(n306[1]), .CO(n51470));
    SB_CARRY unary_minus_26_add_3_7 (.CI(n51588), .I0(GND_net), .I1(n1_adj_5101[5]), 
            .CO(n51589));
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[4]), 
            .I3(n51587), .O(n436[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n306[0]), .I3(GND_net), 
            .O(n356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_6 (.CI(n51587), .I0(GND_net), .I1(n1_adj_5101[4]), 
            .CO(n51588));
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[3]), 
            .I3(n51586), .O(n436[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n51586), .I0(GND_net), .I1(n1_adj_5101[3]), 
            .CO(n51587));
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[2]), 
            .I3(n51585), .O(n436[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n51585), .I0(GND_net), .I1(n1_adj_5101[2]), 
            .CO(n51586));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[1]), 
            .I3(n51584), .O(n436[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_5_lut (.I0(GND_net), .I1(n20538[2]), .I2(n344_adj_4867), 
            .I3(n52890), .O(n20454[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_5 (.CI(n52890), .I0(n20538[2]), .I1(n344_adj_4867), 
            .CO(n52891));
    SB_LUT4 add_6434_14_lut (.I0(GND_net), .I1(n19222[11]), .I2(n980), 
            .I3(n51729), .O(n18858[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n51584), .I0(GND_net), .I1(n1_adj_5101[1]), 
            .CO(n51585));
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n306[0]), .CO(n51469));
    SB_LUT4 add_6434_13_lut (.I0(GND_net), .I1(n19222[10]), .I2(n907), 
            .I3(n51728), .O(n18858[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_13 (.CI(n51728), .I0(n19222[10]), .I1(n907), .CO(n51729));
    SB_LUT4 add_6434_12_lut (.I0(GND_net), .I1(n19222[9]), .I2(n834), 
            .I3(n51727), .O(n18858[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_12 (.CI(n51727), .I0(n19222[9]), .I1(n834), .CO(n51728));
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5101[0]), 
            .I3(VCC_net), .O(n436[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_4_lut (.I0(GND_net), .I1(n20538[1]), .I2(n271_adj_4864), 
            .I3(n52889), .O(n20454[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n1[23]), .I3(n51468), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5101[0]), 
            .CO(n51584));
    SB_LUT4 add_6434_11_lut (.I0(GND_net), .I1(n19222[8]), .I2(n761), 
            .I3(n51726), .O(n18858[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_11 (.CI(n51726), .I0(n19222[8]), .I1(n761), .CO(n51727));
    SB_LUT4 add_6434_10_lut (.I0(GND_net), .I1(n19222[7]), .I2(n688), 
            .I3(n51725), .O(n18858[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n1[22]), .I3(n51467), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n356[23]), .I1(GND_net), .I2(n1_adj_5100[23]), 
            .I3(n51583), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[22]), 
            .I3(n51582), .O(n382[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_10 (.CI(n51725), .I0(n19222[7]), .I1(n688), .CO(n51726));
    SB_CARRY add_6567_4 (.CI(n52889), .I0(n20538[1]), .I1(n271_adj_4864), 
            .CO(n52890));
    SB_LUT4 add_6434_9_lut (.I0(GND_net), .I1(n19222[6]), .I2(n615), .I3(n51724), 
            .O(n18858[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n51582), .I0(GND_net), .I1(n1_adj_5100[22]), 
            .CO(n51583));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[21]), 
            .I3(n51581), .O(n382[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_3_lut (.I0(GND_net), .I1(n20538[0]), .I2(n198_adj_4857), 
            .I3(n52888), .O(n20454[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_9 (.CI(n51724), .I0(n19222[6]), .I1(n615), .CO(n51725));
    SB_CARRY unary_minus_20_add_3_23 (.CI(n51581), .I0(GND_net), .I1(n1_adj_5100[21]), 
            .CO(n51582));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[20]), 
            .I3(n51580), .O(n382[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_3 (.CI(n52888), .I0(n20538[0]), .I1(n198_adj_4857), 
            .CO(n52889));
    SB_LUT4 add_6434_8_lut (.I0(GND_net), .I1(n19222[5]), .I2(n542), .I3(n51723), 
            .O(n18858[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n51580), .I0(GND_net), .I1(n1_adj_5100[20]), 
            .CO(n51581));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[19]), 
            .I3(n51579), .O(n382[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_2_lut (.I0(GND_net), .I1(n56_adj_4853), .I2(n125_adj_4852), 
            .I3(GND_net), .O(n20454[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_8 (.CI(n51723), .I0(n19222[5]), .I1(n542), .CO(n51724));
    SB_LUT4 add_6434_7_lut (.I0(GND_net), .I1(n19222[4]), .I2(n469), .I3(n51722), 
            .O(n18858[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n51579), .I0(GND_net), .I1(n1_adj_5100[19]), 
            .CO(n51580));
    SB_CARRY add_6434_7 (.CI(n51722), .I0(n19222[4]), .I1(n469), .CO(n51723));
    SB_CARRY add_9_24 (.CI(n51467), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n1[22]), .CO(n51468));
    SB_LUT4 add_6434_6_lut (.I0(GND_net), .I1(n19222[3]), .I2(n396_adj_4849), 
            .I3(n51721), .O(n18858[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[18]), 
            .I3(n51578), .O(n382[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_2 (.CI(GND_net), .I0(n56_adj_4853), .I1(n125_adj_4852), 
            .CO(n52888));
    SB_CARRY add_6434_6 (.CI(n51721), .I0(n19222[3]), .I1(n396_adj_4849), 
            .CO(n51722));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n51578), .I0(GND_net), .I1(n1_adj_5100[18]), 
            .CO(n51579));
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n1[21]), .I3(n51466), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[17]), 
            .I3(n51577), .O(n382[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6434_5_lut (.I0(GND_net), .I1(n19222[2]), .I2(n323), .I3(n51720), 
            .O(n18858[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6471_13_lut (.I0(GND_net), .I1(n19677[10]), .I2(n910_adj_4842), 
            .I3(n52887), .O(n19390[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n51466), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n1[21]), .CO(n51467));
    SB_LUT4 add_6471_12_lut (.I0(GND_net), .I1(n19677[9]), .I2(n837_adj_4841), 
            .I3(n52886), .O(n19390[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_12 (.CI(n52886), .I0(n19677[9]), .I1(n837_adj_4841), 
            .CO(n52887));
    SB_LUT4 add_6471_11_lut (.I0(GND_net), .I1(n19677[8]), .I2(n764_adj_4836), 
            .I3(n52885), .O(n19390[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n51577), .I0(GND_net), .I1(n1_adj_5100[17]), 
            .CO(n51578));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[16]), 
            .I3(n51576), .O(n382[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_11 (.CI(n52885), .I0(n19677[8]), .I1(n764_adj_4836), 
            .CO(n52886));
    SB_LUT4 add_6471_10_lut (.I0(GND_net), .I1(n19677[7]), .I2(n691_adj_4831), 
            .I3(n52884), .O(n19390[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_5 (.CI(n51720), .I0(n19222[2]), .I1(n323), .CO(n51721));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n51576), .I0(GND_net), .I1(n1_adj_5100[16]), 
            .CO(n51577));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[15]), 
            .I3(n51575), .O(n382[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_10 (.CI(n52884), .I0(n19677[7]), .I1(n691_adj_4831), 
            .CO(n52885));
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n1[20]), .I3(n51465), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6434_4_lut (.I0(GND_net), .I1(n19222[1]), .I2(n250), .I3(n51719), 
            .O(n18858[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n51575), .I0(GND_net), .I1(n1_adj_5100[15]), 
            .CO(n51576));
    SB_CARRY add_6434_4 (.CI(n51719), .I0(n19222[1]), .I1(n250), .CO(n51720));
    SB_CARRY add_9_22 (.CI(n51465), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n1[20]), .CO(n51466));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[14]), 
            .I3(n51574), .O(n382[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6471_9_lut (.I0(GND_net), .I1(n19677[6]), .I2(n618_adj_4827), 
            .I3(n52883), .O(n19390[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6434_3_lut (.I0(GND_net), .I1(n19222[0]), .I2(n177), .I3(n51718), 
            .O(n18858[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_3 (.CI(n51718), .I0(n19222[0]), .I1(n177), .CO(n51719));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n51574), .I0(GND_net), .I1(n1_adj_5100[14]), 
            .CO(n51575));
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n1[19]), .I3(n51464), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[13]), 
            .I3(n51573), .O(n382[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6434_2_lut (.I0(GND_net), .I1(n35_adj_4823), .I2(n104), 
            .I3(GND_net), .O(n18858[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6434_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_9 (.CI(n52883), .I0(n19677[6]), .I1(n618_adj_4827), 
            .CO(n52884));
    SB_CARRY unary_minus_20_add_3_15 (.CI(n51573), .I0(GND_net), .I1(n1_adj_5100[13]), 
            .CO(n51574));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[12]), 
            .I3(n51572), .O(n382[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6434_2 (.CI(GND_net), .I0(n35_adj_4823), .I1(n104), .CO(n51718));
    SB_CARRY add_9_21 (.CI(n51464), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n1[19]), .CO(n51465));
    SB_LUT4 add_6471_8_lut (.I0(GND_net), .I1(n19677[5]), .I2(n545_adj_4820), 
            .I3(n52882), .O(n19390[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n1[18]), .I3(n51463), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n51572), .I0(GND_net), .I1(n1_adj_5100[12]), 
            .CO(n51573));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[11]), 
            .I3(n51571), .O(n382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6203_21_lut (.I0(GND_net), .I1(n15358[18]), .I2(GND_net), 
            .I3(n51955), .O(n14518[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_8 (.CI(n52882), .I0(n19677[5]), .I1(n545_adj_4820), 
            .CO(n52883));
    SB_LUT4 add_6471_7_lut (.I0(GND_net), .I1(n19677[4]), .I2(n472_adj_4816), 
            .I3(n52881), .O(n19390[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n51463), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n1[18]), .CO(n51464));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n1[17]), .I3(n51462), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n51571), .I0(GND_net), .I1(n1_adj_5100[11]), 
            .CO(n51572));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[10]), 
            .I3(n51570), .O(n382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6203_20_lut (.I0(GND_net), .I1(n15358[17]), .I2(GND_net), 
            .I3(n51954), .O(n14518[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n51570), .I0(GND_net), .I1(n1_adj_5100[10]), 
            .CO(n51571));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[9]), 
            .I3(n51569), .O(n382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_20 (.CI(n51954), .I0(n15358[17]), .I1(GND_net), 
            .CO(n51955));
    SB_CARRY unary_minus_20_add_3_11 (.CI(n51569), .I0(GND_net), .I1(n1_adj_5100[9]), 
            .CO(n51570));
    SB_LUT4 add_6203_19_lut (.I0(GND_net), .I1(n15358[16]), .I2(GND_net), 
            .I3(n51953), .O(n14518[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_19 (.CI(n51953), .I0(n15358[16]), .I1(GND_net), 
            .CO(n51954));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[8]), 
            .I3(n51568), .O(n382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n51462), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n1[17]), .CO(n51463));
    SB_LUT4 add_6203_18_lut (.I0(GND_net), .I1(n15358[15]), .I2(GND_net), 
            .I3(n51952), .O(n14518[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n1[16]), .I3(n51461), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_18 (.CI(n51952), .I0(n15358[15]), .I1(GND_net), 
            .CO(n51953));
    SB_LUT4 add_6203_17_lut (.I0(GND_net), .I1(n15358[14]), .I2(GND_net), 
            .I3(n51951), .O(n14518[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n51568), .I0(GND_net), .I1(n1_adj_5100[8]), 
            .CO(n51569));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[7]), 
            .I3(n51567), .O(n382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51584_4_lut (.I0(n27_adj_5074), .I1(n15_adj_5073), .I2(n13_adj_5072), 
            .I3(n11_adj_5071), .O(n67758));
    defparam i51584_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n51567), .I0(GND_net), .I1(n1_adj_5100[7]), 
            .CO(n51568));
    SB_CARRY add_6203_17 (.CI(n51951), .I0(n15358[14]), .I1(GND_net), 
            .CO(n51952));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[6]), 
            .I3(n51566), .O(n382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6203_16_lut (.I0(GND_net), .I1(n15358[13]), .I2(n1105_adj_4803), 
            .I3(n51950), .O(n14518[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n51566), .I0(GND_net), .I1(n1_adj_5100[6]), 
            .CO(n51567));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[5]), 
            .I3(n51565), .O(n382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_16 (.CI(n51950), .I0(n15358[13]), .I1(n1105_adj_4803), 
            .CO(n51951));
    SB_CARRY unary_minus_20_add_3_7 (.CI(n51565), .I0(GND_net), .I1(n1_adj_5100[5]), 
            .CO(n51566));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[4]), 
            .I3(n51564), .O(n382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n51564), .I0(GND_net), .I1(n1_adj_5100[4]), 
            .CO(n51565));
    SB_LUT4 add_6203_15_lut (.I0(GND_net), .I1(n15358[12]), .I2(n1032_adj_4800), 
            .I3(n51949), .O(n14518[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_15 (.CI(n51949), .I0(n15358[12]), .I1(n1032_adj_4800), 
            .CO(n51950));
    SB_LUT4 add_6203_14_lut (.I0(GND_net), .I1(n15358[11]), .I2(n959_adj_4799), 
            .I3(n51948), .O(n14518[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[3]), 
            .I3(n51563), .O(n382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_14 (.CI(n51948), .I0(n15358[11]), .I1(n959_adj_4799), 
            .CO(n51949));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n51563), .I0(GND_net), .I1(n1_adj_5100[3]), 
            .CO(n51564));
    SB_LUT4 add_6459_13_lut (.I0(GND_net), .I1(n19534[10]), .I2(n910), 
            .I3(n51709), .O(n19222[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6203_13_lut (.I0(GND_net), .I1(n15358[10]), .I2(n886_adj_4795), 
            .I3(n51947), .O(n14518[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_7 (.CI(n52881), .I0(n19677[4]), .I1(n472_adj_4816), 
            .CO(n52882));
    SB_LUT4 add_6471_6_lut (.I0(GND_net), .I1(n19677[3]), .I2(n399_adj_4794), 
            .I3(n52880), .O(n19390[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_13 (.CI(n51947), .I0(n15358[10]), .I1(n886_adj_4795), 
            .CO(n51948));
    SB_LUT4 add_6203_12_lut (.I0(GND_net), .I1(n15358[9]), .I2(n813_adj_4793), 
            .I3(n51946), .O(n14518[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_12 (.CI(n51946), .I0(n15358[9]), .I1(n813_adj_4793), 
            .CO(n51947));
    SB_LUT4 add_6203_11_lut (.I0(GND_net), .I1(n15358[8]), .I2(n740_adj_4792), 
            .I3(n51945), .O(n14518[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_11 (.CI(n51945), .I0(n15358[8]), .I1(n740_adj_4792), 
            .CO(n51946));
    SB_LUT4 add_6203_10_lut (.I0(GND_net), .I1(n15358[7]), .I2(n667_adj_4791), 
            .I3(n51944), .O(n14518[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_10 (.CI(n51944), .I0(n15358[7]), .I1(n667_adj_4791), 
            .CO(n51945));
    SB_LUT4 add_6203_9_lut (.I0(GND_net), .I1(n15358[6]), .I2(n594_adj_4789), 
            .I3(n51943), .O(n14518[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_18 (.CI(n51461), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n1[16]), .CO(n51462));
    SB_CARRY add_6471_6 (.CI(n52880), .I0(n19677[3]), .I1(n399_adj_4794), 
            .CO(n52881));
    SB_CARRY add_6203_9 (.CI(n51943), .I0(n15358[6]), .I1(n594_adj_4789), 
            .CO(n51944));
    SB_LUT4 add_6203_8_lut (.I0(GND_net), .I1(n15358[5]), .I2(n521_adj_4788), 
            .I3(n51942), .O(n14518[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_8 (.CI(n51942), .I0(n15358[5]), .I1(n521_adj_4788), 
            .CO(n51943));
    SB_LUT4 add_6203_7_lut (.I0(GND_net), .I1(n15358[4]), .I2(n448_adj_4785), 
            .I3(n51941), .O(n14518[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[2]), 
            .I3(n51562), .O(n382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_7 (.CI(n51941), .I0(n15358[4]), .I1(n448_adj_4785), 
            .CO(n51942));
    SB_LUT4 add_6203_6_lut (.I0(GND_net), .I1(n15358[3]), .I2(n375_adj_4781), 
            .I3(n51940), .O(n14518[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_6 (.CI(n51940), .I0(n15358[3]), .I1(n375_adj_4781), 
            .CO(n51941));
    SB_LUT4 add_6203_5_lut (.I0(GND_net), .I1(n15358[2]), .I2(n302_adj_4780), 
            .I3(n51939), .O(n14518[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_5 (.CI(n51939), .I0(n15358[2]), .I1(n302_adj_4780), 
            .CO(n51940));
    SB_LUT4 add_6471_5_lut (.I0(GND_net), .I1(n19677[2]), .I2(n326_adj_4779), 
            .I3(n52879), .O(n19390[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6471_5 (.CI(n52879), .I0(n19677[2]), .I1(n326_adj_4779), 
            .CO(n52880));
    SB_LUT4 add_6471_4_lut (.I0(GND_net), .I1(n19677[1]), .I2(n253_adj_4778), 
            .I3(n52878), .O(n19390[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n51562), .I0(GND_net), .I1(n1_adj_5100[2]), 
            .CO(n51563));
    SB_CARRY add_6471_4 (.CI(n52878), .I0(n19677[1]), .I1(n253_adj_4778), 
            .CO(n52879));
    SB_LUT4 add_6203_4_lut (.I0(GND_net), .I1(n15358[1]), .I2(n229_adj_4777), 
            .I3(n51938), .O(n14518[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_4 (.CI(n51938), .I0(n15358[1]), .I1(n229_adj_4777), 
            .CO(n51939));
    SB_LUT4 add_6471_3_lut (.I0(GND_net), .I1(n19677[0]), .I2(n180_adj_4775), 
            .I3(n52877), .O(n19390[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5100[1]), 
            .I3(n51561), .O(n405)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6203_3_lut (.I0(GND_net), .I1(n15358[0]), .I2(n156_adj_4770), 
            .I3(n51937), .O(n14518[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6203_3 (.CI(n51937), .I0(n15358[0]), .I1(n156_adj_4770), 
            .CO(n51938));
    SB_CARRY add_6471_3 (.CI(n52877), .I0(n19677[0]), .I1(n180_adj_4775), 
            .CO(n52878));
    SB_LUT4 add_6203_2_lut (.I0(GND_net), .I1(n14_adj_4769), .I2(n83_adj_4768), 
            .I3(GND_net), .O(n14518[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6203_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6471_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_4767), 
            .I3(GND_net), .O(n19390[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6471_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6459_12_lut (.I0(GND_net), .I1(n19534[9]), .I2(n837), 
            .I3(n51708), .O(n19222[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_12 (.CI(n51708), .I0(n19534[9]), .I1(n837), .CO(n51709));
    SB_CARRY add_6471_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_4767), .CO(n52877));
    SB_CARRY add_6203_2 (.CI(GND_net), .I0(n14_adj_4769), .I1(n83_adj_4768), 
            .CO(n51937));
    SB_LUT4 add_6513_11_lut (.I0(GND_net), .I1(n20117[8]), .I2(n770), 
            .I3(n51936), .O(n19918[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_12_lut (.I0(GND_net), .I1(n19918[9]), .I2(n840_adj_4766), 
            .I3(n52876), .O(n19677[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6513_10_lut (.I0(GND_net), .I1(n20117[7]), .I2(n697), 
            .I3(n51935), .O(n19918[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_11_lut (.I0(GND_net), .I1(n19918[8]), .I2(n767_adj_4765), 
            .I3(n52875), .O(n19677[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_10 (.CI(n51935), .I0(n20117[7]), .I1(n697), .CO(n51936));
    SB_LUT4 add_6459_11_lut (.I0(GND_net), .I1(n19534[8]), .I2(n764), 
            .I3(n51707), .O(n19222[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_11 (.CI(n52875), .I0(n19918[8]), .I1(n767_adj_4765), 
            .CO(n52876));
    SB_LUT4 add_6513_9_lut (.I0(GND_net), .I1(n20117[6]), .I2(n624), .I3(n51934), 
            .O(n19918[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_10_lut (.I0(GND_net), .I1(n19918[7]), .I2(n694_adj_4763), 
            .I3(n52874), .O(n19677[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_10 (.CI(n52874), .I0(n19918[7]), .I1(n694_adj_4763), 
            .CO(n52875));
    SB_CARRY add_6513_9 (.CI(n51934), .I0(n20117[6]), .I1(n624), .CO(n51935));
    SB_LUT4 add_6513_8_lut (.I0(GND_net), .I1(n20117[5]), .I2(n551), .I3(n51933), 
            .O(n19918[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_9_lut (.I0(GND_net), .I1(n19918[6]), .I2(n621_adj_4762), 
            .I3(n52873), .O(n19677[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_8 (.CI(n51933), .I0(n20117[5]), .I1(n551), .CO(n51934));
    SB_LUT4 add_6513_7_lut (.I0(GND_net), .I1(n20117[4]), .I2(n478), .I3(n51932), 
            .O(n19918[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_9 (.CI(n52873), .I0(n19918[6]), .I1(n621_adj_4762), 
            .CO(n52874));
    SB_CARRY add_6513_7 (.CI(n51932), .I0(n20117[4]), .I1(n478), .CO(n51933));
    SB_CARRY add_6459_11 (.CI(n51707), .I0(n19534[8]), .I1(n764), .CO(n51708));
    SB_LUT4 add_6493_8_lut (.I0(GND_net), .I1(n19918[5]), .I2(n548_adj_4759), 
            .I3(n52872), .O(n19677[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6459_10_lut (.I0(GND_net), .I1(n19534[7]), .I2(n691), 
            .I3(n51706), .O(n19222[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6513_6_lut (.I0(GND_net), .I1(n20117[3]), .I2(n405_c), 
            .I3(n51931), .O(n19918[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_6 (.CI(n51931), .I0(n20117[3]), .I1(n405_c), .CO(n51932));
    SB_LUT4 add_6513_5_lut (.I0(GND_net), .I1(n20117[2]), .I2(n332_adj_4755), 
            .I3(n51930), .O(n19918[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_10 (.CI(n51706), .I0(n19534[7]), .I1(n691), .CO(n51707));
    SB_CARRY add_6493_8 (.CI(n52872), .I0(n19918[5]), .I1(n548_adj_4759), 
            .CO(n52873));
    SB_LUT4 add_6459_9_lut (.I0(GND_net), .I1(n19534[6]), .I2(n618), .I3(n51705), 
            .O(n19222[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_5 (.CI(n51930), .I0(n20117[2]), .I1(n332_adj_4755), 
            .CO(n51931));
    SB_CARRY unary_minus_20_add_3_3 (.CI(n51561), .I0(GND_net), .I1(n1_adj_5100[1]), 
            .CO(n51562));
    SB_LUT4 add_6513_4_lut (.I0(GND_net), .I1(n20117[1]), .I2(n259_adj_4754), 
            .I3(n51929), .O(n19918[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n37361), .I1(GND_net), .I2(n1_adj_5100[0]), 
            .I3(VCC_net), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_6513_4 (.CI(n51929), .I0(n20117[1]), .I1(n259_adj_4754), 
            .CO(n51930));
    SB_CARRY add_6459_9 (.CI(n51705), .I0(n19534[6]), .I1(n618), .CO(n51706));
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5100[0]), 
            .CO(n51561));
    SB_LUT4 add_6513_3_lut (.I0(GND_net), .I1(n20117[0]), .I2(n186_adj_4752), 
            .I3(n51928), .O(n19918[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[23]), 
            .I3(n51560), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_3 (.CI(n51928), .I0(n20117[0]), .I1(n186_adj_4752), 
            .CO(n51929));
    SB_LUT4 add_6513_2_lut (.I0(GND_net), .I1(n44_adj_4751), .I2(n113_adj_4750), 
            .I3(GND_net), .O(n19918[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6513_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6513_2 (.CI(GND_net), .I0(n44_adj_4751), .I1(n113_adj_4750), 
            .CO(n51928));
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[22]), 
            .I3(n51559), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_7_lut (.I0(GND_net), .I1(n19918[4]), .I2(n475_adj_4749), 
            .I3(n52871), .O(n19677[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6459_8_lut (.I0(GND_net), .I1(n19534[5]), .I2(n545), .I3(n51704), 
            .O(n19222[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n1[15]), .I3(n51460), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_24 (.CI(n51559), .I0(GND_net), .I1(n1_adj_5099[22]), 
            .CO(n51560));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[21]), 
            .I3(n51558), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_8 (.CI(n51704), .I0(n19534[5]), .I1(n545), .CO(n51705));
    SB_LUT4 add_6459_7_lut (.I0(GND_net), .I1(n19534[4]), .I2(n472), .I3(n51703), 
            .O(n19222[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_7 (.CI(n52871), .I0(n19918[4]), .I1(n475_adj_4749), 
            .CO(n52872));
    SB_CARRY add_6459_7 (.CI(n51703), .I0(n19534[4]), .I1(n472), .CO(n51704));
    SB_CARRY unary_minus_13_add_3_23 (.CI(n51558), .I0(GND_net), .I1(n1_adj_5099[21]), 
            .CO(n51559));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[20]), 
            .I3(n51557), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n51557), .I0(GND_net), .I1(n1_adj_5099[20]), 
            .CO(n51558));
    SB_LUT4 add_6459_6_lut (.I0(GND_net), .I1(n19534[3]), .I2(n399), .I3(n51702), 
            .O(n19222[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_6 (.CI(n51702), .I0(n19534[3]), .I1(n399), .CO(n51703));
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[19]), 
            .I3(n51556), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_21 (.CI(n51556), .I0(GND_net), .I1(n1_adj_5099[19]), 
            .CO(n51557));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[18]), 
            .I3(n51555), .O(n188)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n51555), .I0(GND_net), .I1(n1_adj_5099[18]), 
            .CO(n51556));
    SB_LUT4 add_6459_5_lut (.I0(GND_net), .I1(n19534[2]), .I2(n326), .I3(n51701), 
            .O(n19222[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[17]), 
            .I3(n51554), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_5 (.CI(n51701), .I0(n19534[2]), .I1(n326), .CO(n51702));
    SB_LUT4 add_6493_6_lut (.I0(GND_net), .I1(n19918[3]), .I2(n402_adj_4743), 
            .I3(n52870), .O(n19677[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_19 (.CI(n51554), .I0(GND_net), .I1(n1_adj_5099[17]), 
            .CO(n51555));
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[16]), 
            .I3(n51553), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_18 (.CI(n51553), .I0(GND_net), .I1(n1_adj_5099[16]), 
            .CO(n51554));
    SB_CARRY add_6493_6 (.CI(n52870), .I0(n19918[3]), .I1(n402_adj_4743), 
            .CO(n52871));
    SB_LUT4 add_6459_4_lut (.I0(GND_net), .I1(n19534[1]), .I2(n253), .I3(n51700), 
            .O(n19222[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[15]), 
            .I3(n51552), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_5_lut (.I0(GND_net), .I1(n19918[2]), .I2(n329), .I3(n52869), 
            .O(n19677[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_4 (.CI(n51700), .I0(n19534[1]), .I1(n253), .CO(n51701));
    SB_CARRY unary_minus_13_add_3_17 (.CI(n51552), .I0(GND_net), .I1(n1_adj_5099[15]), 
            .CO(n51553));
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[14]), 
            .I3(n51551), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_5 (.CI(n52869), .I0(n19918[2]), .I1(n329), .CO(n52870));
    SB_CARRY unary_minus_13_add_3_16 (.CI(n51551), .I0(GND_net), .I1(n1_adj_5099[14]), 
            .CO(n51552));
    SB_LUT4 add_6459_3_lut (.I0(GND_net), .I1(n19534[0]), .I2(n180), .I3(n51699), 
            .O(n19222[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_4_lut (.I0(GND_net), .I1(n19918[1]), .I2(n256), .I3(n52868), 
            .O(n19677[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6459_3 (.CI(n51699), .I0(n19534[0]), .I1(n180), .CO(n51700));
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[13]), 
            .I3(n51550), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_15 (.CI(n51550), .I0(GND_net), .I1(n1_adj_5099[13]), 
            .CO(n51551));
    SB_CARRY add_6493_4 (.CI(n52868), .I0(n19918[1]), .I1(n256), .CO(n52869));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[12]), 
            .I3(n51549), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6459_2_lut (.I0(GND_net), .I1(n38_adj_4734), .I2(n107_adj_4733), 
            .I3(GND_net), .O(n19222[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6459_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_3_lut (.I0(GND_net), .I1(n19918[0]), .I2(n183), .I3(n52867), 
            .O(n19677[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n51549), .I0(GND_net), .I1(n1_adj_5099[12]), 
            .CO(n51550));
    SB_CARRY add_6459_2 (.CI(GND_net), .I0(n38_adj_4734), .I1(n107_adj_4733), 
            .CO(n51699));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[11]), 
            .I3(n51548), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_13 (.CI(n51548), .I0(GND_net), .I1(n1_adj_5099[11]), 
            .CO(n51549));
    SB_CARRY add_6493_3 (.CI(n52867), .I0(n19918[0]), .I1(n183), .CO(n52868));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[10]), 
            .I3(n51547), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6573_7_lut (.I0(GND_net), .I1(n61143), .I2(n490), .I3(n51698), 
            .O(n20502[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6493_2_lut (.I0(GND_net), .I1(n41_adj_4711), .I2(n110), 
            .I3(GND_net), .O(n19677[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6493_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_12 (.CI(n51547), .I0(GND_net), .I1(n1_adj_5099[10]), 
            .CO(n51548));
    SB_LUT4 add_6573_6_lut (.I0(GND_net), .I1(n20573[3]), .I2(n417), .I3(n51697), 
            .O(n20502[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[9]), 
            .I3(n51546), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6493_2 (.CI(GND_net), .I0(n41_adj_4711), .I1(n110), .CO(n52867));
    SB_CARRY unary_minus_13_add_3_11 (.CI(n51546), .I0(GND_net), .I1(n1_adj_5099[9]), 
            .CO(n51547));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[8]), 
            .I3(n51545), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6573_6 (.CI(n51697), .I0(n20573[3]), .I1(n417), .CO(n51698));
    SB_LUT4 add_6573_5_lut (.I0(GND_net), .I1(n20576), .I2(n344), .I3(n51696), 
            .O(n20502[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n51545), .I0(GND_net), .I1(n1_adj_5099[8]), 
            .CO(n51546));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[7]), 
            .I3(n51544), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n51544), .I0(GND_net), .I1(n1_adj_5099[7]), 
            .CO(n51545));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[6]), 
            .I3(n51543), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6573_5 (.CI(n51696), .I0(n20576), .I1(n344), .CO(n51697));
    SB_CARRY unary_minus_13_add_3_8 (.CI(n51543), .I0(GND_net), .I1(n1_adj_5099[6]), 
            .CO(n51544));
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[5]), 
            .I3(n51542), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[2] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n356[7]), .I1(n356[16]), .I2(n33_adj_5070), 
            .I3(GND_net), .O(n12_adj_5086));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n356[5]), .I1(n356[6]), .I2(n13_adj_5072), 
            .I3(GND_net), .O(n10_adj_5087));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i30_3_lut (.I0(n12_adj_5086), .I1(n356[17]), .I2(n35_adj_5069), 
            .I3(GND_net), .O(n30_adj_5088));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_13_add_3_7 (.CI(n51542), .I0(GND_net), .I1(n1_adj_5099[5]), 
            .CO(n51543));
    SB_CARRY add_9_17 (.CI(n51460), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n1[15]), .CO(n51461));
    SB_LUT4 i52484_4_lut (.I0(n13_adj_5072), .I1(n11_adj_5071), .I2(n9_adj_5075), 
            .I3(n67793), .O(n68658));
    defparam i52484_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52476_4_lut (.I0(n19_adj_5077), .I1(n17_adj_5076), .I2(n15_adj_5073), 
            .I3(n68658), .O(n68650));
    defparam i52476_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n1[14]), .I3(n51459), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53476_4_lut (.I0(n25_adj_5065), .I1(n23_adj_5063), .I2(n21_adj_5078), 
            .I3(n68650), .O(n69651));
    defparam i53476_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52868_4_lut (.I0(n31_adj_5067), .I1(n29_adj_5066), .I2(n27_adj_5074), 
            .I3(n69651), .O(n69043));
    defparam i52868_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[1] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53569_4_lut (.I0(n37_adj_5068), .I1(n35_adj_5069), .I2(n33_adj_5070), 
            .I3(n69043), .O(n69744));
    defparam i53569_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n356[9]), .I1(n356[21]), .I2(n43_adj_5062), 
            .I3(GND_net), .O(n16_adj_5089));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53137_3_lut (.I0(n6_adj_5090), .I1(n356[10]), .I2(n21_adj_5078), 
            .I3(GND_net), .O(n69312));   // verilog/motorControl.v(52[14:29])
    defparam i53137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53138_3_lut (.I0(n69312), .I1(n356[11]), .I2(n23_adj_5063), 
            .I3(GND_net), .O(n69313));   // verilog/motorControl.v(52[14:29])
    defparam i53138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n356[4]), .I1(n356[8]), .I2(n17_adj_5076), 
            .I3(GND_net), .O(n8_adj_5091));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i24_3_lut (.I0(n16_adj_5089), .I1(n356[22]), .I2(n45_adj_5061), 
            .I3(GND_net), .O(n24_adj_5092));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51559_4_lut (.I0(n43_adj_5062), .I1(n25_adj_5065), .I2(n23_adj_5063), 
            .I3(n67772), .O(n67733));
    defparam i51559_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53002_4_lut (.I0(n24_adj_5092), .I1(n8_adj_5091), .I2(n45_adj_5061), 
            .I3(n67731), .O(n69177));   // verilog/motorControl.v(52[14:29])
    defparam i53002_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52026_3_lut (.I0(n69313), .I1(n356[12]), .I2(n25_adj_5065), 
            .I3(GND_net), .O(n68200));   // verilog/motorControl.v(52[14:29])
    defparam i52026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i4_4_lut (.I0(PWMLimit[0]), .I1(n379), .I2(PWMLimit[1]), 
            .I3(n356[0]), .O(n4_adj_5093));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_6573_4_lut (.I0(GND_net), .I1(n20577), .I2(n271), .I3(n51695), 
            .O(n20502[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6573_4 (.CI(n51695), .I0(n20577), .I1(n271), .CO(n51696));
    SB_LUT4 i53127_3_lut (.I0(n4_adj_5093), .I1(n356[13]), .I2(n27_adj_5074), 
            .I3(GND_net), .O(n69302));   // verilog/motorControl.v(52[14:29])
    defparam i53127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53128_3_lut (.I0(n69302), .I1(n356[14]), .I2(n29_adj_5066), 
            .I3(GND_net), .O(n69303));   // verilog/motorControl.v(52[14:29])
    defparam i53128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51576_4_lut (.I0(n33_adj_5070), .I1(n31_adj_5067), .I2(n29_adj_5066), 
            .I3(n67758), .O(n67750));
    defparam i51576_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53422_4_lut (.I0(n30_adj_5088), .I1(n10_adj_5087), .I2(n35_adj_5069), 
            .I3(n67744), .O(n69597));   // verilog/motorControl.v(52[14:29])
    defparam i53422_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52028_3_lut (.I0(n69303), .I1(n356[15]), .I2(n31_adj_5067), 
            .I3(GND_net), .O(n68202));   // verilog/motorControl.v(52[14:29])
    defparam i52028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53638_4_lut (.I0(n68202), .I1(n69597), .I2(n35_adj_5069), 
            .I3(n67750), .O(n69813));   // verilog/motorControl.v(52[14:29])
    defparam i53638_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53639_3_lut (.I0(n69813), .I1(n356[18]), .I2(n37_adj_5068), 
            .I3(GND_net), .O(n69814));   // verilog/motorControl.v(52[14:29])
    defparam i53639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53614_3_lut (.I0(n69814), .I1(n356[19]), .I2(n39_adj_5059), 
            .I3(GND_net), .O(n69789));   // verilog/motorControl.v(52[14:29])
    defparam i53614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51561_4_lut (.I0(n43_adj_5062), .I1(n41_adj_5060), .I2(n39_adj_5059), 
            .I3(n69744), .O(n67735));
    defparam i51561_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53311_4_lut (.I0(n68200), .I1(n69177), .I2(n45_adj_5061), 
            .I3(n67733), .O(n69486));   // verilog/motorControl.v(52[14:29])
    defparam i53311_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52034_3_lut (.I0(n69789), .I1(n356[20]), .I2(n41_adj_5060), 
            .I3(GND_net), .O(n68208));   // verilog/motorControl.v(52[14:29])
    defparam i52034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53522_4_lut (.I0(n68208), .I1(n69486), .I2(n45_adj_5061), 
            .I3(n67735), .O(n69697));   // verilog/motorControl.v(52[14:29])
    defparam i53522_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_9_16 (.CI(n51459), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n1[14]), .CO(n51460));
    SB_LUT4 add_6573_3_lut (.I0(GND_net), .I1(n20573[0]), .I2(n198), .I3(n51694), 
            .O(n20502[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6573_3 (.CI(n51694), .I0(n20573[0]), .I1(n198), .CO(n51695));
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[4]), 
            .I3(n51541), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6573_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_4700), 
            .I3(GND_net), .O(n20502[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6573_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53523_3_lut (.I0(n69697), .I1(PWMLimit[23]), .I2(n356[23]), 
            .I3(GND_net), .O(n409));   // verilog/motorControl.v(52[14:29])
    defparam i53523_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n51541), .I0(GND_net), .I1(n1_adj_5099[4]), 
            .CO(n51542));
    SB_LUT4 i51671_4_lut (.I0(n356[6]), .I1(n356[5]), .I2(n382[6]), .I3(n382[5]), 
            .O(n67845));
    defparam i51671_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i52531_3_lut (.I0(n356[7]), .I1(n67845), .I2(n382[7]), .I3(GND_net), 
            .O(n68706));
    defparam i52531_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i27_rep_148_2_lut (.I0(n356[13]), .I1(n382[13]), 
            .I2(GND_net), .I3(GND_net), .O(n71257));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i27_rep_148_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52515_4_lut (.I0(n356[14]), .I1(n71257), .I2(n382[14]), .I3(n68706), 
            .O(n68690));
    defparam i52515_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_142_2_lut (.I0(n356[15]), .I1(n382[15]), 
            .I2(GND_net), .I3(GND_net), .O(n71251));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i31_rep_142_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6573_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_4700), .CO(n51694));
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n382[7]), .I1(n382[16]), .I2(n356[16]), 
            .I3(GND_net), .O(n12_adj_5095));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51641_4_lut (.I0(n356[16]), .I1(n356[7]), .I2(n382[16]), 
            .I3(n382[7]), .O(n67815));
    defparam i51641_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n382[5]), .I1(n382[6]), .I2(n356[6]), 
            .I3(GND_net), .O(n10_adj_4563));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_5095), .I1(n382[17]), .I2(n356[17]), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51663_4_lut (.I0(n356[8]), .I1(n356[4]), .I2(n382[8]), .I3(n382[4]), 
            .O(n67837));
    defparam i51663_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i52527_3_lut (.I0(n356[9]), .I1(n67837), .I2(n382[9]), .I3(GND_net), 
            .O(n68702));
    defparam i52527_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i21_rep_161_2_lut (.I0(n356[10]), .I1(n382[10]), 
            .I2(GND_net), .I3(GND_net), .O(n71270));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i21_rep_161_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52523_4_lut (.I0(n356[11]), .I1(n71270), .I2(n382[11]), .I3(n68702), 
            .O(n68698));
    defparam i52523_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i25_rep_156_2_lut (.I0(n356[12]), .I1(n382[12]), 
            .I2(GND_net), .I3(GND_net), .O(n71265));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i25_rep_156_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n382[9]), .I1(n382[21]), .I2(n356[21]), 
            .I3(GND_net), .O(n16_adj_5096));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51625_4_lut (.I0(n356[21]), .I1(n356[9]), .I2(n382[21]), 
            .I3(n382[9]), .O(n67799));
    defparam i51625_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n382[4]), .I1(n382[8]), .I2(n356[8]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_5096), .I1(n382[22]), .I2(n356[22]), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51675_4_lut (.I0(n356[3]), .I1(n356[2]), .I2(n382[3]), .I3(n382[2]), 
            .O(n67849));
    defparam i51675_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i9_rep_187_2_lut (.I0(n356[4]), .I1(n382[4]), .I2(GND_net), 
            .I3(GND_net), .O(n71296));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i9_rep_187_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51673_4_lut (.I0(n356[5]), .I1(n71296), .I2(n382[5]), .I3(n67849), 
            .O(n67847));
    defparam i51673_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i13_rep_180_2_lut (.I0(n356[6]), .I1(n382[6]), .I2(GND_net), 
            .I3(GND_net), .O(n71289));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i13_rep_180_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52902_4_lut (.I0(n356[7]), .I1(n71289), .I2(n382[7]), .I3(n67847), 
            .O(n69077));
    defparam i52902_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i17_rep_183_2_lut (.I0(n356[8]), .I1(n382[8]), .I2(GND_net), 
            .I3(GND_net), .O(n71292));   // verilog/motorControl.v(51[33:53])
    defparam LessThan_21_i17_rep_183_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52529_4_lut (.I0(n356[9]), .I1(n71292), .I2(n382[9]), .I3(n69077), 
            .O(n68704));
    defparam i52529_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i53257_4_lut (.I0(n356[11]), .I1(n71270), .I2(n382[11]), .I3(n68704), 
            .O(n69432));
    defparam i53257_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51655_4_lut (.I0(n356[13]), .I1(n71265), .I2(n382[13]), .I3(n69432), 
            .O(n67829));
    defparam i51655_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5099[3]), 
            .I3(n51540), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_5 (.CI(n51540), .I0(GND_net), .I1(n1_adj_5099[3]), 
            .CO(n51541));
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_5017));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5016));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_5015));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4988));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3844[0] ));   // verilog/motorControl.v(47[18] 49[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51619_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n356[3]), .I2(n356[2]), 
            .I3(PWMLimit[2]), .O(n67793));   // verilog/motorControl.v(52[14:29])
    defparam i51619_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4987));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_23_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n356[3]), 
            .I2(n356[2]), .I3(GND_net), .O(n6_adj_5090));   // verilog/motorControl.v(52[14:29])
    defparam LessThan_23_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4986));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4985));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4984));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4983));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4982));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6034_2_lut_4_lut (.I0(control_update), .I1(n69697), .I2(PWMLimit[23]), 
            .I3(n356[23]), .O(n12028));
    defparam i6034_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 i51557_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n356[21]), .I2(PWMLimit[9]), 
            .I3(n356[9]), .O(n67731));
    defparam i51557_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4975));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51570_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n356[16]), .I2(PWMLimit[7]), 
            .I3(n356[7]), .O(n67744));
    defparam i51570_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4963));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4962));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4958));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4955));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_5056));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4940));   // verilog/motorControl.v(50[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36883_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_5097), 
            .I3(n20598[1]), .O(n6_adj_4878));   // verilog/motorControl.v(50[18:24])
    defparam i36883_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_963 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n20598[1]), 
            .I3(n4_adj_5097), .O(n20538[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_963.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_964 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n20598[0]), 
            .I3(n51141), .O(n20538[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_964.LUT_INIT = 16'h8778;
    SB_LUT4 i36875_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n51141), 
            .I3(n20598[0]), .O(n4_adj_5097));   // verilog/motorControl.v(50[18:24])
    defparam i36875_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i36862_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n20538[0]));   // verilog/motorControl.v(50[18:24])
    defparam i36862_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36864_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n51141));   // verilog/motorControl.v(50[18:24])
    defparam i36864_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut_4_lut_adj_965 (.I0(\Kp[3] ), .I1(n1[19]), .I2(n20638[1]), 
            .I3(n4_adj_5098), .O(n20598[2]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_965.LUT_INIT = 16'h8778;
    SB_LUT4 i36788_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[19]), .I2(n4_adj_5098), 
            .I3(n20638[1]), .O(n6_adj_4886));   // verilog/motorControl.v(50[18:24])
    defparam i36788_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i36742_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n51002), 
            .I3(n20662[0]), .O(n4_adj_4887));   // verilog/motorControl.v(50[18:24])
    defparam i36742_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_966 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n20662[0]), 
            .I3(n51002), .O(n20638[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_966.LUT_INIT = 16'h8778;
    SB_LUT4 i36729_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n20638[0]));   // verilog/motorControl.v(50[18:24])
    defparam i36729_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36731_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n51002));   // verilog/motorControl.v(50[18:24])
    defparam i36731_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_5054));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36767_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n20598[0]));   // verilog/motorControl.v(50[18:24])
    defparam i36767_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_5053));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_5052));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_5051));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_5050));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_5049));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36780_3_lut_4_lut (.I0(n62_adj_4883), .I1(n131_adj_4882), .I2(n204_adj_4881), 
            .I3(n20638[0]), .O(n4_adj_5098));   // verilog/motorControl.v(50[18:24])
    defparam i36780_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut_adj_967 (.I0(n62_adj_4883), .I1(n131_adj_4882), 
            .I2(n204_adj_4881), .I3(n20638[0]), .O(n20598[1]));   // verilog/motorControl.v(50[18:24])
    defparam i1_3_lut_4_lut_adj_967.LUT_INIT = 16'h8778;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_5048));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_5047));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51859_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n68033));
    defparam i51859_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51058_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n67232));
    defparam i51058_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51502_2_lut_4_lut (.I0(n356[21]), .I1(n436[21]), .I2(n356[9]), 
            .I3(n436[9]), .O(n67676));
    defparam i51502_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51522_2_lut_4_lut (.I0(n356[16]), .I1(n436[16]), .I2(n356[7]), 
            .I3(n436[7]), .O(n67696));
    defparam i51522_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51269_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n67443));
    defparam i51269_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51325_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n67499));
    defparam i51325_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_5038));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3844[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5037));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_5035));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_5034));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_5033));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5032));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51703_2_lut_4_lut (.I0(deadband[17]), .I1(n356[17]), .I2(deadband[8]), 
            .I3(n356[8]), .O(n67877));
    defparam i51703_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51839_2_lut_4_lut (.I0(deadband[9]), .I1(n356[9]), .I2(deadband[5]), 
            .I3(n356[5]), .O(n68013));
    defparam i51839_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5031));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_5030));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_5029));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_5028));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5027));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5026));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_5025));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3844[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_5024));   // verilog/motorControl.v(50[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (GND_net, n3358, pwm_out, clk32MHz, VCC_net, reset, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n3358;
    output pwm_out;
    input clk32MHz;
    input VCC_net;
    input reset;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire n52653;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n52654, n58008, n52652, n48, n58046, n52651, n58080, 
        n52650, n58118, n52649, n58152, n52648, n58240, n52647, 
        n58342, n52646, n58476, n52645, n58574, n52644, n58576, 
        n52643, pwm_out_N_706, n58578, n52642, n58572, n57700, n57720, 
        n57740, n57760, n57782, n57806, n57832, n57854, n57884, 
        n57908, n57944, n57974, n39, n41, n45, n43, n29, n31, 
        n37, n23, n25, n35, n11, n13, n15, n27, n33, n9, 
        n17, n19, n21, n67684, n67670, n12, n30, n67705, n68582, 
        n68574, n69609, n69005, n69738, n6, n69342, n69343, n16, 
        n24, n67619, n8, n67596, n69157, n68156, n4, n69338, 
        n69339, n67657, n10, n67655, n69579, n68158, n69803, n69804, 
        n69802, n67632, n69476, n68164, n69685, n60972, n18, n21_adj_4557, 
        n20, n24_adj_4558, n19_adj_4559, n52664, n52663, n52662, 
        n52661, n52660, n52659, n52658, n52657, n52656, n52655;
    
    SB_CARRY pwm_counter_2049_add_4_14 (.CI(n52653), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n52654));
    SB_LUT4 pwm_counter_2049_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n52652), .O(n58008)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_13 (.CI(n52652), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n52653));
    SB_LUT4 pwm_counter_2049_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n52651), .O(n58046)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_12 (.CI(n52651), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n52652));
    SB_LUT4 pwm_counter_2049_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n52650), .O(n58080)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_11 (.CI(n52650), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n52651));
    SB_LUT4 pwm_counter_2049_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n52649), .O(n58118)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_10 (.CI(n52649), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n52650));
    SB_LUT4 pwm_counter_2049_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n52648), .O(n58152)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_9 (.CI(n52648), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n52649));
    SB_LUT4 pwm_counter_2049_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n52647), .O(n58240)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_8 (.CI(n52647), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n52648));
    SB_LUT4 pwm_counter_2049_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n52646), .O(n58342)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_7 (.CI(n52646), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n52647));
    SB_LUT4 pwm_counter_2049_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n52645), .O(n58476)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_6 (.CI(n52645), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n52646));
    SB_LUT4 pwm_counter_2049_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n52644), .O(n58574)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_5 (.CI(n52644), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n52645));
    SB_LUT4 pwm_counter_2049_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n52643), .O(n58576)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_4 (.CI(n52643), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n52644));
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n3358), .D(pwm_out_N_706));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_2049_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n52642), .O(n58578)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_3 (.CI(n52642), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n52643));
    SB_LUT4 pwm_counter_2049_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n58572)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n52642));
    SB_DFFR pwm_counter_2049__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n58572), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n57700), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n57720), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n57740), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n57760), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n57782), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n57806), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n57832), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n57854), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n57884), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n57908), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n57944), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n57974), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n58008), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n58046), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n58080), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n58118), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n58152), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n58240), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n58342), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n58476), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n58574), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n58576), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2049__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n58578), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51510_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n67684));
    defparam i51510_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51496_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n67670));
    defparam i51496_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52408_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n67705), 
            .O(n68582));
    defparam i52408_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52400_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n68582), 
            .O(n68574));
    defparam i52400_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53434_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n68574), 
            .O(n69609));
    defparam i53434_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52830_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n69609), 
            .O(n69005));
    defparam i52830_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53563_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69005), 
            .O(n69738));
    defparam i53563_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53167_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n69342));   // verilog/pwm.v(21[8:24])
    defparam i53167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53168_3_lut (.I0(n69342), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n69343));   // verilog/pwm.v(21[8:24])
    defparam i53168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51445_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n67684), 
            .O(n67619));
    defparam i51445_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52982_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n67596), 
            .O(n69157));   // verilog/pwm.v(21[8:24])
    defparam i52982_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51982_3_lut (.I0(n69343), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n68156));   // verilog/pwm.v(21[8:24])
    defparam i51982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53163_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n69338));   // verilog/pwm.v(21[8:24])
    defparam i53163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53164_3_lut (.I0(n69338), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n69339));   // verilog/pwm.v(21[8:24])
    defparam i53164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51483_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n67670), 
            .O(n67657));
    defparam i51483_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53404_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n67655), 
            .O(n69579));   // verilog/pwm.v(21[8:24])
    defparam i53404_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51984_3_lut (.I0(n69339), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n68158));   // verilog/pwm.v(21[8:24])
    defparam i51984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53628_4_lut (.I0(n68158), .I1(n69579), .I2(n35), .I3(n67657), 
            .O(n69803));   // verilog/pwm.v(21[8:24])
    defparam i53628_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53629_3_lut (.I0(n69803), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n69804));   // verilog/pwm.v(21[8:24])
    defparam i53629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53627_3_lut (.I0(n69804), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n69802));   // verilog/pwm.v(21[8:24])
    defparam i53627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51458_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n69738), 
            .O(n67632));
    defparam i51458_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53301_4_lut (.I0(n68156), .I1(n69157), .I2(n45), .I3(n67619), 
            .O(n69476));   // verilog/pwm.v(21[8:24])
    defparam i53301_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51990_3_lut (.I0(n69802), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n68164));   // verilog/pwm.v(21[8:24])
    defparam i51990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53510_4_lut (.I0(n68164), .I1(n69476), .I2(n45), .I3(n67632), 
            .O(n69685));   // verilog/pwm.v(21[8:24])
    defparam i53510_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53511_3_lut (.I0(n69685), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_706));   // verilog/pwm.v(21[8:24])
    defparam i53511_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n60972));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[17]), .I1(n60972), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i5_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[15]), .I2(pwm_counter[18]), 
            .I3(pwm_counter[16]), .O(n21_adj_4557));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n21_adj_4557), .I1(pwm_counter[19]), .I2(n18), 
            .I3(pwm_counter[14]), .O(n24_adj_4558));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[13]), .I1(pwm_counter[12]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4559));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4559), .I2(n24_adj_4558), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_counter_2049_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n52664), .O(n57700)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2049_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n52663), .O(n57720)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_24 (.CI(n52663), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n52664));
    SB_LUT4 pwm_counter_2049_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n52662), .O(n57740)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_23 (.CI(n52662), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n52663));
    SB_LUT4 pwm_counter_2049_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n52661), .O(n57760)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_22 (.CI(n52661), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n52662));
    SB_LUT4 pwm_counter_2049_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n52660), .O(n57782)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_21 (.CI(n52660), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n52661));
    SB_LUT4 pwm_counter_2049_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n52659), .O(n57806)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_20 (.CI(n52659), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n52660));
    SB_LUT4 pwm_counter_2049_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n52658), .O(n57832)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_19 (.CI(n52658), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n52659));
    SB_LUT4 pwm_counter_2049_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n52657), .O(n57854)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_18 (.CI(n52657), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n52658));
    SB_LUT4 pwm_counter_2049_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n52656), .O(n57884)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_17 (.CI(n52656), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n52657));
    SB_LUT4 pwm_counter_2049_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n52655), .O(n57908)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_16 (.CI(n52655), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n52656));
    SB_LUT4 pwm_counter_2049_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n52654), .O(n57944)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2049_add_4_15 (.CI(n52654), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n52655));
    SB_LUT4 pwm_counter_2049_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n52653), .O(n57974)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2049_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51531_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n67705));   // verilog/pwm.v(21[8:24])
    defparam i51531_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51422_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n67596));
    defparam i51422_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51481_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n67655));
    defparam i51481_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
