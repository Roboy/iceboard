// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Oct 30 19:28:15 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    inout PIN_9 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    inout PIN_10 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    inout PIN_11 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_1, PIN_7_c_0, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(67[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(68[12:17])
    
    wire blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(151[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(152[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(189[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(190[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(191[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(192[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(193[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(194[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(196[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(197[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(198[22:35])
    
    wire n41317;
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(200[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(225[22:33])
    
    wire n5961, n5960, n5957, n5956, n5923;
    wire [7:0]color_23__N_164;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n1172, n1166, n1258, n1257, n1256, n1255, n1254, n8, 
        blink_N_255, n1253, n43329;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105, n40668, n40660, n40654, n1252;
    wire [31:0]motor_state_23__N_106;
    wire [24:0]displacement_23__N_229;
    wire [23:0]displacement_23__N_80;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n42390, n6045, n6044, n6043, n6042, n6041, n6040, n6039, 
        n6038, n6037, n6036, n6035, n6067, n6066, n6065, n6064, 
        n6063, n6062, n6061, n6060, n6059, n6058, n6057, n6056, 
        n1251, n1250, n42285, n6055, n6054, n6081, n6080, n6079, 
        n6078, n6074, n42281;
    wire [3:0]state_3__N_362;
    
    wire n42280, n28325;
    wire [31:0]one_wire_N_513;
    
    wire n42276, n28324, n3008, n3007, n3006, n4442, n35679, n2825, 
        n2823, n2821, n2819, n2817, n3015_adj_4671, n99, n98, 
        n97, n89, n1184, n3005, n3004, n15, n17111, n57, n55, 
        n68, n60, n61, n56, n3003, n3002, n4648, n15_adj_4672, 
        n4670, n15_adj_4673, n3001, n3000, n2999, n58, n2998, 
        n2997, n2996, n2995, n2968, n42268, n63, n94, n93, n92, 
        n91, n2967, n2966, n2965, n2964, n2963, n2962, n2961, 
        n2960, n2959, n2958, n2957, n2956, n2955, n2954, n2953, 
        n2952, n2951, n2950, n2949, n2948, n2947, n2946, n2945, 
        n90, n87, n42263, n672, n671, n670, n669, n668, n667, 
        n666, n665, n664, n663, n662, n661, n660, n659, n658, 
        n657, n656, n655, n654, n653, n652, n651, n650, n649, 
        n648, n1158, n33461, n88, n86, n96, n1157;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n28125, n5970, n5994, n5993, n5992, n5991, n5990, n5988, 
        n28323, n10, n81, n72, n1156, n5987, n5986, n5985, n6007, 
        n6006, n6005, n6004, n6003, n6002, n6001, n3, n4, n5, 
        n6, n7, n8_adj_4674, n9, n10_adj_4675, n11, n12, n13, 
        n14, n15_adj_4676, n16, n17, n18, n19, n20, n21, n22, 
        n23, n24, n25, n1155, n1154, n1153, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n28322, n28321;
    wire [7:0]\data_in_frame[24] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n1152, n1151, n2, n28124, n122;
    wire [31:0]\FRAME_MATCHER.state_31__N_2661 ;
    
    wire n28123, n28320, n28122, n28319, n28121, n5927, n5926, 
        n28318, n28317, n28316, n28315, n42214, n42213, n41307, 
        n28120, n28119, n42210, n42208, n28118, n28314, n28313, 
        n28117, n28116, n28115, n28312, n28311, n95, n28114, n28310, 
        n42205, n28113, n28112, n28309, n28308, n42201, n42267, 
        n788, n28307, n28306, n28305, n28304, n28111, n28110, 
        n28109, n28303, n28302, n4_adj_4677, n28301, n28108, n28107, 
        n28300, n42186, n28106, n28105, n28299, n28104, n42182, 
        n28298, n28297, n28296, n28103, n28295, n28294, n28293, 
        n42275, n5925, n15851, n42176, n42174, n42172, n28292, 
        n42170, n42168, n28291, n42167, n15883, n28290, n28102, 
        n28101, n28100, n28099, n28098, n28289, n42320, n28097, 
        n28096, n28095, n28288, n28094, n42398, n35625, n28287, 
        n28286, n42148, n28285, n28284, n28283, n15871, n28282, 
        n28281, n28280, n35687, n28279, n28278, n28277, n28276, 
        n28275, n28274, n28273, n35635, n35590, n28272, n27847, 
        n28271, n28270, n28269, n28268, n27846, n28267, n28266, 
        n28265, n28264, n15866, n42283, n28263, n15863, n42143, 
        n28262, n42141, n15860, n27845, n28261, n15857, n43694, 
        n2957_adj_4678, n15854, n6_adj_4679, n22_adj_4680, n28260, 
        n19_adj_4681, n18_adj_4682, n16_adj_4683, n1319, n1320, n3894, 
        n35671, n40596, n41289, n41573, n15845, n28259, n28258, 
        n28257, n41283, n42101, n42099, n35523, n35521, n28256, 
        n28060, n41833, n41575, n42095, n42215, n41272, n15880, 
        n42217, n42219, n28255, n15817, n42075, n27844, n28059, 
        n15812, n42073, n28058, n27843, n15808, n42069, n42067, 
        n28057, n42065, n41264, n41262, n41663, n42064, n15804, 
        n15801, n41029, n28254, n28056, n28253, n28252, n28055, 
        n28251, n28250, n41974, n28054, n28053, n5921, n28249, 
        n1321, n1322, \FRAME_MATCHER.i_31__N_2621 , \FRAME_MATCHER.i_31__N_2625 , 
        n17743, n17742, n17741, n17740, n17739, n17738, n17737, 
        n17736, n17735, n17734, n17733, n17732, n17731, n17730, 
        n17729, n17728, n17727, n17726, n17725, n17724, n17723, 
        n17722, n17721, n17720, n17719, n17718, n17717, n17716, 
        n17714, n17713, n17712, n17711, n17710, n17709, n17708, 
        n17707, n17706, n17705, n17704, n17703, n17702, n17701, 
        n17700, n17699, n17698, n17697, n17696, n17695, n17694, 
        n17693, n17692, n17691, n17690, n17689, n17688, n17687, 
        n17686, n17685, n17684, n17683, n17682, n17681, n17680, 
        n17679, n17678, n17677, n17676, n17675, n17674, n17673, 
        n17672, n17671, n17670, n17669, n17668, n17667, n17666, 
        n17665, n17664, n17663, n17662, n17661, n17660, n17659, 
        n17658, n17657, n17656, n17655, n17654, n17653, n17652, 
        n17651, n17650, n17649, n17648, n17647, n17646, n17645, 
        n17644, n17643, n17642, n17641, n17640, n17639, n17638, 
        n17637, n17636, n17635, n17634, n17633, n17632, n17631, 
        n17630, n17629, n17628, n17627, n17626, n17625, n17624, 
        n17623, n17622, n17621, n17620, n17619, n17618, n17617, 
        n17616, n17615, n17614, n17613, n17612, n17611, n17610, 
        n17609, n17608, n17607, n17606, n17605, n17604, n17603, 
        n17602, n17601, n17600, n17599, n17598, n17597, n17596, 
        n17595, n17594, n17593, n17592, n17591, n17590, n17589, 
        n17588, n17587, n17586, n17585, n17584, n17583, n17582, 
        n17581, n17580, n17579, n17578, n17577, n17576, n17575, 
        n17574, n17573, n17572, n17571, n17570, n17569, n17568, 
        n17567, n17566, n17565, n17564, n17563, n17562, n17561, 
        n17560, n17559, n17558, n17557, n17555, n17554, n17553, 
        n17552, n17551, n17550, n17549, n17548, n17547, n17546, 
        n17545, n17544, n17543, n17542, n17541, n17540, n17539, 
        n17538, n17537, n17536, n17535, n17534, n17533, n17532, 
        n17531, n17530, n17529, n17528, n17527, n17526, n17525, 
        n42030, n558, n534, n533, n41254, n41252, n511, n510, 
        n1125, n1124, n1123, n1122, n1121, n1120, n1425, n1424, 
        n1423, n1422, n1421, n1420, n1419, n1418, n1417, n1085, 
        n28248, n41962, n393, n392, n1354, n1351, n17523, n1349, 
        n1353, n1352, n1358, n1357, n1356, n1355, n369, n17522, 
        n17521, n17520, n17519, n17518, n17517, n17516, n17515, 
        n17514, n17513, n17512, n17511, n17510, n17509, n17508, 
        n17507, n17506, n17505, n17504, n17503, n17502, n17501, 
        n28247, n28246, n17493, n17492, n17491, n28245, n28244, 
        n1058, n1057, n1056, n1055, n1054, n41958, n1053, n1052, 
        n41242, n5920, n1025, n1024, n1023, n1022, n1021, n5952, 
        n5951, n5949, n5948, n5947, n5946, n5945, n5944, n5943, 
        n5942, n5966, n5965, n71, n28243, n73, n83, n84, n28052, 
        n41951, n28051, n28242, n41839, n28241, n28240, n28239, 
        n28238, n28237, n28236, n28235, n28234, n28233, n28050, 
        n28049, n28048, n28047, n28046, n28045, n28232, n28044, 
        n41937, n41240, n20_adj_4684, n18_adj_4685, n41236, n16_adj_4686, 
        n17490, n28043, n35653, n28042, n6076, n6077, n28041, 
        n28231, n41232, n28230, n28229, n80, n82, n28040, n5924, 
        n1350, n15797, n17489, n28228, n28039, n8_adj_4687, n28227, 
        n41928, n6_adj_4688, n42068, n28226, n4372, n4371, n4370, 
        n4369, n4368, n4367, n4366, n4365, n4364, n4363, n4362, 
        n4361, n4360, n4359, n4358, n4357, n4356, n4355, n4354, 
        n4353, n28225, n28224, n4_adj_4689, n4352, n4351, n4350, 
        n4349, n63_adj_4690, n59, n44, n43, n42, n41, n40, n38, 
        n8_adj_4691, n17488, n17487, n17486, n17485, n17484, n17483, 
        n17482, n17481, n17480, n17479, n17478, n17477, n62, quadA_debounced, 
        quadB_debounced, count_enable, n11_adj_4692, n28223, n7_adj_4693, 
        n10_adj_4694, n39, n9_adj_4695, n37, n36, n8_adj_4696, n7_adj_4697, 
        n5964, n5963, n5962, n5959, n5958, n34, n33, n28222, 
        n6_adj_4698, quadA_debounced_adj_4699, quadB_debounced_adj_4700, 
        count_enable_adj_4701, n15794, n17476, n17475, n17474, n17473, 
        n17472, n17471, n17470, n75, n17469, n3_adj_4702, n28221, 
        n53, n3018, n3017, n3016, n3015, n3014, n3013, n3012, 
        n3011, n3010, n3009, n249, n248, n27, n64, n85, n22_adj_4703, 
        n4_adj_4704, n17468, n79, n78, n17467, n17466, n17465, 
        n17464, n17463, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n66, n69, n17462, n33441, n33443, n17452, n34135, n5919, 
        n5933, n5932, n5931, n28220, n17446, n28219, n1325, n1324, 
        n1323, n224, n33445, n17431, n17429, n35692, n3_adj_4705, 
        n17428;
    wire [2:0]r_SM_Main_adj_5379;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5381;   // verilog/uart_tx.v(33[16:27])
    
    wire n28218;
    wire [2:0]r_SM_Main_2__N_3579;
    
    wire n28217, n17427, n17426, n17425, n17424, n33453, n33455, 
        n28992, n28991, n28990, n28989, n28988, n17417, n33457, 
        n17413, n17412, n17411, n17410, n33459, n28987, n28216, 
        n28986, n28985, n28984, n28983;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n33463, n28982, n17403, n28981, n54;
    wire [1:0]reg_B_adj_5390;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17402, n17401, n28980, n17399, n17398, n28979, n28978, 
        n15791, n17396, n28977, n17395, n17394, n17393, n17392, 
        n33465, n28976, n74, n5971, n28975, n28974, n28973, n33467, 
        n28972, n28971, n28970, n4_adj_4713, n28215, n5969, n28969, 
        n28968, n28967, n28966, n33469, n28965, n28964, n33471, 
        n15_adj_4714, n28963, n28962, n6_adj_4715, n5_adj_4716, n4_adj_4717, 
        n28961, n28960, n28959, n28958, n28957, n29, n28956, n28955, 
        n28954, n33473, n33475, n28953, n28952, n28951, n9_adj_4718, 
        n28950, n8_adj_4719, n28949, n7_adj_4720, n41218, n28948, 
        n28947, n28946, n33477, n28945, n5997, n41216, n15_adj_4721, 
        n14_adj_4722, n13_adj_4723, n28944, n28943, n28942, n12_adj_4724, 
        n28941, n11_adj_4725, n28940, n28939, n28938, n28937, n28936, 
        n28935, n33483, n70, n5996, n28934, n1382, n17_adj_4726, 
        n28933, n16_adj_4727, n28932, n28931, n28930, n28929, n28928, 
        n41214, n33485, n77, n28927, n28926, n24_adj_4728, n23_adj_4729, 
        n22_adj_4730, n21_adj_4731, n20_adj_4732, n19_adj_4733, n18_adj_4734, 
        n28925, n28924, n28923, n33487, n33489, n65, n28922, n15626, 
        n28921, n28920, n28919, n1283, n6075, n33491, n67, n28918, 
        n28917, n28916, n28915, n28914, n28913, n28912, n28911, 
        n28910, n28909, n25_adj_4735, n28908, n15788, n28907, n28906, 
        n28905, n28904, n28903, n28902, n28901, n28900, n28899, 
        n28898, n28897, n5995, n33493, n33495, n28896, n28895, 
        n28894, n28893, n28892, n28891, n28890, n28889, n28888, 
        n5989, n1318, n28887, n28886, n5984, n4_adj_4736, n28885, 
        n28884, n33497, n28883, n28882, n28881, n28880, n28879, 
        n28878, n28877, n33499, n17343, n17342, n28876, n17341, 
        n28875, n17338, n28874, n34179, n28873, n12_adj_4737, n13_adj_4738, 
        n14_adj_4739, n15_adj_4740, n16_adj_4741, n17_adj_4742, n18_adj_4743, 
        n19_adj_4744, n20_adj_4745, n21_adj_4746, n22_adj_4747, n23_adj_4748, 
        n24_adj_4749, n25_adj_4750, n986, n28872, n13263, n958, 
        n957, n956, n955, n954, n953, n783, n784, n785, n41589, 
        n806, n807, n35588, n914, n915, n916, n917, n918, n938, 
        n939, n884, n1043, n1044, n1045, n1046, n1047, n1048, 
        n1067, n1068, n41591, n41868, n5912, n5913, n5914, n5915, 
        n5916, n28871, n855, n28870, n852, n28869, n1169, n1170, 
        n1171, n1172_adj_4751, n1173, n1174, n1175, n41864, n1193, 
        n1194, n28868, n28867, n1292, n1293, n1294, n1295, n1296, 
        n1297, n1298, n1299, n41861, n1316, n1317, n41862, n42307, 
        n5934, n5935, n5936, n5937, n5938, n5939, n1412, n1413, 
        n1414, n1415, n1416, n1417_adj_4752, n1418_adj_4753, n1419_adj_4754, 
        n1420_adj_4755, n1436, n1437, n40564, n28866, n28865, n749, 
        n748, n746, n1529, n1530, n1531, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1553, n1554, n28864, n28863, 
        n28862, n28861, n28860, n28859, n28858, n28857, n28856, 
        n28855, n41856, n1643, n1644, n1645, n1646, n1647, n1648, 
        n1649, n1650, n1651, n1652, n1653, n28854, n1667, n1668, 
        n28853, n28852, n26, n24_adj_4756, n22_adj_4757, n43090, 
        n43093, n43096, n43099, n28851, n5972, n5973, n5974, n5975, 
        n5976, n5977, n5978, n5979, n5980, n5981, n28850, n3453, 
        n3454, n3455, n3456, n3457, n3458, n43102, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n3452, n28849, n28848, n1778, n1779, n28847, 
        n41847, n35527, n35529, n28846, n28845, n28844, n28843, 
        n28842, n28841, n28840, n28839, n28838, n28837, n28836, 
        n28835, n28834, n28833, n28832, n28831, n18067, n1862, 
        n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
        n1871, n1872, n1873, n1874, n18066, n18064, n18063, n18062, 
        n1886, n1887, n18061, n18060, n18059, n18058, n18057, 
        n18056, n18055, n18054, n18053, n18052, n18051, n18050, 
        n18049, n18048, n18047, n6008, n6009, n6010, n6011, n6012, 
        n6013, n6014, n6032, n18046, n18045, n18044, n18043, n28830, 
        n28829, n1967, n1968, n1969, n1970, n1971, n1972, n1973, 
        n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1991, 
        n1992, n18042, n18041, n18040, n18039, n41855, n10627, 
        n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
        n6025, n6026, n6027, n6028, n6029, n6030, n6031, n3360, 
        n28828, n3362, n18038, n28827, n2069, n2070, n2071, n2072, 
        n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
        n2081, n2082, n2083, n3358, n3357, n3356, n3355, n3354, 
        n3353, n3352, n3351, n3350, n2093, n2094, n18036, n33435, 
        n3348, n3347, n3346, n3345, n3344, n3343, n3342, n3341, 
        n18031, n18030, n18029, n6046, n6047, n6048, n6049, n6050, 
        n6051, n18_adj_4758, n3334, n3335, n3336, n3337, n3338, 
        n3339, n3340, n33433, n16_adj_4759, n2168, n2169, n2170, 
        n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
        n2179, n2180, n2181, n2182, n2183, n3333, n3332, n3331, 
        n3330, n3329, n33431, n2192, n2193, n18022, n13_adj_4760, 
        n41852, n18_adj_4761, n18020, n28826, n6068, n6069, n6070, 
        n6071, n6186, n28825, n28824, n2264, n2265, n2266, n2267, 
        n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
        n2276, n2277, n2278, n2279, n2280, n2288, n2289, n28823, 
        n28822, n6082, n6083, n6084, n6085, n6086, n6087, n6088, 
        n6089, n6090, n6091, n6092, n18012, n6114, n6137, n18011, 
        n6161, n18010, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
        n2371, n2372, n2373, n2374, n18009, n18008, n2381, n2382, 
        n18007, n18006, n18005, n6095, n6096, n6097, n6098, n6099, 
        n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
        n6108, n6109, n6110, n6111, n6112, n6113, n2447, n2448, 
        n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
        n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
        n2465, n2471, n2472, n18004, n18003, n28821, n6117, n6118, 
        n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
        n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, 
        n6135, n6136, n18002, n3263, n41851, n18001, n18000, n2534, 
        n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
        n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
        n2551, n2552, n2553, n28820, n2558, n2559, n17999, n28214, 
        n28819, n3257, n3256, n3255, n17998, n6140, n6141, n6142, 
        n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, 
        n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, 
        n6159, n6160, n3253, n3254, n17997, n2618, n2619, n2620, 
        n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
        n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
        n2637, n2638, n3252, n3251, n3250, n2642, n2643, n17996, 
        n28818, n28817, n28816, n3248, n3247, n6164, n6165, n6166, 
        n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
        n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, 
        n6183, n6184, n6185, n3246, n2699, n2700, n2701, n2702, 
        n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
        n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
        n2719, n2720, n3245, n3244, n2723, n2724, n17995, n3243, 
        n41671, n3242, n2777, n2798, n2799, n3241, n2801, n2802, 
        n17994, n28815, n28814, n17993, n17992, n17991, n17990, 
        n17988, n17987, n17986, n17985, n17984, n17983, n17982, 
        n17981, n17980, n28213, n3239, n3238, n3237, n3236, n3235, 
        n3234, n3233, n3232, n3231, n3230, n3225, n3224, n3223, 
        n3222, n3221, n3220, n3219, n3218, n3217, n3216, n3215, 
        n42309, n17979, n17978, n17977, n28813, n28812, n3214, 
        n28811, n28810, n3213, n3212, n28809, n28808, n28807, 
        n3211, n3210, n28806, n3209, n3208, n3207, n3206, n28805, 
        n3205, n3204, n28804, n28803, n3203, n3202, n3201, n17976, 
        n17975, n17974, n17973, n17972, n17971, n17970, n17969, 
        n17968, n17967, n17966, n17965, n17964, n17963, n17962, 
        n17961, n17960, n17959, n17958, n17957, n17956, n17955, 
        n17954, n17953, n17952, n17951, n17950, n17949, n17948, 
        n17947, n3200, n3199, n17946, n28802, n17945, n17944, 
        n17943, n28801, n17942, n17941, n17940, n17939, n17938, 
        n17937, n17936, n17935, n28800, n28799, n28798, n28797, 
        n28796, n28795, n3164, n28794, n3158, n3157, n3156, n3155, 
        n17058, n3154, n3153, n3152, n3151, n3150, n3149, n17052, 
        n3148, n3147, n3146, n3145, n3144, n3143, n3142, n3141, 
        n3140, n3139, n3138, n3137, n3136, n17314, n3135, n3134, 
        n17189, n3133, n3132, n3131, n3125, n3124, n3123, n3122, 
        n3121, n3120, n3119, n3118, n3117, n3116, n3115, n3114, 
        n3113, n3112, n3111, n3110, n3109, n3108, n3107, n3106, 
        n3105, n17311, n3104, n15734, n17008, n3103, n3102, n3101, 
        n3100, n3065, n28793, n3058, n3057, n3056, n3055, n3054, 
        n3053, n3052, n3051, n3050, n3049, n3048, n3047, n28792, 
        n28212, n28791, n5922, n3046, n3045, n3044, n3043, n3042, 
        n3041, n3040, n3039, n3038, n3037, n3036, n3035, n3034, 
        n3033, n3032, n3025, n3024, n3023, n3022, n3021, n3020, 
        n3019, n3018_adj_4762, n3017_adj_4763, n41613, n28790, n40534, 
        n28789, n40531, n28788, n40529, n28787, n40527, n41887, 
        n41139, n41857, n28786, n28785, n28784, n28783, n41617, 
        n28782, n3016_adj_4764, n41135, n28781, n15778, n15774, 
        n15744, n33_adj_4765, n32, n31, n30, n29_adj_4766, n28, 
        n27_adj_4767, n26_adj_4768, n25_adj_4769, n24_adj_4770, n23_adj_4771, 
        n22_adj_4772, n21_adj_4773, n20_adj_4774, n19_adj_4775, n18_adj_4776, 
        n17_adj_4777, n16_adj_4778, n15_adj_4779, n14_adj_4780, n13_adj_4781, 
        n12_adj_4782, n3014_adj_4783, n3013_adj_4784, n3012_adj_4785, 
        n3011_adj_4786, n3010_adj_4787, n3009_adj_4788, n28780, n3008_adj_4789, 
        n3007_adj_4790, n28779, n28778, n3006_adj_4791, n28777, n3005_adj_4792, 
        n3004_adj_4793, n3003_adj_4794, n3002_adj_4795, n3001_adj_4796, 
        n26_adj_4797, n28776, n28775, n28774, n28773, n2966_adj_4798, 
        n36_adj_4799, n35, n28772, n34_adj_4800, n33_adj_4801, n2958_adj_4802, 
        n2957_adj_4803, n2956_adj_4804, n2955_adj_4805, n2954_adj_4806, 
        n2953_adj_4807, n2952_adj_4808, n2951_adj_4809, n2950_adj_4810, 
        n2949_adj_4811, n2948_adj_4812, n2947_adj_4813, n2946_adj_4814, 
        n2945_adj_4815, n2944, n2943, n2942, n31_adj_4816, n2941, 
        n2940, n2939, n2938, n2937, n2936, n28771, n2935, n2934, 
        n28770, n28769, n2933, n28768, n28767, n28766, n28765, 
        n28764, n28763, n28762, n2925, n2924, n2923, n2922, n2921, 
        n2920, n2919, n2918, n2917, n2916, n2915, n2914, n2913, 
        n24_adj_4817, n2912, n2911, n2910, n2909, n2908, n2907, 
        n2906, n2905, n2904, n2903, n2902, n28761, n28760, n28759, 
        n28758, n28757, n28756, n28755, n28754, n28753, n28752, 
        n2867, n28751, n2858, n2857, n2856, n2855, n2854, n2853, 
        n2852, n2851, n28750, n2850, n2849, n28749, n28748, n2848, 
        n28747, n2847, n2846, n2845, n2844, n2843, n2842, n2841, 
        n2840, n2839, n2838, n7_adj_4818, n2837, n2836, n2835, 
        n2834, n28746, n28745, n28744, n28743, n2824, n28742, 
        n2822, n28741, n2820, n28740, n2818, n2816, n2815, n2814, 
        n35595, n2813, n2812, n2811, n2810, n2809, n2808, n2807, 
        n2806, n2805, n2804, n2803, n34_adj_4819, n33_adj_4820, 
        n32_adj_4821, n2768, n28739, n28738, n31_adj_4822, n30_adj_4823, 
        n2758, n2757, n2756, n2755, n2754, n2753, n2752, n2751, 
        n2750, n2749, n2748, n2747, n2746, n11_adj_4824, n10_adj_4825, 
        n9_adj_4826, n8_adj_4827, n7_adj_4828, n6_adj_4829, n5_adj_4830, 
        n4_adj_4831, n3_adj_4832, n28737, n1778_adj_4833, n2743, n1844, 
        n1813, n1845, n1814, n1846, n1815, n1847, n1816, n1848, 
        n1817, n1849, n1818, n1850, n1819, n1851, n1820, n1852, 
        n1821, n1853, n1822, n1854, n1823, n1855, n1824, n1856, 
        n1825, n1857, n1858, n41123, n3240, n2744, n2745, n134, 
        n135, n136, n137, n138, n139, n140, n141, n142, n143, 
        n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, 
        n162, n163, n164, n165, n1745, n1746, n1747, n1748, 
        n1749, n1750, n1751, n1752, n1753, n1754_adj_4834, n1755_adj_4835, 
        n1756_adj_4836, n1757_adj_4837, n1758_adj_4838, n2742, n1714, 
        n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
        n1723, n1724, n1725, n2741, n2739, n2738, n2737, n2736, 
        n2735, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1646_adj_4839, n28736, n1647_adj_4840, 
        n1679, n1648_adj_4841, n1649_adj_4842, n28_adj_4843, n1650_adj_4844, 
        n1651_adj_4845, n1652_adj_4846, n1653_adj_4847, n1654, n1655, 
        n1656, n1657, n1658, n2740, n40516, n6_adj_4848, n36881, 
        n40489, n1615, n1553_adj_4849, n1554_adj_4850, n1555, n1556, 
        n1557, n1558, n41065, n28735, n1580, n1523, n1524, n1525, 
        n1547, n1548, n1549, n1550, n1551, n1552, n41893, n33479, 
        n33481, n17249, n17248, n28211, n28210, n28209, n28208, 
        n28734, n1481, n27_adj_4851, n5_adj_4852, n1225, n1224, 
        n1223, n1222, n1221, n1220, n1219, n1516, n1517, n1518, 
        n1519, n1520, n1521, n1522, n1453, n1454, n1455, n1456, 
        n1457, n1458, n28207, n28206, n28205, n1448, n1451, n1449, 
        n1452, n1450, n2669, n28733, n2658, n2657, n2656, n2655, 
        n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647, 
        n2646, n2645, n2644, n28732, n46, n2643_adj_4853, n2642_adj_4854, 
        n2641, n2640, n2639, n2638_adj_4855, n2637_adj_4856, n2636_adj_4857, 
        n16_adj_4858, n26_adj_4859, n2625_adj_4860, n2624_adj_4861, 
        n2623_adj_4862, n5950, n2622_adj_4863, n2621_adj_4864, n2620_adj_4865, 
        n2619_adj_4866, n2618_adj_4867, n2617, n2616, n2615, n2614, 
        n2613, n2612, n2611, n2610, n2609, n2608, n2607, n2606, 
        n2605, n11_adj_4868, n10_adj_4869, n28731, n2570, n28730, 
        n2558_adj_4870, n2557, n2556, n2555, n2554, n2553_adj_4871, 
        n2552_adj_4872, n2551_adj_4873, n2550_adj_4874, n2549_adj_4875, 
        n2548_adj_4876, n2547_adj_4877, n2546_adj_4878, n2545_adj_4879, 
        n2544_adj_4880, n2543_adj_4881, n2542_adj_4882, n2541_adj_4883, 
        n2540_adj_4884, n2539_adj_4885, n2538_adj_4886, n2537_adj_4887, 
        n25_adj_4888, n2525, n2524, n2523, n2522, n2521, n2520, 
        n2519, n2518, n2517, n2516, n2515, n2514, n2513, n2512, 
        n2511, n2510, n2509, n2508, n2507, n2506, n2_adj_4889, 
        n3_adj_4890, n4_adj_4891, n5_adj_4892, n6_adj_4893, n7_adj_4894, 
        n8_adj_4895, n9_adj_4896, n10_adj_4897, n11_adj_4898, n12_adj_4899, 
        n13_adj_4900, n14_adj_4901, n15_adj_4902, n16_adj_4903, n17_adj_4904, 
        n18_adj_4905, n19_adj_4906, n20_adj_4907, n21_adj_4908, n22_adj_4909, 
        n23_adj_4910, n24_adj_4911, n25_adj_4912, n2_adj_4913, n3_adj_4914, 
        n4_adj_4915, n5_adj_4916, n6_adj_4917, n7_adj_4918, n8_adj_4919, 
        n9_adj_4920, n10_adj_4921, n11_adj_4922, n12_adj_4923, n13_adj_4924, 
        n14_adj_4925, n15_adj_4926, n16_adj_4927, n17_adj_4928, n18_adj_4929, 
        n19_adj_4930, n20_adj_4931, n21_adj_4932, n22_adj_4933, n23_adj_4934, 
        n24_adj_4935, n25_adj_4936, n2471_adj_4937, n28729, n2458_adj_4938, 
        n2457_adj_4939, n2456_adj_4940, n2455_adj_4941, n2454_adj_4942, 
        n2453_adj_4943, n2452_adj_4944, n2451_adj_4945, n2450_adj_4946, 
        n2449_adj_4947, n2448_adj_4948, n2447_adj_4949, n2446, n2445, 
        n2444, n2443, n28728, n44_adj_4950, n2442, n2441, n2440, 
        n2439, n2438, n2425, n2424, n2423, n2422, n2421, n2420, 
        n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, 
        n2411, n2410, n2409, n2408, n2407, n41653, n28727, n42_adj_4951, 
        n42074, n2372_adj_4952, n28726, n41035, n2358_adj_4953, n2357_adj_4954, 
        n2356, n2355, n2354, n2353, n2352, n2351, n2350, n2349, 
        n2348, n2347, n2346, n2345, n2344, n2343, n2342, n2341, 
        n2340, n2339, n42282, n28725, n40_adj_4955, n42_adj_4956, 
        n44_adj_4957, n45, n2325, n2324, n2323, n2322, n2321, 
        n2320, n2319, n2318, n2317, n2316, n2315, n2314, n2313, 
        n2312, n2311, n2310, n2309, n2308, n28724, n38_adj_4958, 
        n40_adj_4959, n42_adj_4960, n43_adj_4961, n41661, n42072, 
        n2273_adj_4962, n28723, n28722, n28721, n2258, n2257, n2256, 
        n2255, n2254, n2253, n2252, n2251, n2250, n2249, n2248, 
        n2247, n2246, n2245, n2244, n2243, n2242, n2241, n2240, 
        n28720, n28719, n28718, n36_adj_4963, n38_adj_4964, n40_adj_4965, 
        n41_adj_4966, n42269, n2225, n2224, n2223, n2222, n2221, 
        n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, 
        n2212, n2211, n2210, n2209, n28717, n28716, n34_adj_4967, 
        n36_adj_4968, n38_adj_4969, n39_adj_4970, n41_adj_4971, n43_adj_4972, 
        n44_adj_4973, n45_adj_4974, n41665, n2174_adj_4975, n28715, 
        n41891, n2158, n2157, n2156, n2155, n2154, n2153, n2152, 
        n2151, n2150, n2149, n2148, n2147, n2146, n2145, n2144, 
        n2143, n28714, n32_adj_4976, n34_adj_4977, n37_adj_4978, n39_adj_4979, 
        n41_adj_4980, n42066, n43_adj_4981, n41931, n2142, n2141, 
        n28713, n28712, n2125, n2124, n2123, n2122, n2121, n2120, 
        n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, 
        n2111, n2110, n28711, n30_adj_4982, n31_adj_4983, n32_adj_4984, 
        n33_adj_4985, n34_adj_4986, n35_adj_4987, n37_adj_4988, n39_adj_4989, 
        n41_adj_4990, n42_adj_4991, n43_adj_4992, n45_adj_4993, n2075_adj_4994, 
        n28710, n28709, n28_adj_4995, n29_adj_4996, n30_adj_4997, 
        n31_adj_4998, n32_adj_4999, n33_adj_5000, n35_adj_5001, n37_adj_5002, 
        n39_adj_5003, n40_adj_5004, n41_adj_5005, n43_adj_5006, n42183, 
        n42354, n41013, n2058, n2057, n2056, n2055, n2054, n2053, 
        n2052, n2051, n2050, n2049, n2048, n2047, n2046, n2045, 
        n2044, n2043, n2042, n28708, n26_adj_5007, n27_adj_5008, 
        n28_adj_5009, n29_adj_5010, n30_adj_5011, n31_adj_5012, n33_adj_5013, 
        n35_adj_5014, n37_adj_5015, n38_adj_5016, n39_adj_5017, n41_adj_5018, 
        n42364, n2025, n2024, n2023, n2022, n2021, n2020, n2019, 
        n2018, n2017, n2016, n2015, n2014, n2013, n2012, n2011, 
        n28707, n40457, n24_adj_5019, n25_adj_5020, n26_adj_5021, 
        n27_adj_5022, n28_adj_5023, n29_adj_5024, n30_adj_5025, n31_adj_5026, 
        n32_adj_5027, n33_adj_5028, n35_adj_5029, n36_adj_5030, n37_adj_5031, 
        n39_adj_5032, n1976_adj_5033, n28706, n40455, n22_adj_5034, 
        n23_adj_5035, n24_adj_5036, n25_adj_5037, n26_adj_5038, n27_adj_5039, 
        n28_adj_5040, n29_adj_5041, n30_adj_5042, n31_adj_5043, n33_adj_5044, 
        n34_adj_5045, n35_adj_5046, n37_adj_5047, n39_adj_5048, n42207, 
        n41_adj_5049, n43_adj_5050, n41681, n42059, n42181, n28705, 
        n1958, n1957, n1956, n1955, n1954, n1953, n1952, n28704, 
        n20_adj_5051, n21_adj_5052, n22_adj_5053, n23_adj_5054, n24_adj_5055, 
        n25_adj_5056, n26_adj_5057, n27_adj_5058, n28_adj_5059, n29_adj_5060, 
        n31_adj_5061, n32_adj_5062, n33_adj_5063, n35_adj_5064, n37_adj_5065, 
        n42209, n39_adj_5066, n41_adj_5067, n41943, n42273, n1951, 
        n1950, n1949, n1948, n1947, n1946, n1945, n1944, n3349, 
        n1943, n28703, n40451, n18_adj_5068, n19_adj_5069, n20_adj_5070, 
        n21_adj_5071, n22_adj_5072, n23_adj_5073, n24_adj_5074, n25_adj_5075, 
        n26_adj_5076, n27_adj_5077, n29_adj_5078, n30_adj_5079, n31_adj_5080, 
        n33_adj_5081, n35_adj_5082, n37_adj_5083, n39_adj_5084, n41_adj_5085, 
        n43_adj_5086, n45_adj_5087, n41945, n1925, n1924, n1923, 
        n1922, n1921, n1920, n1919, n1918, n1917, n1916, n1915, 
        n1914, n1913, n28702, n16_adj_5088, n17_adj_5089, n18_adj_5090, 
        n19_adj_5091, n20_adj_5092, n21_adj_5093, n22_adj_5094, n23_adj_5095, 
        n25_adj_5096, n27_adj_5097, n28_adj_5098, n29_adj_5099, n31_adj_5100, 
        n33_adj_5101, n35_adj_5102, n37_adj_5103, n39_adj_5104, n41_adj_5105, 
        n41683, n43_adj_5106, n1912, n28701, n28700, n14_adj_5107, 
        n16_adj_5108, n17_adj_5109, n18_adj_5110, n19_adj_5111, n20_adj_5112, 
        n21_adj_5113, n22_adj_5114, n23_adj_5115, n25_adj_5116, n26_adj_5117, 
        n27_adj_5118, n29_adj_5119, n31_adj_5120, n33_adj_5121, n42144, 
        n35_adj_5122, n37_adj_5123, n42046, n39_adj_5124, n40_adj_5125, 
        n41_adj_5126, n43_adj_5127, n45_adj_5128, n42146, n28699, 
        n12_adj_5129, n14_adj_5130, n15_adj_5131, n16_adj_5132, n17_adj_5133, 
        n18_adj_5134, n19_adj_5135, n20_adj_5136, n21_adj_5137, n23_adj_5138, 
        n24_adj_5139, n25_adj_5140, n27_adj_5141, n29_adj_5142, n31_adj_5143, 
        n42284, n33_adj_5144, n35_adj_5145, n37_adj_5146, n38_adj_5147, 
        n39_adj_5148, n41_adj_5149, n41687, n43_adj_5150, n42033, 
        n1877, n28698, n28697, n10_adj_5151, n12_adj_5152, n13_adj_5153, 
        n14_adj_5154, n15_adj_5155, n16_adj_5156, n17_adj_5157, n18_adj_5158, 
        n19_adj_5159, n21_adj_5160, n22_adj_5161, n23_adj_5162, n25_adj_5163, 
        n27_adj_5164, n29_adj_5165, n30_adj_5166, n31_adj_5167, n33_adj_5168, 
        n34_adj_5169, n35_adj_5170, n36_adj_5171, n37_adj_5172, n39_adj_5173, 
        n41_adj_5174, n41867, n3258, n28696, n8_adj_5175, n10_adj_5176, 
        n11_adj_5177, n12_adj_5178, n13_adj_5179, n14_adj_5180, n15_adj_5181, 
        n16_adj_5182, n17_adj_5183, n19_adj_5184, n20_adj_5185, n21_adj_5186, 
        n23_adj_5187, n25_adj_5188, n41863, n27_adj_5189, n29_adj_5190, 
        n31_adj_5191, n33_adj_5192, n34_adj_5193, n35_adj_5194, n37_adj_5195, 
        n39_adj_5196, n41689, n42027, n3249, n28695, n6_adj_5197, 
        n8_adj_5198, n9_adj_5199, n10_adj_5200, n11_adj_5201, n12_adj_5202, 
        n13_adj_5203, n14_adj_5204, n15_adj_5205, n17_adj_5206, n19_adj_5207, 
        n21_adj_5208, n23_adj_5209, n41858, n25_adj_5210, n41691, 
        n27_adj_5211, n29_adj_5212, n31_adj_5213, n32_adj_5214, n33_adj_5215, 
        n35_adj_5216, n37_adj_5217, n28694, n4_adj_5218, n6_adj_5219, 
        n7_adj_5220, n8_adj_5221, n9_adj_5222, n10_adj_5223, n11_adj_5224, 
        n12_adj_5225, n13_adj_5226, n15_adj_5227, n16_adj_5228, n17_adj_5229, 
        n19_adj_5230, n21_adj_5231, n23_adj_5232, n24_adj_5233, n25_adj_5234, 
        n27_adj_5235, n42022, n29_adj_5236, n30_adj_5237, n31_adj_5238, 
        n33_adj_5239, n35_adj_5240, n37_adj_5241, n42155, n39_adj_5242, 
        n40_adj_5243, n41_adj_5244, n43_adj_5245, n45_adj_5246, n42157, 
        n34067, n28204, n5910, n5911, n5900, n5901, n5902, n5903, 
        n5904, n5905, n5906, n17180, n28693, n5893, n5894, n5895, 
        n5896, n5897, n28692, n28691, n40995, n28690, n28689, 
        n28688, n28687, n42_adj_5247, n41_adj_5248, n40_adj_5249, 
        n41983, n28686, n28685, n28684, n39_adj_5250, n28683, n6_adj_5251, 
        n28682, n35641, n28681, n28680, n28679, n37_adj_5252, n28678, 
        n36_adj_5253, n28677, n28203, n28202, n40965, n28676, n28675, 
        n28201, n40960, n24520, n28674, n40427, n28673, n40409, 
        n28672, n28671, n40401, n40397, n33451, n30_adj_5254, n19_adj_5255, 
        n40390, n40388, n33439, n28670, n35327, n11_adj_5256, n33429, 
        n28669, n28668, n28667, n40939, n42053, n5_adj_5257, n35548, 
        n28666, n41657, n40933, n28665, n40931, n28664, n28663, 
        n12_adj_5258, n28662, n28661, n28660, n28659, n28658, n43211, 
        n13_adj_5259, n42161, n28657, n28656, n40916, n28655, n28654, 
        n11_adj_5260, n28653, n28652, n28651, n30070, n28650, n28649, 
        n28648, n28647, n28646, n40374, n28645, n40900, n28644, 
        n28643, n28642, n28641, n28200, n28640, n28199, n28198, 
        n28639, n42287, n28638, n28637, n28636, n28635, n9001, 
        n28634, n28197, n40370, n40884, n28196, n28633, n28632, 
        n40881, n41523, n28631, n40879, n28630, n40876, n28629, 
        n28628, n28627, n41395, n28626, n28625, n28624, n10199, 
        n10198, n10197, n10196, n10195, n10194, n13_adj_5261, n11_adj_5262, 
        n24628, n28623, n28622, n28621, n28620, n28619, n28618, 
        n28617, n28616, n28615, n28614, n28613, n8936, n28612, 
        n28611, n35557, n28610, n28609, n28608, n28607, n28606, 
        n28605, n42366, n28604, n28603, n28190, n28602, n28601, 
        n28600, n28599, n40865, n40861, n28189, n40856, n28188, 
        n41503, n2_adj_5263, n40852, n40845, n35775, n40841, n42054, 
        n15785, n27890, n43086, n40802, n40798, n41991, n42316, 
        n42399, n40792, n3_adj_5264, n40351, n40786, n40784, n35658, 
        n27889, n42051, n40770, n28187, n40764, n27888, n35517, 
        n42368, n40754, n40748, n40746, n40743, n27887, n41995, 
        n40739, n38149, n40734, n27886, n42040, n28186, n40278, 
        n40277, n40276, n40275, n40274, n40273, n42039, n10_adj_5265, 
        n41892, n28185, n28534, n28533, n27885, n5892, n5909, 
        n42397, n5930, n34_adj_5266, n37976, n28532, n28531, n31_adj_5267, 
        n5955, n38143, n37972, n30_adj_5268, n28_adj_5269, n22_adj_5270, 
        n21_adj_5271, n6000, n28530, n40341, n40339, n40335, n40333, 
        n40258, n40330, n40629, n40256, n40316, n28529, n40644, 
        n40254, n40306, n40253, n40252, n40251, n40250, n40249, 
        n41997, n40248, n40247, n40246, n40245, n40244, n40243, 
        n40242, n40241, n40240, n40239, n40238, n40237, n40236, 
        n40235, n40234, n42296, n28528, n28527, n28526, n28525, 
        n28524, n28523, n40233, n40232, n28522, n40231, n28521, 
        n28520, n28519, n27884, n40230, n28518, n41757, n40229, 
        n40228, n28517, n28516, n28515, n28514, n40227, n40226, 
        n40225, n40224, n40223, n41888, n28513, n28512, n40218, 
        n28511, n40217, n35976, n41769, n42028, n28510, n28509, 
        n2_adj_5272, n3_adj_5273, n4_adj_5274, n5_adj_5275, n6_adj_5276, 
        n7_adj_5277, n8_adj_5278, n9_adj_5279, n10_adj_5280, n11_adj_5281, 
        n12_adj_5282, n13_adj_5283, n14_adj_5284, n15_adj_5285, n16_adj_5286, 
        n17_adj_5287, n18_adj_5288, n19_adj_5289, n20_adj_5290, n21_adj_5291, 
        n22_adj_5292, n23_adj_5293, n24_adj_5294, n25_adj_5295, n26_adj_5296, 
        n27_adj_5297, n28_adj_5298, n29_adj_5299, n30_adj_5300, n31_adj_5301, 
        n32_adj_5302, n33_adj_5303, n28508, n28507, n28506, n27883, 
        n28505, n28504, n28503, n28502, n28501, n35578, n28500, 
        n28499, n28498, n28497, n28496, n28495, n35565, n28494, 
        n28493, n28492, n28491, n35278, n28490, n28489, n27882, 
        n28488, n28487, n28486, n28485, n28484, n24450, n28483, 
        n28482, n28481, n28480, n28479, n28478, n28477, n27881, 
        n28476, n28475, n28474, n28473, n28472, n28471, n28470, 
        n29821, n6_adj_5304, n28469, n29820, n28468, n28467, n29819, 
        n29818, n29817, n28466, n29816, n28465, n28464, n29815, 
        n28463, n28462, n35573, n28461, n28460, n28459, n28458, 
        n29814, n29813, n29812, n28457, n28456, n28455, n29811, 
        n29810, n29809, n28454, n28453, n28452, n28451, n28450, 
        n29808, n29807, n28449, n28448, n28447, n28446, n28445, 
        n28444, n42025, n29806, n29805, n28443, n28442, n28441, 
        n28440, n29804, n28439, n29803, n42395, n37832, n28438, 
        n28437, n28436, n35620, n28435, n29802, n28434, n28433, 
        n28432, n35551, n28431, n29801, n29800, n29799, n35462, 
        n28430, n28429, n28428, n28427, n28426, n29798, n28425, 
        n28424, n28423, n28422, n28421, n28420, n28419, n28418, 
        n28417, n28416, n28415, n28414, n35424, n28413, n28412, 
        n28411, n29797, n35420, n28410, n28409, n29796, n28408, 
        n28407, n28406, n28405, n28404, n28403, n28402, n42304, 
        n28401, n28400, n42394, n28399, n28398, n28397, n23653, 
        n28396, n28395, n28394, n28393, n28392, n28391, n28390, 
        n28389, n28388, n29795, n28387, n28386, n29794, n29793, 
        n29792, n28385, n28384, n29791, n28383, n28382, n35299, 
        n35295, n28381, n28380, n28379, n28378, n40177, n28377, 
        n28376, n28141, n28140, n6_adj_5305, n4_adj_5306, n28139, 
        n28138, n37728, n28375, n28374, n2_adj_5307, n28137, n28136, 
        n2_adj_5308, n28373, n4_adj_5309, n28372, n28371, n28370, 
        n28369, n28368, n28367, n28366, n42013, n28365, n28364, 
        n28363, n28362, n28361, n28360, n35608, n28359, n28358, 
        n28357, n28356, n28355, n28354, n28353, n28352, n28351, 
        n28135, n28350, n28349, n28348, n37688, n28347, n37686, 
        n28346, n37684, n28345, n28344, n28343, n28342, n37678, 
        n28341, n28340, n28339, n28338, n28337, n28336, n28335, 
        n28334, n28333, n28332, n28331, n28330, n28329, n28328, 
        n28327, n28326, n24391, n37664, n37660, n41429, n41435, 
        n15_adj_5310, n14_adj_5311, n37614, n37612, n37610, n41884, 
        n43164, n34001, n40298, n37586, n34037, n40296, n43156, 
        n43152, n5_adj_5312, n37570, n37566, n36877, n40290, n43147, 
        n36115, n34173, n34177, n40285, n41883, n42303, n37474, 
        n41807, n30_adj_5313, n29_adj_5314, n28_adj_5315, n27_adj_5316, 
        n18_adj_5317, n41809, n42021, n42029, n40_adj_5318, n39_adj_5319, 
        n47, n38_adj_5320, n46_adj_5321, n37_adj_5322, n43_adj_5323, 
        n41_adj_5324, n40_adj_5325, n35_adj_5326, n34_adj_5327, n39_adj_5328, 
        n38_adj_5329, n34_adj_5330, n27_adj_5331, n34675, n28_adj_5332, 
        n26_adj_5333, n24_adj_5334, n19_adj_5335, n16_adj_5336, n42386, 
        n24_adj_5337, n22_adj_5338, n20_adj_5339, n42393, n42391, 
        n16_adj_5340, n42387, n42045, n42371, n42370, n42367, n42365, 
        n36887, n42355, n42353, n42345, n42344, n42335;
    
    VCC i2 (.Y(VCC_net));
    SB_IO ID1_input (.PACKAGE_PIN(PIN_10), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID1_input.PIN_TYPE = 6'b000001;
    defparam ID1_input.PULLUP = 1'b1;
    defparam ID1_input.NEG_TRIGGER = 1'b0;
    defparam ID1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO ID2_input (.PACKAGE_PIN(PIN_11), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID2_input.PIN_TYPE = 6'b000001;
    defparam ID2_input.PULLUP = 1'b1;
    defparam ID2_input.NEG_TRIGGER = 1'b0;
    defparam ID2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_CARRY div_46_unary_minus_2_add_3_13 (.CI(n28713), .I0(GND_net), .I1(n14_adj_4925), 
            .CO(n28714));
    SB_LUT4 i22_3_lut (.I0(bit_ctr[22]), .I1(n40243), .I2(n4442), .I3(GND_net), 
            .O(n33475));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_DFF h2_56 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_57 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF dir_61 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 i33511_4_lut (.I0(n35_adj_5145), .I1(n33_adj_5144), .I2(n31_adj_5143), 
            .I3(n41589), .O(n40341));
    defparam i33511_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i1194_3_lut_3_lut (.I0(n1778), .I1(n5976), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i12_4_lut (.I0(n666), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_5129));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35207_3_lut (.I0(n12_adj_5129), .I1(n87), .I2(n35_adj_5145), 
            .I3(GND_net), .O(n42039));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35207_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n28646), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_22 (.CI(n28646), .I0(n3039), .I1(VCC_net), 
            .CO(n28647));
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .bit_ctr({bit_ctr}), .VCC_net(VCC_net), 
            .n40238(n40238), .GND_net(GND_net), .n19(n19_adj_5255), .timer({timer}), 
            .n33435(n33435), .n33465(n33465), .n33467(n33467), .n33469(n33469), 
            .n33471(n33471), .n33473(n33473), .n33475(n33475), .n33477(n33477), 
            .n33429(n33429), .n33431(n33431), .n33443(n33443), .n33445(n33445), 
            .n33451(n33451), .n33453(n33453), .n33455(n33455), .n33457(n33457), 
            .n33497(n33497), .n33493(n33493), .n33495(n33495), .n33489(n33489), 
            .n33491(n33491), .n33485(n33485), .n33487(n33487), .n33479(n33479), 
            .n33481(n33481), .n33483(n33483), .n33463(n33463), .n33461(n33461), 
            .n33433(n33433), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n40237(n40237), .n40231(n40231), .\state_3__N_362[1] (state_3__N_362[1]), 
            .\state[1] (state[1]), .n1166(n1166), .\state[0] (state[0]), 
            .n4442(n4442), .n40236(n40236), .n40245(n40245), .n40234(n40234), 
            .n24628(n24628), .start(start), .n15744(n15744), .\one_wire_N_513[10] (one_wire_N_513[10]), 
            .\one_wire_N_513[8] (one_wire_N_513[8]), .\one_wire_N_513[5] (one_wire_N_513[5]), 
            .\one_wire_N_513[11] (one_wire_N_513[11]), .\one_wire_N_513[7] (one_wire_N_513[7]), 
            .\one_wire_N_513[9] (one_wire_N_513[9]), .\one_wire_N_513[6] (one_wire_N_513[6]), 
            .n35327(n35327), .n33459(n33459), .n33441(n33441), .n33439(n33439), 
            .n17493(n17493), .n17492(n17492), .n17491(n17491), .n17490(n17490), 
            .n17489(n17489), .n17488(n17488), .n17487(n17487), .n17486(n17486), 
            .n17485(n17485), .n17484(n17484), .n17483(n17483), .n17482(n17482), 
            .n17481(n17481), .n17480(n17480), .n17479(n17479), .n17478(n17478), 
            .n17477(n17477), .n17476(n17476), .n17475(n17475), .n17474(n17474), 
            .n17473(n17473), .n17472(n17472), .n17471(n17471), .n17470(n17470), 
            .n17469(n17469), .n17468(n17468), .n17467(n17467), .n17466(n17466), 
            .n17465(n17465), .n17464(n17464), .n17463(n17463), .n35462(n35462), 
            .n40230(n40230), .n35424(n35424), .n36115(n36115), .n17431(n17431), 
            .n40228(n40228), .n17008(n17008), .n35420(n35420), .PIN_8_c(PIN_8_c), 
            .n36877(n36877), .n40227(n40227), .n11(n11_adj_5256), .n40244(n40244), 
            .n33499(n33499), .n17248(n17248), .n40223(n40223), .n40235(n40235), 
            .n40224(n40224), .n40254(n40254), .n40253(n40253), .n40252(n40252), 
            .n40251(n40251), .n40226(n40226), .n40225(n40225), .n40250(n40250), 
            .n40249(n40249), .n40233(n40233), .n40248(n40248), .n40247(n40247), 
            .n40246(n40246), .n40243(n40243), .n40229(n40229), .n40232(n40232), 
            .n40242(n40242), .n40241(n40241), .n40240(n40240), .n40239(n40239), 
            .\color[2] (color[2]), .\color[3] (color[3]), .\color[4] (color[4]), 
            .\color[1] (color[1]), .n24520(n24520)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(98[10] 104[2])
    SB_IO ID0_input (.PACKAGE_PIN(PIN_9), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID0_input.PIN_TYPE = 6'b000001;
    defparam ID0_input.PULLUP = 1'b1;
    defparam ID0_input.NEG_TRIGGER = 1'b0;
    defparam ID0_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n28645), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4926), .I3(n28712), .O(n15_adj_4721)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_21 (.CI(n28645), .I0(n3040), .I1(VCC_net), 
            .CO(n28646));
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n28644), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_20 (.CI(n28644), .I0(n3041), .I1(VCC_net), 
            .CO(n28645));
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n28643), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_15 (.CI(n28910), .I0(n2046), .I1(VCC_net), 
            .CO(n28911));
    SB_CARRY rem_4_add_2055_19 (.CI(n28643), .I0(n3042), .I1(VCC_net), 
            .CO(n28644));
    SB_LUT4 div_46_LessThan_1606_i38_3_lut (.I0(n20_adj_5136), .I1(n83), 
            .I2(n43_adj_5150), .I3(GND_net), .O(n38_adj_5147));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35208_3_lut (.I0(n42039), .I1(n86), .I2(n37_adj_5146), .I3(GND_net), 
            .O(n42040));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35208_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_46_unary_minus_2_add_3_12 (.CI(n28712), .I0(GND_net), .I1(n15_adj_4926), 
            .CO(n28713));
    SB_LUT4 div_46_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4927), .I3(n28711), .O(n16_adj_4727)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_11 (.CI(n28711), .I0(GND_net), .I1(n16_adj_4927), 
            .CO(n28712));
    SB_LUT4 div_46_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4928), .I3(n28710), .O(n17_adj_4726)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n28909), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n28642), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_10 (.CI(n28710), .I0(GND_net), .I1(n17_adj_4928), 
            .CO(n28711));
    SB_CARRY rem_4_add_2055_18 (.CI(n28642), .I0(n3043), .I1(VCC_net), 
            .CO(n28643));
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n28641), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33505_4_lut (.I0(n41_adj_5149), .I1(n39_adj_5148), .I2(n37_adj_5146), 
            .I3(n40339), .O(n40335));
    defparam i33505_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35201_4_lut (.I0(n38_adj_5147), .I1(n18_adj_5134), .I2(n43_adj_5150), 
            .I3(n40333), .O(n42033));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35201_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_1385_14 (.CI(n28909), .I0(n2047), .I1(VCC_net), 
            .CO(n28910));
    SB_LUT4 i35130_3_lut (.I0(n42040), .I1(n85), .I2(n39_adj_5148), .I3(GND_net), 
            .O(n41962));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35130_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1199_3_lut_3_lut (.I0(n1778), .I1(n5981), .I2(n659), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n28908), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4929), .I3(n28709), .O(n18_adj_4734)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_13 (.CI(n28908), .I0(n2048), .I1(VCC_net), 
            .CO(n28909));
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n28907), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_9 (.CI(n28709), .I0(GND_net), .I1(n18_adj_4929), 
            .CO(n28710));
    SB_CARRY rem_4_add_2055_17 (.CI(n28641), .I0(n3044), .I1(VCC_net), 
            .CO(n28642));
    SB_LUT4 div_46_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4930), .I3(n28708), .O(n19_adj_4733)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_12 (.CI(n28907), .I0(n2049), .I1(VCC_net), 
            .CO(n28908));
    SB_CARRY div_46_unary_minus_2_add_3_8 (.CI(n28708), .I0(GND_net), .I1(n19_adj_4930), 
            .CO(n28709));
    SB_LUT4 div_46_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4931), .I3(n28707), .O(n20_adj_4732)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n28906), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_11 (.CI(n28906), .I0(n2050), .I1(VCC_net), 
            .CO(n28907));
    SB_CARRY div_46_unary_minus_2_add_3_7 (.CI(n28707), .I0(GND_net), .I1(n20_adj_4931), 
            .CO(n28708));
    SB_LUT4 div_46_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4932), .I3(n28706), .O(n21_adj_4731)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n28640), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_6 (.CI(n28706), .I0(GND_net), .I1(n21_adj_4932), 
            .CO(n28707));
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n28905), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4933), .I3(n28705), .O(n22_adj_4730)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_10 (.CI(n28905), .I0(n2051), .I1(VCC_net), 
            .CO(n28906));
    SB_CARRY div_46_unary_minus_2_add_3_5 (.CI(n28705), .I0(GND_net), .I1(n22_adj_4933), 
            .CO(n28706));
    SB_CARRY rem_4_add_2055_16 (.CI(n28640), .I0(n3045), .I1(VCC_net), 
            .CO(n28641));
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n28904), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4934), .I3(n28704), .O(n23_adj_4729)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n28639), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_15 (.CI(n28639), .I0(n3046), .I1(VCC_net), 
            .CO(n28640));
    SB_CARRY rem_4_add_1385_9 (.CI(n28904), .I0(n2052), .I1(VCC_net), 
            .CO(n28905));
    SB_CARRY div_46_unary_minus_2_add_3_4 (.CI(n28704), .I0(GND_net), .I1(n23_adj_4934), 
            .CO(n28705));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n28638), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4935), .I3(n28703), .O(n24_adj_4728)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_14 (.CI(n28638), .I0(n3047), .I1(VCC_net), 
            .CO(n28639));
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n28637), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_13 (.CI(n28637), .I0(n3048), .I1(VCC_net), 
            .CO(n28638));
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n28636), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_12 (.CI(n28636), .I0(n3049), .I1(VCC_net), 
            .CO(n28637));
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n28903), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_3 (.CI(n28703), .I0(GND_net), .I1(n24_adj_4935), 
            .CO(n28704));
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n28635), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_8 (.CI(n28903), .I0(n2053), .I1(VCC_net), 
            .CO(n28904));
    SB_LUT4 div_46_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4936), .I3(VCC_net), .O(n25_adj_4735)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n28902), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4936), 
            .CO(n28703));
    SB_CARRY rem_4_add_2055_11 (.CI(n28635), .I0(n3050), .I1(VCC_net), 
            .CO(n28636));
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n28634), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_10 (.CI(n28634), .I0(n3051), .I1(VCC_net), 
            .CO(n28635));
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n28633), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_9 (.CI(n28633), .I0(n3052), .I1(VCC_net), 
            .CO(n28634));
    SB_CARRY rem_4_add_1385_7 (.CI(n28902), .I0(n2054), .I1(GND_net), 
            .CO(n28903));
    SB_LUT4 div_46_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4889), .I3(n28702), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n28632), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4890), .I3(n28701), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n28901), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_6 (.CI(n28901), .I0(n2055), .I1(GND_net), 
            .CO(n28902));
    SB_CARRY div_46_unary_minus_4_add_3_24 (.CI(n28701), .I0(GND_net), .I1(n3_adj_4890), 
            .CO(n28702));
    SB_CARRY rem_4_add_2055_8 (.CI(n28632), .I0(n3053), .I1(VCC_net), 
            .CO(n28633));
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n28631), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n28900), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4891), .I3(n28700), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_7 (.CI(n28631), .I0(n3054), .I1(GND_net), 
            .CO(n28632));
    SB_CARRY div_46_unary_minus_4_add_3_23 (.CI(n28700), .I0(GND_net), .I1(n4_adj_4891), 
            .CO(n28701));
    SB_CARRY rem_4_add_1385_5 (.CI(n28900), .I0(n2056), .I1(VCC_net), 
            .CO(n28901));
    SB_LUT4 div_46_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4892), .I3(n28699), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n28899), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_22 (.CI(n28699), .I0(GND_net), .I1(n5_adj_4892), 
            .CO(n28700));
    SB_CARRY rem_4_add_1385_4 (.CI(n28899), .I0(n2057), .I1(VCC_net), 
            .CO(n28900));
    SB_LUT4 div_46_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4893), .I3(n28698), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n28630), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(n28898), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_21 (.CI(n28698), .I0(GND_net), .I1(n6_adj_4893), 
            .CO(n28699));
    SB_LUT4 div_46_i1193_3_lut_3_lut (.I0(n1778), .I1(n5975), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2055_6 (.CI(n28630), .I0(n3055), .I1(GND_net), 
            .CO(n28631));
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n28629), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_5 (.CI(n28629), .I0(n3056), .I1(VCC_net), 
            .CO(n28630));
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n28628), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_4 (.CI(n28628), .I0(n3057), .I1(VCC_net), 
            .CO(n28629));
    SB_CARRY rem_4_add_1385_3 (.CI(n28898), .I0(n2058), .I1(GND_net), 
            .CO(n28899));
    SB_LUT4 div_46_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4894), .I3(n28697), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2158), .I1(VCC_net), 
            .CO(n28898));
    SB_CARRY div_46_unary_minus_4_add_3_20 (.CI(n28697), .I0(GND_net), .I1(n7_adj_4894), 
            .CO(n28698));
    SB_LUT4 rem_4_add_1452_20_lut (.I0(n2174_adj_4975), .I1(n2141), .I2(VCC_net), 
            .I3(n28897), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1452_19_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n28896), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4895), .I3(n28696), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_19 (.CI(n28696), .I0(GND_net), .I1(n8_adj_4895), 
            .CO(n28697));
    SB_LUT4 div_46_LessThan_1606_i24_3_lut (.I0(n16_adj_5132), .I1(n91), 
            .I2(n27_adj_5141), .I3(GND_net), .O(n24_adj_5139));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35450_4_lut (.I0(n24_adj_5139), .I1(n14_adj_5130), .I2(n27_adj_5141), 
            .I3(n40351), .O(n42282));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35450_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35451_3_lut (.I0(n42282), .I1(n90), .I2(n29_adj_5142), .I3(GND_net), 
            .O(n42283));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35451_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1452_19 (.CI(n28896), .I0(n2142), .I1(VCC_net), 
            .CO(n28897));
    SB_LUT4 i35340_3_lut (.I0(n42283), .I1(n89), .I2(n31_adj_5143), .I3(GND_net), 
            .O(n42172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35340_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(n28627), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35007_4_lut (.I0(n41_adj_5149), .I1(n39_adj_5148), .I2(n37_adj_5146), 
            .I3(n40341), .O(n41839));
    defparam i35007_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35477_4_lut (.I0(n41962), .I1(n42033), .I2(n43_adj_5150), 
            .I3(n40335), .O(n42309));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35477_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35316_3_lut (.I0(n42172), .I1(n88), .I2(n33_adj_5144), .I3(GND_net), 
            .O(n42148));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35316_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4896), .I3(n28695), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35538_4_lut (.I0(n42148), .I1(n42309), .I2(n43_adj_5150), 
            .I3(n41839), .O(n42370));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35538_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n28895), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35539_3_lut (.I0(n42370), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n42371));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35539_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4905));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut (.I0(n42371), .I1(n15866), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5126));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5128));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4904));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12988_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13263), .I3(GND_net), .O(n17717));   // verilog/coms.v(126[12] 292[6])
    defparam i12988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5124));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4732), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n665));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_3 (.CI(n28627), .I0(n3058), .I1(GND_net), 
            .CO(n28628));
    SB_LUT4 div_46_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5127));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1188_3_lut_3_lut (.I0(n1778), .I1(n5970), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5121));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_DFF color__i1 (.Q(color[1]), .C(LED_c), .D(n18022));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_LUT4 div_46_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5122));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_DFF color__i2 (.Q(color[2]), .C(LED_c), .D(n18029));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_DFF color__i3 (.Q(color[3]), .C(LED_c), .D(n18030));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_DFF color__i4 (.Q(color[4]), .C(LED_c), .D(n18031));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_LUT4 i13003_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13263), .I3(GND_net), .O(n17732));   // verilog/coms.v(126[12] 292[6])
    defparam i13003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13004_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13263), .I3(GND_net), .O(n17733));   // verilog/coms.v(126[12] 292[6])
    defparam i13004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4901));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22_3_lut_adj_1714 (.I0(bit_ctr[21]), .I1(n40242), .I2(n4442), 
            .I3(GND_net), .O(n33473));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1714.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5118));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1715 (.I0(bit_ctr[20]), .I1(n40241), .I2(n4442), 
            .I3(GND_net), .O(n33471));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1715.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1716 (.I0(bit_ctr[19]), .I1(n40240), .I2(n4442), 
            .I3(GND_net), .O(n33469));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1716.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5119));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1190_3_lut_3_lut (.I0(n1778), .I1(n5972), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5120));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1717 (.I0(bit_ctr[18]), .I1(n40239), .I2(n4442), 
            .I3(GND_net), .O(n33467));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1717.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4900));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12989_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13263), .I3(GND_net), .O(n17718));   // verilog/coms.v(126[12] 292[6])
    defparam i12989_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3158), .I1(VCC_net), 
            .CO(n28627));
    SB_LUT4 rem_4_add_2122_30_lut (.I0(n3164), .I1(n3131), .I2(VCC_net), 
            .I3(n28626), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5109));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5111));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4903));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n28625), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_29 (.CI(n28625), .I0(n3132), .I1(VCC_net), 
            .CO(n28626));
    SB_LUT4 div_46_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5113));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n28624), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5115));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2122_28 (.CI(n28624), .I0(n3133), .I1(VCC_net), 
            .CO(n28625));
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n28623), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5116));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5123));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33558_4_lut (.I0(n37_adj_5123), .I1(n25_adj_5116), .I2(n23_adj_5115), 
            .I3(n21_adj_5113), .O(n40388));
    defparam i33558_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12990_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13263), .I3(GND_net), .O(n17719));   // verilog/coms.v(126[12] 292[6])
    defparam i12990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12991_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13263), .I3(GND_net), .O(n17720));   // verilog/coms.v(126[12] 292[6])
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12992_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13263), .I3(GND_net), .O(n17721));   // verilog/coms.v(126[12] 292[6])
    defparam i12992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12993_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13263), .I3(GND_net), .O(n17722));   // verilog/coms.v(126[12] 292[6])
    defparam i12993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34291_4_lut (.I0(n19_adj_5111), .I1(n17_adj_5109), .I2(n2373), 
            .I3(n98), .O(n41123));
    defparam i34291_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i12994_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13263), .I3(GND_net), .O(n17723));   // verilog/coms.v(126[12] 292[6])
    defparam i12994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34785_4_lut (.I0(n25_adj_5116), .I1(n23_adj_5115), .I2(n21_adj_5113), 
            .I3(n41123), .O(n41617));
    defparam i34785_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i12995_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13263), .I3(GND_net), .O(n17724));   // verilog/coms.v(126[12] 292[6])
    defparam i12995_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2122_27 (.CI(n28623), .I0(n3134), .I1(VCC_net), 
            .CO(n28624));
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n28622), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_26 (.CI(n28622), .I0(n3135), .I1(VCC_net), 
            .CO(n28623));
    SB_LUT4 i34781_4_lut (.I0(n31_adj_5120), .I1(n29_adj_5119), .I2(n27_adj_5118), 
            .I3(n41617), .O(n41613));
    defparam i34781_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i12996_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13263), .I3(GND_net), .O(n17725));   // verilog/coms.v(126[12] 292[6])
    defparam i12996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33567_4_lut (.I0(n37_adj_5123), .I1(n35_adj_5122), .I2(n33_adj_5121), 
            .I3(n41613), .O(n40397));
    defparam i33567_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i12997_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13263), .I3(GND_net), .O(n17726));   // verilog/coms.v(126[12] 292[6])
    defparam i12997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12998_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13263), .I3(GND_net), .O(n17727));   // verilog/coms.v(126[12] 292[6])
    defparam i12998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i14_4_lut (.I0(n665), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_5107));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4902));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35213_3_lut (.I0(n14_adj_5107), .I1(n87), .I2(n37_adj_5123), 
            .I3(GND_net), .O(n42045));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35213_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35214_3_lut (.I0(n42045), .I1(n86), .I2(n39_adj_5124), .I3(GND_net), 
            .O(n42046));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35214_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1545_i40_3_lut (.I0(n22_adj_5114), .I1(n83), 
            .I2(n45_adj_5128), .I3(GND_net), .O(n40_adj_5125));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33544_4_lut (.I0(n43_adj_5127), .I1(n41_adj_5126), .I2(n39_adj_5124), 
            .I3(n40388), .O(n40374));
    defparam i33544_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34851_4_lut (.I0(n40_adj_5125), .I1(n20_adj_5112), .I2(n45_adj_5128), 
            .I3(n40370), .O(n41683));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34851_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35126_3_lut (.I0(n42046), .I1(n85), .I2(n41_adj_5126), .I3(GND_net), 
            .O(n41958));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35126_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_46_unary_minus_4_add_3_18 (.CI(n28695), .I0(GND_net), .I1(n9_adj_4896), 
            .CO(n28696));
    SB_LUT4 div_46_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4899));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4898));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1452_18 (.CI(n28895), .I0(n2143), .I1(VCC_net), 
            .CO(n28896));
    SB_LUT4 div_46_LessThan_1545_i26_3_lut (.I0(n18_adj_5110), .I1(n91), 
            .I2(n29_adj_5119), .I3(GND_net), .O(n26_adj_5117));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35448_4_lut (.I0(n26_adj_5117), .I1(n16_adj_5108), .I2(n29_adj_5119), 
            .I3(n40427), .O(n42280));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35448_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35449_3_lut (.I0(n42280), .I1(n90), .I2(n31_adj_5120), .I3(GND_net), 
            .O(n42281));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35449_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35342_3_lut (.I0(n42281), .I1(n89), .I2(n33_adj_5121), .I3(GND_net), 
            .O(n42174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35342_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35015_4_lut (.I0(n43_adj_5127), .I1(n41_adj_5126), .I2(n39_adj_5124), 
            .I3(n40397), .O(n41847));
    defparam i35015_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35312_4_lut (.I0(n41958), .I1(n41683), .I2(n45_adj_5128), 
            .I3(n40374), .O(n42144));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35312_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35311_3_lut (.I0(n42174), .I1(n88), .I2(n35_adj_5122), .I3(GND_net), 
            .O(n42143));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35311_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35314_4_lut (.I0(n42143), .I1(n42144), .I2(n45_adj_5128), 
            .I3(n41847), .O(n42146));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35314_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n42146), .I1(n15883), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1588_3_lut_3_lut (.I0(n2381), .I1(n6079), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4897));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13005_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13263), .I3(GND_net), .O(n17734));   // verilog/coms.v(126[12] 292[6])
    defparam i13005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n28894), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5103));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5106));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5105));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(207[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n28621), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_25 (.CI(n28621), .I0(n3136), .I1(VCC_net), 
            .CO(n28622));
    SB_LUT4 div_46_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5104));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4733), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n664));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5100));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13006_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13263), .I3(GND_net), .O(n17735));   // verilog/coms.v(126[12] 292[6])
    defparam i13006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5101));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5102));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5097));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5099));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5091));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n28620), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5093));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2122_24 (.CI(n28620), .I0(n3137), .I1(VCC_net), 
            .CO(n28621));
    SB_LUT4 div_46_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5095));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5096));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13007_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13263), .I3(GND_net), .O(n17736));   // verilog/coms.v(126[12] 292[6])
    defparam i13007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n28619), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13008_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17737));   // verilog/coms.v(126[12] 292[6])
    defparam i13008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12999_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13263), .I3(GND_net), .O(n17728));   // verilog/coms.v(126[12] 292[6])
    defparam i12999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13000_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13263), .I3(GND_net), .O(n17729));   // verilog/coms.v(126[12] 292[6])
    defparam i13000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5089));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33704_4_lut (.I0(n23_adj_5095), .I1(n21_adj_5093), .I2(n19_adj_5091), 
            .I3(n17_adj_5089), .O(n40534));
    defparam i33704_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33697_4_lut (.I0(n29_adj_5099), .I1(n27_adj_5097), .I2(n25_adj_5096), 
            .I3(n40534), .O(n40527));
    defparam i33697_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35061_4_lut (.I0(n35_adj_5102), .I1(n33_adj_5101), .I2(n31_adj_5100), 
            .I3(n40527), .O(n41893));
    defparam i35061_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13009_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17738));   // verilog/coms.v(126[12] 292[6])
    defparam i13009_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1452_17 (.CI(n28894), .I0(n2144), .I1(VCC_net), 
            .CO(n28895));
    SB_LUT4 i13010_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17739));   // verilog/coms.v(126[12] 292[6])
    defparam i13010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1482_i16_4_lut (.I0(n664), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_5088));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35221_3_lut (.I0(n16_adj_5088), .I1(n87), .I2(n39_adj_5104), 
            .I3(GND_net), .O(n42053));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35221_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13011_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17740));   // verilog/coms.v(126[12] 292[6])
    defparam i13011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13001_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13263), .I3(GND_net), .O(n17730));   // verilog/coms.v(126[12] 292[6])
    defparam i13001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31_adj_4816));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1269_3_lut_3_lut (.I0(n1886), .I1(n5995), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13012_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17741));   // verilog/coms.v(126[12] 292[6])
    defparam i13012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35222_3_lut (.I0(n42053), .I1(n86), .I2(n41_adj_5105), .I3(GND_net), 
            .O(n42054));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35222_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13013_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17742));   // verilog/coms.v(126[12] 292[6])
    defparam i13013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n28893), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_16 (.CI(n28893), .I0(n2145), .I1(VCC_net), 
            .CO(n28894));
    SB_LUT4 i34303_4_lut (.I0(n41_adj_5105), .I1(n39_adj_5104), .I2(n27_adj_5097), 
            .I3(n40531), .O(n41135));
    defparam i34303_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34849_3_lut (.I0(n22_adj_5094), .I1(n93), .I2(n27_adj_5097), 
            .I3(GND_net), .O(n41681));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34849_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13014_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17743));   // verilog/coms.v(126[12] 292[6])
    defparam i13014_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13002_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13263), .I3(GND_net), .O(n17731));   // verilog/coms.v(126[12] 292[6])
    defparam i13002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35119_3_lut (.I0(n42054), .I1(n85), .I2(n43_adj_5106), .I3(GND_net), 
            .O(n41951));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35119_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1268_3_lut_3_lut (.I0(n1886), .I1(n5994), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1482_i28_3_lut (.I0(n20_adj_5092), .I1(n91), 
            .I2(n31_adj_5100), .I3(GND_net), .O(n28_adj_5098));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35443_4_lut (.I0(n28_adj_5098), .I1(n18_adj_5090), .I2(n31_adj_5100), 
            .I3(n40516), .O(n42275));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35443_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35444_3_lut (.I0(n42275), .I1(n90), .I2(n33_adj_5101), .I3(GND_net), 
            .O(n42276));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35444_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35344_3_lut (.I0(n42276), .I1(n89), .I2(n35_adj_5102), .I3(GND_net), 
            .O(n42176));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35344_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34307_4_lut (.I0(n41_adj_5105), .I1(n39_adj_5104), .I2(n37_adj_5103), 
            .I3(n41893), .O(n41139));
    defparam i34307_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35219_4_lut (.I0(n41951), .I1(n41681), .I2(n43_adj_5106), 
            .I3(n41135), .O(n42051));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35219_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_i1259_3_lut_3_lut (.I0(n1886), .I1(n5985), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35309_3_lut (.I0(n42176), .I1(n88), .I2(n37_adj_5103), .I3(GND_net), 
            .O(n42141));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35309_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35471_4_lut (.I0(n42141), .I1(n42051), .I2(n43_adj_5106), 
            .I3(n41139), .O(n42303));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35471_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35472_3_lut (.I0(n42303), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n42304));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35472_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n42304), .I1(n15880), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n28892), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_23 (.CI(n28619), .I0(n3138), .I1(VCC_net), 
            .CO(n28620));
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n28618), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_15 (.CI(n28892), .I0(n2146), .I1(VCC_net), 
            .CO(n28893));
    SB_LUT4 div_46_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4897), .I3(n28694), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_22 (.CI(n28618), .I0(n3139), .I1(VCC_net), 
            .CO(n28619));
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n28891), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_17 (.CI(n28694), .I0(GND_net), .I1(n10_adj_4897), 
            .CO(n28695));
    SB_CARRY rem_4_add_1452_14 (.CI(n28891), .I0(n2147), .I1(VCC_net), 
            .CO(n28892));
    SB_LUT4 div_46_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4898), .I3(n28693), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n28890), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_13 (.CI(n28890), .I0(n2148), .I1(VCC_net), 
            .CO(n28891));
    SB_CARRY div_46_unary_minus_4_add_3_16 (.CI(n28693), .I0(GND_net), .I1(n11_adj_4898), 
            .CO(n28694));
    SB_LUT4 div_46_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4899), .I3(n28692), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n28889), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_15 (.CI(n28692), .I0(GND_net), .I1(n12_adj_4899), 
            .CO(n28693));
    SB_CARRY rem_4_add_1452_12 (.CI(n28889), .I0(n2149), .I1(VCC_net), 
            .CO(n28890));
    SB_LUT4 i22_3_lut_adj_1720 (.I0(bit_ctr[17]), .I1(n40238), .I2(n4442), 
            .I3(GND_net), .O(n33465));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1720.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut (.I0(n40275), .I1(byte_transmit_counter[3]), .I2(n24391), 
            .I3(GND_net), .O(n34135));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1258_3_lut_3_lut (.I0(n1886), .I1(n5984), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5084));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5087));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5086));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5085));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n28888), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n28617), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_21 (.CI(n28617), .I0(n3140), .I1(VCC_net), 
            .CO(n28618));
    SB_LUT4 div_46_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4900), .I3(n28691), .O(n63_adj_4690)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_11 (.CI(n28888), .I0(n2150), .I1(VCC_net), 
            .CO(n28889));
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n28616), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_20 (.CI(n28616), .I0(n3141), .I1(VCC_net), 
            .CO(n28617));
    SB_CARRY div_46_unary_minus_4_add_3_14 (.CI(n28691), .I0(GND_net), .I1(n13_adj_4900), 
            .CO(n28692));
    SB_LUT4 div_46_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4901), .I3(n28690), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n28615), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_19 (.CI(n28615), .I0(n3142), .I1(VCC_net), 
            .CO(n28616));
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n28614), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_18 (.CI(n28614), .I0(n3143), .I1(VCC_net), 
            .CO(n28615));
    SB_LUT4 div_46_i1267_3_lut_3_lut (.I0(n1886), .I1(n5993), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5081));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5082));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n28613), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_17 (.CI(n28613), .I0(n3144), .I1(VCC_net), 
            .CO(n28614));
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n28612), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n28612), .I0(n3145), .I1(VCC_net), 
            .CO(n28613));
    SB_LUT4 div_46_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5083));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n28611), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_15 (.CI(n28611), .I0(n3146), .I1(VCC_net), 
            .CO(n28612));
    SB_LUT4 div_46_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4734), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n663));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n28610), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_14 (.CI(n28610), .I0(n3147), .I1(VCC_net), 
            .CO(n28611));
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n28609), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_13 (.CI(n28609), .I0(n3148), .I1(VCC_net), 
            .CO(n28610));
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n28608), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_12 (.CI(n28608), .I0(n3149), .I1(VCC_net), 
            .CO(n28609));
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n28607), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n28887), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_11 (.CI(n28607), .I0(n3150), .I1(VCC_net), 
            .CO(n28608));
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n28606), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_10 (.CI(n28606), .I0(n3151), .I1(VCC_net), 
            .CO(n28607));
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n28605), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_10 (.CI(n28887), .I0(n2151), .I1(VCC_net), 
            .CO(n28888));
    SB_CARRY div_46_unary_minus_4_add_3_13 (.CI(n28690), .I0(GND_net), .I1(n14_adj_4901), 
            .CO(n28691));
    SB_CARRY rem_4_add_2122_9 (.CI(n28605), .I0(n3152), .I1(VCC_net), 
            .CO(n28606));
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n28604), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_8 (.CI(n28604), .I0(n3153), .I1(VCC_net), 
            .CO(n28605));
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n28603), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_7 (.CI(n28603), .I0(n3154), .I1(GND_net), 
            .CO(n28604));
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n28602), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_6 (.CI(n28602), .I0(n3155), .I1(GND_net), 
            .CO(n28603));
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n28601), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_3_lut_adj_1721 (.I0(byte_transmit_counter[2]), .I1(n40278), 
            .I2(n24391), .I3(GND_net), .O(n34179));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut_adj_1721.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4902), .I3(n28689), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n28886), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_5 (.CI(n28601), .I0(n3156), .I1(VCC_net), 
            .CO(n28602));
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n28600), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_4 (.CI(n28600), .I0(n3157), .I1(VCC_net), 
            .CO(n28601));
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(n28599), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1270_3_lut_3_lut (.I0(n1886), .I1(n5996), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_3 (.CI(n28599), .I0(n3158), .I1(GND_net), 
            .CO(n28600));
    SB_LUT4 div_46_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5078));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5080));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5071));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1452_9 (.CI(n28886), .I0(n2152), .I1(VCC_net), 
            .CO(n28887));
    SB_CARRY div_46_unary_minus_4_add_3_12 (.CI(n28689), .I0(GND_net), .I1(n15_adj_4902), 
            .CO(n28690));
    SB_LUT4 div_46_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5073));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5075));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n28885), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5077));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5069));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33828_4_lut (.I0(n25_adj_5075), .I1(n23_adj_5073), .I2(n21_adj_5071), 
            .I3(n19_adj_5069), .O(n40660));
    defparam i33828_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33812_4_lut (.I0(n31_adj_5080), .I1(n29_adj_5078), .I2(n27_adj_5077), 
            .I3(n40660), .O(n40644));
    defparam i33812_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i1266_3_lut_3_lut (.I0(n1886), .I1(n5992), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3258), .I1(VCC_net), 
            .CO(n28599));
    SB_LUT4 i35151_4_lut (.I0(n37_adj_5083), .I1(n35_adj_5082), .I2(n33_adj_5081), 
            .I3(n40644), .O(n41983));
    defparam i35151_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1417_i18_4_lut (.I0(n663), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_5068));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4903), .I3(n28688), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_11 (.CI(n28688), .I0(GND_net), .I1(n16_adj_4903), 
            .CO(n28689));
    SB_LUT4 i35035_3_lut (.I0(n18_adj_5068), .I1(n87), .I2(n41_adj_5085), 
            .I3(GND_net), .O(n41867));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35035_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35036_3_lut (.I0(n41867), .I1(n86), .I2(n43_adj_5086), .I3(GND_net), 
            .O(n41868));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35036_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1264_3_lut_3_lut (.I0(n1886), .I1(n5990), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1265_3_lut_3_lut (.I0(n1886), .I1(n5991), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1452_8 (.CI(n28885), .I0(n2153), .I1(VCC_net), 
            .CO(n28886));
    SB_LUT4 i34451_4_lut (.I0(n43_adj_5086), .I1(n41_adj_5085), .I2(n29_adj_5078), 
            .I3(n40654), .O(n41283));
    defparam i34451_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1417_i26_3_lut (.I0(n24_adj_5074), .I1(n93), 
            .I2(n29_adj_5078), .I3(GND_net), .O(n26_adj_5076));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34410_3_lut (.I0(n41868), .I1(n85), .I2(n45_adj_5087), .I3(GND_net), 
            .O(n41242));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34410_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n28884), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_7 (.CI(n28884), .I0(n2154), .I1(GND_net), 
            .CO(n28885));
    SB_LUT4 div_46_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4904), .I3(n28687), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_10 (.CI(n28687), .I0(GND_net), .I1(n17_adj_4904), 
            .CO(n28688));
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n28883), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i30_3_lut (.I0(n22_adj_5072), .I1(n91), 
            .I2(n33_adj_5081), .I3(GND_net), .O(n30_adj_5079));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35381_4_lut (.I0(n30_adj_5079), .I1(n20_adj_5070), .I2(n33_adj_5081), 
            .I3(n40629), .O(n42213));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35381_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35382_3_lut (.I0(n42213), .I1(n90), .I2(n35_adj_5082), .I3(GND_net), 
            .O(n42214));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35382_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4905), .I3(n28686), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35263_3_lut (.I0(n42214), .I1(n89), .I2(n37_adj_5083), .I3(GND_net), 
            .O(n42095));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35263_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34457_4_lut (.I0(n43_adj_5086), .I1(n41_adj_5085), .I2(n39_adj_5084), 
            .I3(n41983), .O(n41289));
    defparam i34457_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_i1271_3_lut_3_lut (.I0(n1886), .I1(n5997), .I2(n660), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1452_6 (.CI(n28883), .I0(n2155), .I1(GND_net), 
            .CO(n28884));
    SB_LUT4 i35111_4_lut (.I0(n41242), .I1(n26_adj_5076), .I2(n45_adj_5087), 
            .I3(n41283), .O(n41943));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35111_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34408_3_lut (.I0(n42095), .I1(n88), .I2(n39_adj_5084), .I3(GND_net), 
            .O(n41240));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34408_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35113_4_lut (.I0(n41240), .I1(n41943), .I2(n45_adj_5087), 
            .I3(n41289), .O(n41945));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35113_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i1263_3_lut_3_lut (.I0(n1886), .I1(n5989), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n41945), .I1(n15812), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i1659_3_lut (.I0(n2442), .I1(n2509), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2541_adj_4883));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1657_3_lut (.I0(n2440), .I1(n2507), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2539_adj_4885));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1261_3_lut_3_lut (.I0(n1886), .I1(n5987), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1262_3_lut_3_lut (.I0(n1886), .I1(n5988), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1670_3_lut (.I0(n2453_adj_4943), .I1(n2520), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2552_adj_4872));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n28882), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_5 (.CI(n28882), .I0(n2156), .I1(VCC_net), 
            .CO(n28883));
    SB_LUT4 rem_4_i1668_3_lut (.I0(n2451_adj_4945), .I1(n2518), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2550_adj_4874));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_9 (.CI(n28686), .I0(GND_net), .I1(n18_adj_4905), 
            .CO(n28687));
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n28881), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4906), .I3(n28685), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_8 (.CI(n28685), .I0(GND_net), .I1(n19_adj_4906), 
            .CO(n28686));
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4907), .I3(n28684), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1666_3_lut (.I0(n2449_adj_4947), .I1(n2516), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2548_adj_4876));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1260_3_lut_3_lut (.I0(n1886), .I1(n5986), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1662_3_lut (.I0(n2445), .I1(n2512), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2544_adj_4880));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_4 (.CI(n28881), .I0(n2157), .I1(VCC_net), 
            .CO(n28882));
    SB_LUT4 rem_4_i1667_3_lut (.I0(n2450_adj_4946), .I1(n2517), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2549_adj_4875));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1663_3_lut (.I0(n2446), .I1(n2513), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2545_adj_4879));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1673_3_lut (.I0(n2456_adj_4940), .I1(n2523), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2555));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1661_3_lut (.I0(n2444), .I1(n2511), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2543_adj_4881));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1672_3_lut (.I0(n2455_adj_4941), .I1(n2522), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2554));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1665_3_lut (.I0(n2448_adj_4948), .I1(n2515), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2547_adj_4877));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1671_3_lut (.I0(n2454_adj_4942), .I1(n2521), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2553_adj_4871));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1669_3_lut (.I0(n2452_adj_4944), .I1(n2519), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2551_adj_4873));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1664_3_lut (.I0(n2447_adj_4949), .I1(n2514), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2546_adj_4878));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1660_3_lut (.I0(n2443), .I1(n2510), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2542_adj_4882));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1658_3_lut (.I0(n2441), .I1(n2508), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2540_adj_4884));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1656_3_lut (.I0(n2439), .I1(n2506), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2538_adj_4886));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1675_3_lut (.I0(n2458_adj_4938), .I1(n2525), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2557));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1674_3_lut (.I0(n2457_adj_4939), .I1(n2524), .I2(n2471_adj_4937), 
            .I3(GND_net), .O(n2556));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut (.I0(n31_adj_4816), .I1(n2739), .I2(n24_adj_4817), 
            .I3(n2740), .O(n36_adj_4799));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n2556), .I1(n2557), .I2(n2558_adj_4870), .I3(GND_net), 
            .O(n35595));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i10_4_lut (.I0(n2538_adj_4886), .I1(n2540_adj_4884), .I2(n2537_adj_4887), 
            .I3(n2542_adj_4882), .O(n28_adj_5269));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2546_adj_4878), .I1(n2551_adj_4873), .I2(n2553_adj_4871), 
            .I3(n2547_adj_4877), .O(n31_adj_5267));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n2554), .I1(n2543_adj_4881), .I2(n35595), .I3(n2555), 
            .O(n22_adj_5270));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i12_4_lut (.I0(n2545_adj_4879), .I1(n2549_adj_4875), .I2(n2544_adj_4880), 
            .I3(n2548_adj_4876), .O(n30_adj_5268));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1723 (.I0(n31_adj_5267), .I1(n2550_adj_4874), 
            .I2(n28_adj_5269), .I3(n2552_adj_4872), .O(n34_adj_5266));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(n28880), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_7 (.CI(n28684), .I0(GND_net), .I1(n20_adj_4907), 
            .CO(n28685));
    SB_LUT4 i3_2_lut (.I0(n2539_adj_4885), .I1(n2541_adj_4883), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5271));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i17_4_lut (.I0(n21_adj_5271), .I1(n34_adj_5266), .I2(n30_adj_5268), 
            .I3(n22_adj_5270), .O(n2570));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4771), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558_adj_4870));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4908), .I3(n28683), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_3 (.CI(n28880), .I0(n2158), .I1(GND_net), 
            .CO(n28881));
    SB_CARRY div_46_unary_minus_4_add_3_6 (.CI(n28683), .I0(GND_net), .I1(n21_adj_4908), 
            .CO(n28684));
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2258), .I1(VCC_net), 
            .CO(n28880));
    SB_LUT4 div_46_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5067));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5066));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_21_lut (.I0(n2273_adj_4962), .I1(n2240), .I2(VCC_net), 
            .I3(n28879), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5065));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_20_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n28878), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4909), .I3(n28682), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_20 (.CI(n28878), .I0(n2241), .I1(VCC_net), 
            .CO(n28879));
    SB_LUT4 div_46_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5064));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n28877), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_5 (.CI(n28682), .I0(GND_net), .I1(n22_adj_4909), 
            .CO(n28683));
    SB_LUT4 div_46_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4910), .I3(n28681), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_4 (.CI(n28681), .I0(GND_net), .I1(n23_adj_4910), 
            .CO(n28682));
    SB_LUT4 div_46_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4911), .I3(n28680), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_3 (.CI(n28680), .I0(GND_net), .I1(n24_adj_4911), 
            .CO(n28681));
    SB_CARRY rem_4_add_1519_19 (.CI(n28877), .I0(n2242), .I1(VCC_net), 
            .CO(n28878));
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n28876), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4726), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n662));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4912), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4912), 
            .CO(n28680));
    SB_CARRY rem_4_add_1519_18 (.CI(n28876), .I0(n2243), .I1(VCC_net), 
            .CO(n28877));
    SB_LUT4 rem_4_add_1988_28_lut (.I0(n2966_adj_4798), .I1(n2933), .I2(VCC_net), 
            .I3(n28679), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_27_lut (.I0(GND_net), .I1(n2934), .I2(VCC_net), 
            .I3(n28678), .O(n3001_adj_4796)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_27 (.CI(n28678), .I0(n2934), .I1(VCC_net), 
            .CO(n28679));
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n28875), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_26_lut (.I0(GND_net), .I1(n2935), .I2(VCC_net), 
            .I3(n28677), .O(n3002_adj_4795)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_26 (.CI(n28677), .I0(n2935), .I1(VCC_net), 
            .CO(n28678));
    SB_LUT4 rem_4_add_1988_25_lut (.I0(GND_net), .I1(n2936), .I2(VCC_net), 
            .I3(n28676), .O(n3003_adj_4794)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_17 (.CI(n28875), .I0(n2244), .I1(VCC_net), 
            .CO(n28876));
    SB_CARRY rem_4_add_1988_25 (.CI(n28676), .I0(n2936), .I1(VCC_net), 
            .CO(n28677));
    SB_LUT4 rem_4_add_1988_24_lut (.I0(GND_net), .I1(n2937), .I2(VCC_net), 
            .I3(n28675), .O(n3004_adj_4793)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n28874), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_24 (.CI(n28675), .I0(n2937), .I1(VCC_net), 
            .CO(n28676));
    SB_LUT4 rem_4_add_1988_23_lut (.I0(GND_net), .I1(n2938), .I2(VCC_net), 
            .I3(n28674), .O(n3005_adj_4792)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_16 (.CI(n28874), .I0(n2245), .I1(VCC_net), 
            .CO(n28875));
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n28873), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_15 (.CI(n28873), .I0(n2246), .I1(VCC_net), 
            .CO(n28874));
    SB_CARRY rem_4_add_1988_23 (.CI(n28674), .I0(n2938), .I1(VCC_net), 
            .CO(n28675));
    SB_LUT4 div_46_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5054));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5056));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n28872), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_14 (.CI(n28872), .I0(n2247), .I1(VCC_net), 
            .CO(n28873));
    SB_LUT4 rem_4_add_1988_22_lut (.I0(GND_net), .I1(n2939), .I2(VCC_net), 
            .I3(n28673), .O(n3006_adj_4791)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5058));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n28871), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_22 (.CI(n28673), .I0(n2939), .I1(VCC_net), 
            .CO(n28674));
    SB_CARRY rem_4_add_1519_13 (.CI(n28871), .I0(n2248), .I1(VCC_net), 
            .CO(n28872));
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n28870), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_21_lut (.I0(GND_net), .I1(n2940), .I2(VCC_net), 
            .I3(n28672), .O(n3007_adj_4790)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2058_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), .I3(GND_net), 
            .O(n3132));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_21 (.CI(n28672), .I0(n2940), .I1(VCC_net), 
            .CO(n28673));
    SB_LUT4 div_46_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5060));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2077_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_20_lut (.I0(GND_net), .I1(n2941), .I2(VCC_net), 
            .I3(n28671), .O(n3008_adj_4789)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5061));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_12 (.CI(n28870), .I0(n2249), .I1(VCC_net), 
            .CO(n28871));
    SB_CARRY rem_4_add_1988_20 (.CI(n28671), .I0(n2941), .I1(VCC_net), 
            .CO(n28672));
    SB_LUT4 rem_4_i2076_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n28869), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_11 (.CI(n28869), .I0(n2250), .I1(VCC_net), 
            .CO(n28870));
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n28868), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_19_lut (.I0(GND_net), .I1(n2942), .I2(VCC_net), 
            .I3(n28670), .O(n3009_adj_4788)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5063));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1519_10 (.CI(n28868), .I0(n2251), .I1(VCC_net), 
            .CO(n28869));
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n28867), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1988_19 (.CI(n28670), .I0(n2942), .I1(VCC_net), 
            .CO(n28671));
    SB_CARRY rem_4_add_1519_9 (.CI(n28867), .I0(n2252), .I1(VCC_net), 
            .CO(n28868));
    SB_LUT4 rem_4_add_1988_18_lut (.I0(GND_net), .I1(n2943), .I2(VCC_net), 
            .I3(n28669), .O(n3010_adj_4787)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_18 (.CI(n28669), .I0(n2943), .I1(VCC_net), 
            .CO(n28670));
    SB_LUT4 rem_4_add_1988_17_lut (.I0(GND_net), .I1(n2944), .I2(VCC_net), 
            .I3(n28668), .O(n3011_adj_4786)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n28866), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5052));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33922_4_lut (.I0(n27_adj_5058), .I1(n25_adj_5056), .I2(n23_adj_5054), 
            .I3(n21_adj_5052), .O(n40754));
    defparam i33922_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1988_17 (.CI(n28668), .I0(n2944), .I1(VCC_net), 
            .CO(n28669));
    SB_CARRY rem_4_add_1519_8 (.CI(n28866), .I0(n2253), .I1(VCC_net), 
            .CO(n28867));
    SB_LUT4 rem_4_add_1988_16_lut (.I0(GND_net), .I1(n2945_adj_4815), .I2(VCC_net), 
            .I3(n28667), .O(n3012_adj_4785)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n28865), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33907_4_lut (.I0(n33_adj_5063), .I1(n31_adj_5061), .I2(n29_adj_5060), 
            .I3(n40754), .O(n40739));
    defparam i33907_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1988_16 (.CI(n28667), .I0(n2945_adj_4815), .I1(VCC_net), 
            .CO(n28668));
    SB_LUT4 rem_4_add_1988_15_lut (.I0(GND_net), .I1(n2946_adj_4814), .I2(VCC_net), 
            .I3(n28666), .O(n3013_adj_4784)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_7 (.CI(n28865), .I0(n2254), .I1(GND_net), 
            .CO(n28866));
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i20_4_lut (.I0(n662), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_5051));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1350_i28_3_lut (.I0(n26_adj_5057), .I1(n93), 
            .I2(n31_adj_5061), .I3(GND_net), .O(n28_adj_5059));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1585_3_lut_3_lut (.I0(n2381), .I1(n6076), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2069_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), .I3(GND_net), 
            .O(n3143));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n28864), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_15 (.CI(n28666), .I0(n2946_adj_4814), .I1(VCC_net), 
            .CO(n28667));
    SB_LUT4 rem_4_i2075_3_lut (.I0(n3050), .I1(n3117), .I2(n3065), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_14_lut (.I0(GND_net), .I1(n2947_adj_4813), .I2(VCC_net), 
            .I3(n28665), .O(n3014_adj_4783)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i32_3_lut (.I0(n24_adj_5055), .I1(n91), 
            .I2(n35_adj_5064), .I3(GND_net), .O(n32_adj_5062));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35377_4_lut (.I0(n32_adj_5062), .I1(n22_adj_5053), .I2(n35_adj_5064), 
            .I3(n40734), .O(n42209));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35377_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35378_3_lut (.I0(n42209), .I1(n90), .I2(n37_adj_5065), .I3(GND_net), 
            .O(n42210));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35378_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35267_3_lut (.I0(n42210), .I1(n89), .I2(n39_adj_5066), .I3(GND_net), 
            .O(n42099));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35267_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35159_4_lut (.I0(n39_adj_5066), .I1(n37_adj_5065), .I2(n35_adj_5064), 
            .I3(n40739), .O(n41991));
    defparam i35159_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35441_4_lut (.I0(n28_adj_5059), .I1(n20_adj_5051), .I2(n31_adj_5061), 
            .I3(n40746), .O(n42273));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35441_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_1519_6 (.CI(n28864), .I0(n2255), .I1(GND_net), 
            .CO(n28865));
    SB_LUT4 i34404_3_lut (.I0(n42099), .I1(n88), .I2(n41_adj_5067), .I3(GND_net), 
            .O(n41236));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34404_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35534_4_lut (.I0(n41236), .I1(n42273), .I2(n41_adj_5067), 
            .I3(n41991), .O(n42366));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35534_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35535_3_lut (.I0(n42366), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n42367));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35535_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35484_3_lut (.I0(n42367), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n42316));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35484_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_i2071_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n28863), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n42316), .I1(n15863), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_14 (.CI(n28665), .I0(n2947_adj_4813), .I1(VCC_net), 
            .CO(n28666));
    SB_LUT4 div_46_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5050));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5048));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5049));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5047));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1994_3_lut (.I0(n2937), .I1(n3004_adj_4793), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3036));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1993_3_lut (.I0(n2936), .I1(n3003_adj_4794), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3035));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4727), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n661));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1992_3_lut (.I0(n2935), .I1(n3002_adj_4795), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3034));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1995_3_lut (.I0(n2938), .I1(n3005_adj_4792), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3037));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut (.I0(n40226), .I1(bit_ctr[1]), .I2(n4442), .I3(GND_net), 
            .O(n33435));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5043));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1519_5 (.CI(n28863), .I0(n2256), .I1(VCC_net), 
            .CO(n28864));
    SB_LUT4 rem_4_i1996_3_lut (.I0(n2939), .I1(n3006_adj_4791), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3038));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n28862), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5044));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_13_lut (.I0(GND_net), .I1(n2948_adj_4812), .I2(VCC_net), 
            .I3(n28664), .O(n3015_adj_4671)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_13 (.CI(n28664), .I0(n2948_adj_4812), .I1(VCC_net), 
            .CO(n28665));
    SB_LUT4 rem_4_i1991_3_lut (.I0(n2934), .I1(n3001_adj_4796), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_4 (.CI(n28862), .I0(n2257), .I1(VCC_net), 
            .CO(n28863));
    SB_LUT4 rem_4_add_1988_12_lut (.I0(GND_net), .I1(n2949_adj_4811), .I2(VCC_net), 
            .I3(n28663), .O(n3016_adj_4764)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_55 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 i1_3_lut_adj_1725 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n35687));
    defparam i1_3_lut_adj_1725.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut (.I0(n3042), .I1(n3054), .I2(n35687), .I3(n3055), 
            .O(n30_adj_5254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut.LUT_INIT = 16'heaaa;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14_4_lut (.I0(n3038), .I1(n3048), .I2(n3037), .I3(n3040), 
            .O(n37_adj_5252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5046));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13_4_lut_adj_1726 (.I0(n3034), .I1(n3039), .I2(n3035), .I3(n3036), 
            .O(n36_adj_5253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(n28861), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut (.I0(n37_adj_5252), .I1(n3046), .I2(n30_adj_5254), 
            .I3(n3041), .O(n42_adj_5247));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5037));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i17_4_lut_adj_1727 (.I0(n3051), .I1(n3045), .I2(n3053), .I3(n3049), 
            .O(n40_adj_5249));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut_adj_1727.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1519_3 (.CI(n28861), .I0(n2258), .I1(GND_net), 
            .CO(n28862));
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4953), .I1(VCC_net), 
            .CO(n28861));
    SB_LUT4 i18_4_lut (.I0(n3047), .I1(n36_adj_5253), .I2(n3033), .I3(n3032), 
            .O(n41_adj_5248));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1988_12 (.CI(n28663), .I0(n2949_adj_4811), .I1(VCC_net), 
            .CO(n28664));
    SB_LUT4 i16_4_lut_adj_1728 (.I0(n3043), .I1(n3050), .I2(n3044), .I3(n3052), 
            .O(n39_adj_5250));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_5250), .I1(n41_adj_5248), .I2(n40_adj_5249), 
            .I3(n42_adj_5247), .O(n3065));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1988_11_lut (.I0(GND_net), .I1(n2950_adj_4810), .I2(VCC_net), 
            .I3(n28662), .O(n3017_adj_4763)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5039));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_11 (.CI(n28662), .I0(n2950_adj_4810), .I1(VCC_net), 
            .CO(n28663));
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1586_22_lut (.I0(n2372_adj_4952), .I1(n2339), .I2(VCC_net), 
            .I3(n28860), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5041));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1729 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n35635));
    defparam i1_3_lut_adj_1729.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5035));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4896));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1730 (.I0(n3141), .I1(n3145), .I2(n3142), .I3(n3146), 
            .O(n40));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1988_10_lut (.I0(GND_net), .I1(n2951_adj_4809), .I2(VCC_net), 
            .I3(n28661), .O(n3018_adj_4762)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33970_4_lut (.I0(n29_adj_5041), .I1(n27_adj_5039), .I2(n25_adj_5037), 
            .I3(n23_adj_5035), .O(n40802));
    defparam i33970_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i1340_3_lut_3_lut (.I0(n1991), .I1(n6013), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i5_4_lut (.I0(n3139), .I1(n3154), .I2(n35635), .I3(n3155), 
            .O(n29));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i33960_4_lut (.I0(n35_adj_5046), .I1(n33_adj_5044), .I2(n31_adj_5043), 
            .I3(n40802), .O(n40792));
    defparam i33960_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_1586_21_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n28859), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4797));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_1988_10 (.CI(n28661), .I0(n2951_adj_4809), .I1(VCC_net), 
            .CO(n28662));
    SB_CARRY rem_4_add_1586_21 (.CI(n28859), .I0(n2340), .I1(VCC_net), 
            .CO(n28860));
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n28858), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_9_lut (.I0(GND_net), .I1(n2952_adj_4808), .I2(VCC_net), 
            .I3(n28660), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_9 (.CI(n28660), .I0(n2952_adj_4808), .I1(VCC_net), 
            .CO(n28661));
    SB_LUT4 rem_4_add_1988_8_lut (.I0(GND_net), .I1(n2953_adj_4807), .I2(VCC_net), 
            .I3(n28659), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_20 (.CI(n28858), .I0(n2341), .I1(VCC_net), 
            .CO(n28859));
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n28857), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_8 (.CI(n28659), .I0(n2953_adj_4807), .I1(VCC_net), 
            .CO(n28660));
    SB_LUT4 div_46_LessThan_1281_i22_4_lut (.I0(n661), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_5034));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i14_4_lut_adj_1731 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1331_3_lut_3_lut (.I0(n1991), .I1(n6004), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i20_4_lut (.I0(n29), .I1(n40), .I2(n3140), .I3(n3150), .O(n44));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 rem_4_add_1988_7_lut (.I0(GND_net), .I1(n2954_adj_4806), .I2(GND_net), 
            .I3(n28658), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18_4_lut_adj_1732 (.I0(n3148), .I1(n3144), .I2(n3151), .I3(n3153), 
            .O(n42));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1281_i30_3_lut (.I0(n28_adj_5040), .I1(n93), 
            .I2(n33_adj_5044), .I3(GND_net), .O(n30_adj_5042));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1586_19 (.CI(n28857), .I0(n2342), .I1(VCC_net), 
            .CO(n28858));
    SB_CARRY rem_4_add_1988_7 (.CI(n28658), .I0(n2954_adj_4806), .I1(GND_net), 
            .CO(n28659));
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n28856), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_6_lut (.I0(GND_net), .I1(n2955_adj_4805), .I2(GND_net), 
            .I3(n28657), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_18 (.CI(n28856), .I0(n2343), .I1(VCC_net), 
            .CO(n28857));
    SB_CARRY rem_4_add_1988_6 (.CI(n28657), .I0(n2955_adj_4805), .I1(GND_net), 
            .CO(n28658));
    SB_LUT4 i19_4_lut_adj_1733 (.I0(n3132), .I1(n38), .I2(n26_adj_4797), 
            .I3(n3131), .O(n43));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n28855), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_17 (.CI(n28855), .I0(n2344), .I1(VCC_net), 
            .CO(n28856));
    SB_LUT4 rem_4_add_1988_5_lut (.I0(GND_net), .I1(n2956_adj_4804), .I2(VCC_net), 
            .I3(n28656), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n28656), .I0(n2956_adj_4804), .I1(VCC_net), 
            .CO(n28657));
    SB_LUT4 rem_4_add_1988_4_lut (.I0(GND_net), .I1(n2957_adj_4803), .I2(VCC_net), 
            .I3(n28655), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut_adj_1734 (.I0(n3147), .I1(n3149), .I2(n3152), .I3(n3143), 
            .O(n41));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n28854), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n28854), .I0(n2345), .I1(VCC_net), 
            .CO(n28855));
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n28853), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n3164));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4766), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1328_3_lut_3_lut (.I0(n1991), .I1(n6001), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1330_3_lut_3_lut (.I0(n1991), .I1(n6003), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1281_i34_3_lut (.I0(n26_adj_5038), .I1(n91), 
            .I2(n37_adj_5047), .I3(GND_net), .O(n34_adj_5045));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35375_4_lut (.I0(n34_adj_5045), .I1(n24_adj_5036), .I2(n37_adj_5047), 
            .I3(n40786), .O(n42207));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35375_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35376_3_lut (.I0(n42207), .I1(n90), .I2(n39_adj_5048), .I3(GND_net), 
            .O(n42208));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35376_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35269_3_lut (.I0(n42208), .I1(n89), .I2(n41_adj_5049), .I3(GND_net), 
            .O(n42101));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35269_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35165_4_lut (.I0(n41_adj_5049), .I1(n39_adj_5048), .I2(n37_adj_5047), 
            .I3(n40792), .O(n41997));
    defparam i35165_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35227_4_lut (.I0(n30_adj_5042), .I1(n22_adj_5034), .I2(n33_adj_5044), 
            .I3(n40798), .O(n42059));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35227_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34400_3_lut (.I0(n42101), .I1(n88), .I2(n43_adj_5050), .I3(GND_net), 
            .O(n41232));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34400_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35349_4_lut (.I0(n41232), .I1(n42059), .I2(n43_adj_5050), 
            .I3(n41997), .O(n42181));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35349_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35350_3_lut (.I0(n42181), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n42182));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35350_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i1329_3_lut_3_lut (.I0(n1991), .I1(n6002), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n42182), .I1(n15860), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5029));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1327_3_lut_3_lut (.I0(n1991), .I1(n6000), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1586_3_lut_3_lut (.I0(n2381), .I1(n6077), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4721), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n660));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5028));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5032));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5022));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5024));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5026));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5031));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1736 (.I0(n2744), .I1(n2745), .I2(n2746), .I3(n2751), 
            .O(n34_adj_4800));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5020));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34024_4_lut (.I0(n31_adj_5026), .I1(n29_adj_5024), .I2(n27_adj_5022), 
            .I3(n25_adj_5020), .O(n40856));
    defparam i34024_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i1336_3_lut_3_lut (.I0(n1991), .I1(n6009), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1988_4 (.CI(n28655), .I0(n2957_adj_4803), .I1(VCC_net), 
            .CO(n28656));
    SB_CARRY rem_4_add_1586_15 (.CI(n28853), .I0(n2346), .I1(VCC_net), 
            .CO(n28854));
    SB_LUT4 div_46_LessThan_1210_i36_3_lut (.I0(n28_adj_5023), .I1(n91), 
            .I2(n39_adj_5032), .I3(GND_net), .O(n36_adj_5030));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1210_i24_4_lut (.I0(n660), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_5019));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1210_i32_3_lut (.I0(n30_adj_5025), .I1(n93), 
            .I2(n35_adj_5029), .I3(GND_net), .O(n32_adj_5027));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34013_4_lut (.I0(n37_adj_5031), .I1(n35_adj_5029), .I2(n33_adj_5028), 
            .I3(n40856), .O(n40845));
    defparam i34013_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35373_4_lut (.I0(n36_adj_5030), .I1(n26_adj_5021), .I2(n39_adj_5032), 
            .I3(n40841), .O(n42205));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35373_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34839_4_lut (.I0(n32_adj_5027), .I1(n24_adj_5019), .I2(n35_adj_5029), 
            .I3(n40852), .O(n41671));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34839_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35512_4_lut (.I0(n41671), .I1(n42205), .I2(n39_adj_5032), 
            .I3(n40845), .O(n42344));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35512_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35513_3_lut (.I0(n42344), .I1(n90), .I2(n1865), .I3(GND_net), 
            .O(n42345));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35513_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_983_12_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n27890), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i35464_3_lut (.I0(n42345), .I1(n89), .I2(n1864), .I3(GND_net), 
            .O(n42296));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35464_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n27889), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_11 (.CI(n27889), .I0(n1449), .I1(VCC_net), 
            .CO(n27890));
    SB_LUT4 i35105_3_lut (.I0(n42296), .I1(n88), .I2(n1863), .I3(GND_net), 
            .O(n41937));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35105_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n41937), .I1(n15808), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1655_3_lut_3_lut (.I0(n2471), .I1(n6108), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5015));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_3_lut (.I0(GND_net), .I1(n2958_adj_4802), .I2(GND_net), 
            .I3(n28654), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5014));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1334_3_lut_3_lut (.I0(n1991), .I1(n6007), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4722), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n659));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5018));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5017));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n28852), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n28654), .I0(n2958_adj_4802), .I1(GND_net), 
            .CO(n28655));
    SB_LUT4 div_46_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5010));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1642_3_lut_3_lut (.I0(n2471), .I1(n6095), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5012));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5013));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n27888), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5008));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34068_4_lut (.I0(n33_adj_5013), .I1(n31_adj_5012), .I2(n29_adj_5010), 
            .I3(n27_adj_5008), .O(n40900));
    defparam i34068_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n3058), .I1(VCC_net), 
            .CO(n28654));
    SB_CARRY rem_4_add_1586_14 (.CI(n28852), .I0(n2347), .I1(VCC_net), 
            .CO(n28853));
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n28851), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1335_3_lut_3_lut (.I0(n1991), .I1(n6008), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2055_29_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n28653), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1586_13 (.CI(n28851), .I0(n2348), .I1(VCC_net), 
            .CO(n28852));
    SB_LUT4 rem_4_add_2055_28_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n28652), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i38_3_lut (.I0(n30_adj_5011), .I1(n91), 
            .I2(n41_adj_5018), .I3(GND_net), .O(n38_adj_5016));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1137_i26_4_lut (.I0(n659), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_5007));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35051_3_lut (.I0(n26_adj_5007), .I1(n95), .I2(n33_adj_5013), 
            .I3(GND_net), .O(n41883));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35051_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35052_3_lut (.I0(n41883), .I1(n94), .I2(n35_adj_5014), .I3(GND_net), 
            .O(n41884));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35052_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34052_4_lut (.I0(n39_adj_5017), .I1(n37_adj_5015), .I2(n35_adj_5014), 
            .I3(n40900), .O(n40884));
    defparam i34052_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35369_4_lut (.I0(n38_adj_5016), .I1(n28_adj_5009), .I2(n41_adj_5018), 
            .I3(n40876), .O(n42201));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34386_3_lut (.I0(n41884), .I1(n93), .I2(n37_adj_5015), .I3(GND_net), 
            .O(n41218));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34386_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35532_4_lut (.I0(n41218), .I1(n42201), .I2(n41_adj_5018), 
            .I3(n40884), .O(n42364));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35533_3_lut (.I0(n42364), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n42365));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35533_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35488_3_lut (.I0(n42365), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n42320));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35488_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n42320), .I1(n15857), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n28850), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_28 (.CI(n28652), .I0(n3033), .I1(VCC_net), 
            .CO(n28653));
    SB_LUT4 div_46_i1339_3_lut_3_lut (.I0(n1991), .I1(n6012), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1586_12 (.CI(n28850), .I0(n2349), .I1(VCC_net), 
            .CO(n28851));
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n28651), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n28849), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_27 (.CI(n28651), .I0(n3034), .I1(VCC_net), 
            .CO(n28652));
    SB_LUT4 div_46_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5003));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2189_31_lut (.I0(n3230), .I1(n3230), .I2(n3263), 
            .I3(n28534), .O(n3329)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_31_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_2189_30_lut (.I0(n3231), .I1(n3231), .I2(n3263), 
            .I3(n28533), .O(n3330)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5002));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2189_30 (.CI(n28533), .I0(n3231), .I1(n3263), .CO(n28534));
    SB_CARRY rem_4_add_1586_11 (.CI(n28849), .I0(n2350), .I1(VCC_net), 
            .CO(n28850));
    SB_LUT4 div_46_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5006));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n28650), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_29_lut (.I0(n3232), .I1(n3232), .I2(n3263), 
            .I3(n28532), .O(n3331)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4723), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n658));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5005));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4998));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5000));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5001));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4996));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1643_3_lut_3_lut (.I0(n2471), .I1(n6096), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1644_3_lut_3_lut (.I0(n2471), .I1(n6097), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34107_4_lut (.I0(n35_adj_5001), .I1(n33_adj_5000), .I2(n31_adj_4998), 
            .I3(n29_adj_4996), .O(n40939));
    defparam i34107_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_2189_29 (.CI(n28532), .I0(n3232), .I1(n3263), .CO(n28533));
    SB_LUT4 div_46_LessThan_1062_i40_3_lut (.I0(n32_adj_4999), .I1(n91), 
            .I2(n43_adj_5006), .I3(GND_net), .O(n40_adj_5004));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1062_i28_4_lut (.I0(n658), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4995));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n28848), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_26 (.CI(n28650), .I0(n3035), .I1(VCC_net), 
            .CO(n28651));
    SB_LUT4 i35055_3_lut (.I0(n28_adj_4995), .I1(n95), .I2(n35_adj_5001), 
            .I3(GND_net), .O(n41887));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35055_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1338_3_lut_3_lut (.I0(n1991), .I1(n6011), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35056_3_lut (.I0(n41887), .I1(n94), .I2(n37_adj_5002), .I3(GND_net), 
            .O(n41888));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35056_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2189_28_lut (.I0(n3233), .I1(n3233), .I2(n3263), 
            .I3(n28531), .O(n3332)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_28 (.CI(n28531), .I0(n3233), .I1(n3263), .CO(n28532));
    SB_LUT4 i34101_4_lut (.I0(n41_adj_5005), .I1(n39_adj_5003), .I2(n37_adj_5002), 
            .I3(n40939), .O(n40933));
    defparam i34101_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_2189_27_lut (.I0(n3234), .I1(n3234), .I2(n3263), 
            .I3(n28530), .O(n3333)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_i1647_3_lut_3_lut (.I0(n2471), .I1(n6100), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35351_4_lut (.I0(n40_adj_5004), .I1(n30_adj_4997), .I2(n43_adj_5006), 
            .I3(n40931), .O(n42183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35351_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_i1645_3_lut_3_lut (.I0(n2471), .I1(n6098), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1648_3_lut_3_lut (.I0(n2471), .I1(n6101), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34384_3_lut (.I0(n41888), .I1(n93), .I2(n39_adj_5003), .I3(GND_net), 
            .O(n41216));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34384_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_983_10 (.CI(n27888), .I0(n1450), .I1(VCC_net), 
            .CO(n27889));
    SB_LUT4 i35522_4_lut (.I0(n41216), .I1(n42183), .I2(n43_adj_5006), 
            .I3(n40933), .O(n42354));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35522_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35523_3_lut (.I0(n42354), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n42355));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35523_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i1661_3_lut_3_lut (.I0(n2471), .I1(n6114), .I2(n666), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1646_3_lut_3_lut (.I0(n2471), .I1(n6099), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_27 (.CI(n28530), .I0(n3234), .I1(n3263), .CO(n28531));
    SB_LUT4 i13206_3_lut (.I0(\data_in_frame[24] [0]), .I1(rx_data[0]), 
            .I2(n36887), .I3(GND_net), .O(n17935));   // verilog/coms.v(126[12] 292[6])
    defparam i13206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n42355), .I1(n15804), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hceef;
    SB_LUT4 i13216_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17945));   // verilog/coms.v(126[12] 292[6])
    defparam i13216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13215_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17944));   // verilog/coms.v(126[12] 292[6])
    defparam i13215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13214_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17943));   // verilog/coms.v(126[12] 292[6])
    defparam i13214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n28649), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1650_3_lut_3_lut (.I0(n2471), .I1(n6103), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4989));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4990));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13218_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17947));   // verilog/coms.v(126[12] 292[6])
    defparam i13218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13217_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17946));   // verilog/coms.v(126[12] 292[6])
    defparam i13217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_26_lut (.I0(n3235), .I1(n3235), .I2(n3263), 
            .I3(n28529), .O(n3334)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hCA3A;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1651_3_lut_3_lut (.I0(n2471), .I1(n6104), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1586_10 (.CI(n28848), .I0(n2351), .I1(VCC_net), 
            .CO(n28849));
    SB_CARRY rem_4_add_2055_25 (.CI(n28649), .I0(n3036), .I1(VCC_net), 
            .CO(n28650));
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n28847), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n28648), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_24 (.CI(n28648), .I0(n3037), .I1(VCC_net), 
            .CO(n28649));
    SB_LUT4 i13220_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17949));   // verilog/coms.v(126[12] 292[6])
    defparam i13220_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_26 (.CI(n28529), .I0(n3235), .I1(n3263), .CO(n28530));
    SB_LUT4 rem_4_add_2189_25_lut (.I0(n3236), .I1(n3236), .I2(n3263), 
            .I3(n28528), .O(n3335)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13219_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17948));   // verilog/coms.v(126[12] 292[6])
    defparam i13219_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_25 (.CI(n28528), .I0(n3236), .I1(n3263), .CO(n28529));
    SB_LUT4 rem_4_add_2189_24_lut (.I0(n3237), .I1(n3237), .I2(n3263), 
            .I3(n28527), .O(n3336)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_24 (.CI(n28527), .I0(n3237), .I1(n3263), .CO(n28528));
    SB_LUT4 div_46_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4724), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n657));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_23_lut (.I0(n3238), .I1(n3238), .I2(n3263), 
            .I3(n28526), .O(n3337)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_23 (.CI(n28526), .I0(n3238), .I1(n3263), .CO(n28527));
    SB_LUT4 rem_4_add_2189_22_lut (.I0(n3239), .I1(n3239), .I2(n3263), 
            .I3(n28525), .O(n3338)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_22 (.CI(n28525), .I0(n3239), .I1(n3263), .CO(n28526));
    SB_LUT4 rem_4_add_2189_21_lut (.I0(n3240), .I1(n3240), .I2(n3263), 
            .I3(n28524), .O(n3339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_21 (.CI(n28524), .I0(n3240), .I1(n3263), .CO(n28525));
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n27887), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_20_lut (.I0(n3241), .I1(n3241), .I2(n3263), 
            .I3(n28523), .O(n3340)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_20 (.CI(n28523), .I0(n3241), .I1(n3263), .CO(n28524));
    SB_LUT4 i13222_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17951));   // verilog/coms.v(126[12] 292[6])
    defparam i13222_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1586_9 (.CI(n28847), .I0(n2352), .I1(VCC_net), 
            .CO(n28848));
    SB_LUT4 rem_4_add_2189_19_lut (.I0(n3242), .I1(n3242), .I2(n3263), 
            .I3(n28522), .O(n3341)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n28846), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13221_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17950));   // verilog/coms.v(126[12] 292[6])
    defparam i13221_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_19 (.CI(n28522), .I0(n3242), .I1(n3263), .CO(n28523));
    SB_LUT4 div_46_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4993));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2189_18_lut (.I0(n3243), .I1(n3243), .I2(n3263), 
            .I3(n28521), .O(n3342)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1586_8 (.CI(n28846), .I0(n2353), .I1(VCC_net), 
            .CO(n28847));
    SB_CARRY rem_4_add_2189_18 (.CI(n28521), .I0(n3243), .I1(n3263), .CO(n28522));
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n28845), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_17_lut (.I0(n3244), .I1(n3244), .I2(n3263), 
            .I3(n28520), .O(n3343)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13224_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17953));   // verilog/coms.v(126[12] 292[6])
    defparam i13224_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_17 (.CI(n28520), .I0(n3244), .I1(n3263), .CO(n28521));
    SB_LUT4 rem_4_add_2189_16_lut (.I0(n3245), .I1(n3245), .I2(n3263), 
            .I3(n28519), .O(n3344)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_16 (.CI(n28519), .I0(n3245), .I1(n3263), .CO(n28520));
    SB_LUT4 rem_4_add_2189_15_lut (.I0(n3246), .I1(n3246), .I2(n3263), 
            .I3(n28518), .O(n3345)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_983_9 (.CI(n27887), .I0(n1451), .I1(VCC_net), .CO(n27888));
    SB_CARRY rem_4_add_1586_7 (.CI(n28845), .I0(n2354), .I1(GND_net), 
            .CO(n28846));
    SB_CARRY rem_4_add_2189_15 (.CI(n28518), .I0(n3246), .I1(n3263), .CO(n28519));
    SB_LUT4 rem_4_add_2189_14_lut (.I0(n3247), .I1(n3247), .I2(n3263), 
            .I3(n28517), .O(n3346)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_14 (.CI(n28517), .I0(n3247), .I1(n3263), .CO(n28518));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(n3248), .I1(n3248), .I2(n3263), 
            .I3(n28516), .O(n3347)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_i1657_3_lut_3_lut (.I0(n2471), .I1(n6110), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_13 (.CI(n28516), .I0(n3248), .I1(n3263), .CO(n28517));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(n3249), .I1(n3249), .I2(n3263), 
            .I3(n28515), .O(n3348)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_i1337_3_lut_3_lut (.I0(n1991), .I1(n6010), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n28844), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_12 (.CI(n28515), .I0(n3249), .I1(n3263), .CO(n28516));
    SB_LUT4 i13223_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17952));   // verilog/coms.v(126[12] 292[6])
    defparam i13223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_11_lut (.I0(n3250), .I1(n3250), .I2(n3263), 
            .I3(n28514), .O(n3349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_11 (.CI(n28514), .I0(n3250), .I1(n3263), .CO(n28515));
    SB_LUT4 rem_4_add_2189_10_lut (.I0(n3251), .I1(n3251), .I2(n3263), 
            .I3(n28513), .O(n3350)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13226_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17955));   // verilog/coms.v(126[12] 292[6])
    defparam i13226_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1586_6 (.CI(n28844), .I0(n2355), .I1(GND_net), 
            .CO(n28845));
    SB_CARRY rem_4_add_2189_10 (.CI(n28513), .I0(n3251), .I1(n3263), .CO(n28514));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n27886), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n28843), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_9_lut (.I0(n3252), .I1(n3252), .I2(n3263), 
            .I3(n28512), .O(n3351)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1586_5 (.CI(n28843), .I0(n2356), .I1(VCC_net), 
            .CO(n28844));
    SB_CARRY rem_4_add_2189_9 (.CI(n28512), .I0(n3252), .I1(n3263), .CO(n28513));
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4954), .I2(VCC_net), 
            .I3(n28842), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_8_lut (.I0(n3253), .I1(n3253), .I2(n3263), 
            .I3(n28511), .O(n3352)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_983_8 (.CI(n27886), .I0(n1452), .I1(VCC_net), .CO(n27887));
    SB_CARRY rem_4_add_2189_8 (.CI(n28511), .I0(n3253), .I1(n3263), .CO(n28512));
    SB_LUT4 div_46_i1653_3_lut_3_lut (.I0(n2471), .I1(n6106), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_7_lut (.I0(n3254), .I1(n3254), .I2(n43147), 
            .I3(n28510), .O(n3353)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_2189_7 (.CI(n28510), .I0(n3254), .I1(n43147), .CO(n28511));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(n3255), .I1(n3255), .I2(n43147), 
            .I3(n28509), .O(n3354)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_2189_6 (.CI(n28509), .I0(n3255), .I1(n43147), .CO(n28510));
    SB_CARRY rem_4_add_1586_4 (.CI(n28842), .I0(n2357_adj_4954), .I1(VCC_net), 
            .CO(n28843));
    SB_LUT4 i13225_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17954));   // verilog/coms.v(126[12] 292[6])
    defparam i13225_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_5_lut (.I0(n3256), .I1(n3256), .I2(n3263), 
            .I3(n28508), .O(n3355)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4985));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4988));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2189_5 (.CI(n28508), .I0(n3256), .I1(n3263), .CO(n28509));
    SB_LUT4 div_46_i1652_3_lut_3_lut (.I0(n2471), .I1(n6105), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_4_lut (.I0(n3257), .I1(n3257), .I2(n3263), 
            .I3(n28507), .O(n3356)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_2189_4 (.CI(n28507), .I0(n3257), .I1(n3263), .CO(n28508));
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4953), .I2(GND_net), 
            .I3(n28841), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_3 (.CI(n28841), .I0(n2358_adj_4953), .I1(GND_net), 
            .CO(n28842));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(n3258), .I1(n3258), .I2(n43147), 
            .I3(n28506), .O(n3357)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_2189_3 (.CI(n28506), .I0(n3258), .I1(n43147), .CO(n28507));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4938), .I1(VCC_net), 
            .CO(n28841));
    SB_LUT4 rem_4_add_1653_23_lut (.I0(n2471_adj_4937), .I1(n2438), .I2(VCC_net), 
            .I3(n28840), .O(n2537_adj_4887)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(GND_net), .I1(n2439), .I2(VCC_net), 
            .I3(n28839), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n27885), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_22 (.CI(n28839), .I0(n2439), .I1(VCC_net), 
            .CO(n28840));
    SB_LUT4 rem_4_add_1653_21_lut (.I0(GND_net), .I1(n2440), .I2(VCC_net), 
            .I3(n28838), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_21 (.CI(n28838), .I0(n2440), .I1(VCC_net), 
            .CO(n28839));
    SB_LUT4 rem_4_add_1653_20_lut (.I0(GND_net), .I1(n2441), .I2(VCC_net), 
            .I3(n28837), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3358), .I1(VCC_net), 
            .CO(n28506));
    SB_CARRY rem_4_add_1653_20 (.CI(n28837), .I0(n2441), .I1(VCC_net), 
            .CO(n28838));
    SB_LUT4 rem_4_add_1653_19_lut (.I0(GND_net), .I1(n2442), .I2(VCC_net), 
            .I3(n28836), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_7 (.CI(n27885), .I0(n1453), .I1(VCC_net), .CO(n27886));
    SB_CARRY rem_4_add_1653_19 (.CI(n28836), .I0(n2442), .I1(VCC_net), 
            .CO(n28837));
    SB_LUT4 rem_4_add_1653_18_lut (.I0(GND_net), .I1(n2443), .I2(VCC_net), 
            .I3(n28835), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n27884), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1185_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n28505), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1185_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n28504), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_18 (.CI(n28835), .I0(n2443), .I1(VCC_net), 
            .CO(n28836));
    SB_LUT4 div_46_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4987));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1185_add_4_32 (.CI(n28504), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n28505));
    SB_LUT4 div_46_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4992));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_1185_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n28503), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_31 (.CI(n28503), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n28504));
    SB_CARRY rem_4_add_983_6 (.CI(n27884), .I0(n1454), .I1(GND_net), .CO(n27885));
    SB_LUT4 rem_4_add_1653_17_lut (.I0(GND_net), .I1(n2444), .I2(VCC_net), 
            .I3(n28834), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n27883), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1185_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n28502), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_17 (.CI(n28834), .I0(n2444), .I1(VCC_net), 
            .CO(n28835));
    SB_LUT4 rem_4_add_1653_16_lut (.I0(GND_net), .I1(n2445), .I2(VCC_net), 
            .I3(n28833), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1660_3_lut_3_lut (.I0(n2471), .I1(n6113), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_30 (.CI(n28502), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n28503));
    SB_LUT4 div_46_i1601_3_lut_3_lut (.I0(n2381), .I1(n6092), .I2(n665), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1185_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n28501), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_29 (.CI(n28501), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n28502));
    SB_LUT4 communication_counter_1185_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n28500), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1659_3_lut_3_lut (.I0(n2471), .I1(n6112), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_28 (.CI(n28500), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n28501));
    SB_LUT4 communication_counter_1185_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n28499), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13230_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17959));   // verilog/coms.v(126[12] 292[6])
    defparam i13230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13229_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17958));   // verilog/coms.v(126[12] 292[6])
    defparam i13229_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13228_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17957));   // verilog/coms.v(126[12] 292[6])
    defparam i13228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13227_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17956));   // verilog/coms.v(126[12] 292[6])
    defparam i13227_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4895));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1398_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34861_3_lut (.I0(n1953), .I1(n2020), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13241_3_lut (.I0(encoder0_position[5]), .I1(n3013), .I2(count_enable), 
            .I3(GND_net), .O(n17970));   // quad.v(35[10] 41[6])
    defparam i13241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13240_3_lut (.I0(encoder0_position[4]), .I1(n3014), .I2(count_enable), 
            .I3(GND_net), .O(n17969));   // quad.v(35[10] 41[6])
    defparam i13240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13239_3_lut (.I0(encoder0_position[3]), .I1(n3015), .I2(count_enable), 
            .I3(GND_net), .O(n17968));   // quad.v(35[10] 41[6])
    defparam i13239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13238_3_lut (.I0(encoder0_position[2]), .I1(n3016), .I2(count_enable), 
            .I3(GND_net), .O(n17967));   // quad.v(35[10] 41[6])
    defparam i13238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13237_3_lut (.I0(encoder0_position[1]), .I1(n3017), .I2(count_enable), 
            .I3(GND_net), .O(n17966));   // quad.v(35[10] 41[6])
    defparam i13237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13236_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17965));   // verilog/coms.v(126[12] 292[6])
    defparam i13236_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1185_add_4_27 (.CI(n28499), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n28500));
    SB_LUT4 i13235_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17964));   // verilog/coms.v(126[12] 292[6])
    defparam i13235_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13234_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17963));   // verilog/coms.v(126[12] 292[6])
    defparam i13234_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13233_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17962));   // verilog/coms.v(126[12] 292[6])
    defparam i13233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13332_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1172), .I3(GND_net), .O(n18061));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4983));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13245_3_lut (.I0(encoder0_position[9]), .I1(n3009), .I2(count_enable), 
            .I3(GND_net), .O(n17974));   // quad.v(35[10] 41[6])
    defparam i13245_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_983_5 (.CI(n27883), .I0(n1455), .I1(GND_net), .CO(n27884));
    SB_LUT4 i13244_3_lut (.I0(encoder0_position[8]), .I1(n3010), .I2(count_enable), 
            .I3(GND_net), .O(n17973));   // quad.v(35[10] 41[6])
    defparam i13244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1658_3_lut_3_lut (.I0(n2471), .I1(n6111), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13243_3_lut (.I0(encoder0_position[7]), .I1(n3011), .I2(count_enable), 
            .I3(GND_net), .O(n17972));   // quad.v(35[10] 41[6])
    defparam i13243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1185_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n28498), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13242_3_lut (.I0(encoder0_position[6]), .I1(n3012), .I2(count_enable), 
            .I3(GND_net), .O(n17971));   // quad.v(35[10] 41[6])
    defparam i13242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13253_3_lut (.I0(encoder0_position[17]), .I1(n3001), .I2(count_enable), 
            .I3(GND_net), .O(n17982));   // quad.v(35[10] 41[6])
    defparam i13253_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_16 (.CI(n28833), .I0(n2445), .I1(VCC_net), 
            .CO(n28834));
    SB_LUT4 i34163_4_lut (.I0(n37_adj_4988), .I1(n35_adj_4987), .I2(n33_adj_4985), 
            .I3(n31_adj_4983), .O(n40995));
    defparam i34163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_985_i42_3_lut (.I0(n34_adj_4986), .I1(n91), 
            .I2(n45_adj_4993), .I3(GND_net), .O(n42_adj_4991));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_985_i30_4_lut (.I0(n657), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4982));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35059_3_lut (.I0(n30_adj_4982), .I1(n95), .I2(n37_adj_4988), 
            .I3(GND_net), .O(n41891));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35059_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35060_3_lut (.I0(n41891), .I1(n94), .I2(n39_adj_4989), .I3(GND_net), 
            .O(n41892));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35060_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY communication_counter_1185_add_4_26 (.CI(n28498), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n28499));
    SB_LUT4 i13252_3_lut (.I0(encoder0_position[16]), .I1(n3002), .I2(count_enable), 
            .I3(GND_net), .O(n17981));   // quad.v(35[10] 41[6])
    defparam i13252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13263_3_lut (.I0(encoder1_position[3]), .I1(n2965), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17992));   // quad.v(35[10] 41[6])
    defparam i13263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34133_4_lut (.I0(n43_adj_4992), .I1(n41_adj_4990), .I2(n39_adj_4989), 
            .I3(n40995), .O(n40965));
    defparam i34133_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13262_3_lut (.I0(encoder1_position[2]), .I1(n2966), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17991));   // quad.v(35[10] 41[6])
    defparam i13262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1185_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n28497), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13261_3_lut (.I0(encoder1_position[1]), .I1(n2967), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17990));   // quad.v(35[10] 41[6])
    defparam i13261_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1185_add_4_25 (.CI(n28497), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n28498));
    SB_LUT4 div_46_i1341_3_lut_3_lut (.I0(n1991), .I1(n6014), .I2(n661), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1656_3_lut_3_lut (.I0(n2471), .I1(n6109), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35099_4_lut (.I0(n42_adj_4991), .I1(n32_adj_4984), .I2(n45_adj_4993), 
            .I3(n40960), .O(n41931));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35099_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34382_3_lut (.I0(n41892), .I1(n93), .I2(n41_adj_4990), .I3(GND_net), 
            .O(n41214));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34382_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35437_4_lut (.I0(n41214), .I1(n41931), .I2(n45_adj_4993), 
            .I3(n40965), .O(n42269));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35437_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n42269), .I1(n15854), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1333_3_lut_3_lut (.I0(n1991), .I1(n6006), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1649_3_lut_3_lut (.I0(n2471), .I1(n6102), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1185_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n28496), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4981));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i37_2_lut (.I0(n1417_adj_4752), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4978));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1654_3_lut_3_lut (.I0(n2471), .I1(n6107), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13265_3_lut (.I0(encoder1_position[5]), .I1(n2963), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17994));   // quad.v(35[10] 41[6])
    defparam i13265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13264_3_lut (.I0(encoder1_position[4]), .I1(n2964), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17993));   // quad.v(35[10] 41[6])
    defparam i13264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4980));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13267_3_lut (.I0(encoder1_position[7]), .I1(n2961), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17996));   // quad.v(35[10] 41[6])
    defparam i13267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1332_3_lut_3_lut (.I0(n1991), .I1(n6005), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1713_3_lut_3_lut (.I0(n2558), .I1(n6131), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1699_3_lut_3_lut (.I0(n2558), .I1(n6117), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_24 (.CI(n28496), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n28497));
    SB_LUT4 communication_counter_1185_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n28495), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13266_3_lut (.I0(encoder1_position[6]), .I1(n2962), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17995));   // quad.v(35[10] 41[6])
    defparam i13266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13269_3_lut (.I0(encoder1_position[9]), .I1(n2959), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17998));   // quad.v(35[10] 41[6])
    defparam i13269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4979));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1700_3_lut_3_lut (.I0(n2558), .I1(n6118), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1653_15_lut (.I0(GND_net), .I1(n2446), .I2(VCC_net), 
            .I3(n28832), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_23 (.CI(n28495), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n28496));
    SB_LUT4 communication_counter_1185_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n28494), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4725), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n656));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13268_3_lut (.I0(encoder1_position[8]), .I1(n2960), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17997));   // quad.v(35[10] 41[6])
    defparam i13268_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1185_add_4_22 (.CI(n28494), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n28495));
    SB_LUT4 div_46_i1701_3_lut_3_lut (.I0(n2558), .I1(n6119), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1404_3_lut_3_lut (.I0(n2093), .I1(n6027), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1653_15 (.CI(n28832), .I0(n2446), .I1(VCC_net), 
            .CO(n28833));
    SB_LUT4 communication_counter_1185_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n28493), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1702_3_lut_3_lut (.I0(n2558), .I1(n6120), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1705_3_lut_3_lut (.I0(n2558), .I1(n6123), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_21 (.CI(n28493), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n28494));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(GND_net), .I1(n2447_adj_4949), .I2(VCC_net), 
            .I3(n28831), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1185_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n28492), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13271_3_lut (.I0(encoder1_position[11]), .I1(n2957), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18000));   // quad.v(35[10] 41[6])
    defparam i13271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13270_3_lut (.I0(encoder1_position[10]), .I1(n2958), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17999));   // quad.v(35[10] 41[6])
    defparam i13270_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1185_add_4_20 (.CI(n28492), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n28493));
    SB_LUT4 i13273_3_lut (.I0(encoder1_position[13]), .I1(n2955), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18002));   // quad.v(35[10] 41[6])
    defparam i13273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1185_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n28491), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1703_3_lut_3_lut (.I0(n2558), .I1(n6121), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13272_3_lut (.I0(encoder1_position[12]), .I1(n2956), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18001));   // quad.v(35[10] 41[6])
    defparam i13272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1706_3_lut_3_lut (.I0(n2558), .I1(n6124), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1719_3_lut_3_lut (.I0(n2558), .I1(n6137), .I2(n667), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_906_i32_4_lut (.I0(n656), .I1(n99), .I2(n1420_adj_4755), 
            .I3(n558), .O(n32_adj_4976));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_1653_14 (.CI(n28831), .I0(n2447_adj_4949), .I1(VCC_net), 
            .CO(n28832));
    SB_LUT4 i35234_3_lut (.I0(n32_adj_4976), .I1(n95), .I2(n39_adj_4979), 
            .I3(GND_net), .O(n42066));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35234_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34862_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1704_3_lut_3_lut (.I0(n2558), .I1(n6122), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35235_3_lut (.I0(n42066), .I1(n94), .I2(n41_adj_4980), .I3(GND_net), 
            .O(n42067));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35235_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1708_3_lut_3_lut (.I0(n2558), .I1(n6126), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34181_4_lut (.I0(n41_adj_4980), .I1(n39_adj_4979), .I2(n37_adj_4978), 
            .I3(n40316), .O(n41013));
    defparam i34181_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34833_3_lut (.I0(n34_adj_4977), .I1(n96), .I2(n37_adj_4978), 
            .I3(GND_net), .O(n41665));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34833_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35096_3_lut (.I0(n42067), .I1(n93), .I2(n43_adj_4981), .I3(GND_net), 
            .O(n41928));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35096_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35232_4_lut (.I0(n41928), .I1(n41665), .I2(n43_adj_4981), 
            .I3(n41013), .O(n42064));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35232_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35233_3_lut (.I0(n42064), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n42065));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35233_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY communication_counter_1185_add_4_19 (.CI(n28491), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n28492));
    SB_LUT4 rem_4_add_1653_13_lut (.I0(GND_net), .I1(n2448_adj_4948), .I2(VCC_net), 
            .I3(n28830), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n27882), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1185_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n28490), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n42065), .I1(n15801), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hceef;
    SB_CARRY communication_counter_1185_add_4_18 (.CI(n28490), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n28491));
    SB_LUT4 communication_counter_1185_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n28489), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_17 (.CI(n28489), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n28490));
    SB_LUT4 communication_counter_1185_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n28488), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1709_3_lut_3_lut (.I0(n2558), .I1(n6127), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1399_3_lut_3_lut (.I0(n2093), .I1(n6022), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4970));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1185_add_4_16 (.CI(n28488), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n28489));
    SB_LUT4 i13213_3_lut (.I0(\data_in_frame[24] [7]), .I1(rx_data[7]), 
            .I2(n36887), .I3(GND_net), .O(n17942));   // verilog/coms.v(126[12] 292[6])
    defparam i13213_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 div_46_i1710_3_lut_3_lut (.I0(n2558), .I1(n6128), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 div_46_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4972));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 div_46_i1711_3_lut_3_lut (.I0(n2558), .I1(n6129), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 i15_4_lut (.I0(n2752), .I1(n2748), .I2(n2753), .I3(n2749), 
            .O(n35));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 div_46_i1715_3_lut_3_lut (.I0(n2558), .I1(n6133), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 i13212_3_lut (.I0(\data_in_frame[24] [6]), .I1(rx_data[6]), 
            .I2(n36887), .I3(GND_net), .O(n17941));   // verilog/coms.v(126[12] 292[6])
    defparam i13212_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 div_46_i1401_3_lut_3_lut (.I0(n2093), .I1(n6024), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 i13211_3_lut (.I0(\data_in_frame[24] [5]), .I1(rx_data[5]), 
            .I2(n36887), .I3(GND_net), .O(n17940));   // verilog/coms.v(126[12] 292[6])
    defparam i13211_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 div_46_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4974));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13210_3_lut (.I0(\data_in_frame[24] [4]), .I1(rx_data[4]), 
            .I2(n36887), .I3(GND_net), .O(n17939));   // verilog/coms.v(126[12] 292[6])
    defparam i13210_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 div_46_i1716_3_lut_3_lut (.I0(n2558), .I1(n6134), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 communication_counter_1185_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n28487), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF communication_counter_1185__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_LUT4 rem_4_i1396_3_lut (.I0(n2051), .I1(n2118), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2150));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1395_3_lut (.I0(n2050), .I1(n2117), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1185_add_4_15 (.CI(n28487), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n28488));
    SB_LUT4 i1_3_lut_adj_1742 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n35620));
    defparam i1_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut (.I0(n2046), .I1(n2054), .I2(n35620), .I3(n2055), 
            .O(n16_adj_5340));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i9_4_lut (.I0(n2047), .I1(n2053), .I2(n2048), .I3(n2051), 
            .O(n22_adj_5338));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n2050), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_5339));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1743 (.I0(n2044), .I1(n22_adj_5338), .I2(n16_adj_5340), 
            .I3(n2045), .O(n24_adj_5337));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1744 (.I0(n2049), .I1(n24_adj_5337), .I2(n20_adj_5339), 
            .I3(n2052), .O(n2075_adj_4994));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1745 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n35578));
    defparam i1_3_lut_adj_1745.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1746 (.I0(n2154), .I1(n2147), .I2(n35578), .I3(n2155), 
            .O(n18_adj_4761));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1746.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut_adj_1747 (.I0(n2148), .I1(n2149), .I2(n2150), .I3(n2151), 
            .O(n24_adj_4756));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_4757));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1748 (.I0(n2145), .I1(n24_adj_4756), .I2(n18_adj_4761), 
            .I3(n2146), .O(n26));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_1185_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n28486), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1749 (.I0(n2153), .I1(n26), .I2(n22_adj_4757), 
            .I3(n2152), .O(n2174_adj_4975));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4775), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4894));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4971));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i2015_3_lut (.I0(n2958_adj_4802), .I1(n3025), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1712_3_lut_3_lut (.I0(n2558), .I1(n6130), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2014_3_lut (.I0(n2957_adj_4803), .I1(n3024), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1718_3_lut_3_lut (.I0(n2558), .I1(n6136), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13209_3_lut (.I0(\data_in_frame[24] [3]), .I1(rx_data[3]), 
            .I2(n36887), .I3(GND_net), .O(n17938));   // verilog/coms.v(126[12] 292[6])
    defparam i13209_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1185_add_4_14 (.CI(n28486), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n28487));
    SB_LUT4 div_46_i1397_3_lut_3_lut (.I0(n2093), .I1(n6020), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13208_3_lut (.I0(\data_in_frame[24] [2]), .I1(rx_data[2]), 
            .I2(n36887), .I3(GND_net), .O(n17937));   // verilog/coms.v(126[12] 292[6])
    defparam i13208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1717_3_lut_3_lut (.I0(n2558), .I1(n6135), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1714_3_lut_3_lut (.I0(n2558), .I1(n6132), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1653_13 (.CI(n28830), .I0(n2448_adj_4948), .I1(VCC_net), 
            .CO(n28831));
    SB_LUT4 i13207_3_lut (.I0(\data_in_frame[24] [1]), .I1(rx_data[1]), 
            .I2(n36887), .I3(GND_net), .O(n17936));   // verilog/coms.v(126[12] 292[6])
    defparam i13207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4776), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2013_3_lut (.I0(n2956_adj_4804), .I1(n3023), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4893));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4892));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1653_12_lut (.I0(GND_net), .I1(n2449_adj_4947), .I2(VCC_net), 
            .I3(n28829), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4891));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22_3_lut_adj_1750 (.I0(bit_ctr[3]), .I1(n40244), .I2(n4442), 
            .I3(GND_net), .O(n33477));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1750.LUT_INIT = 16'hacac;
    SB_LUT4 i13334_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1172), .I3(GND_net), .O(n18063));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1334_3_lut (.I0(n1957), .I1(n2024), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2012_3_lut (.I0(n2955_adj_4805), .I1(n3022), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4890));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2011_3_lut (.I0(n2954_adj_4806), .I1(n3021), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4889));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2010_3_lut (.I0(n2953_adj_4807), .I1(n3020), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3052));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2009_3_lut (.I0(n2952_adj_4808), .I1(n3019), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3051));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1707_3_lut_3_lut (.I0(n2558), .I1(n6125), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n655));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13283_3_lut (.I0(encoder1_position[23]), .I1(n2945), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18012));   // quad.v(35[10] 41[6])
    defparam i13283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13282_3_lut (.I0(encoder1_position[22]), .I1(n2946), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18011));   // quad.v(35[10] 41[6])
    defparam i13282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1769_3_lut_3_lut (.I0(n2642), .I1(n6155), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1754_3_lut_3_lut (.I0(n2642), .I1(n6140), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4936));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2008_3_lut (.I0(n2951_adj_4809), .I1(n3018_adj_4762), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3050));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2007_3_lut (.I0(n2950_adj_4810), .I1(n3017_adj_4763), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3049));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2006_3_lut (.I0(n2949_adj_4811), .I1(n3016_adj_4764), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3048));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4935));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2005_3_lut (.I0(n2948_adj_4812), .I1(n3015_adj_4671), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3047));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2004_3_lut (.I0(n2947_adj_4813), .I1(n3014_adj_4783), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3046));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4934));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4933));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1329_3_lut (.I0(n1952), .I1(n2019), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2003_3_lut (.I0(n2946_adj_4814), .I1(n3013_adj_4784), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3045));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4932));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1328_3_lut (.I0(n1951), .I1(n2018), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4931));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4930));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1327_3_lut (.I0(n1950), .I1(n2017), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_12 (.CI(n28829), .I0(n2449_adj_4947), .I1(VCC_net), 
            .CO(n28830));
    SB_CARRY rem_4_add_983_4 (.CI(n27882), .I0(n1456), .I1(VCC_net), .CO(n27883));
    SB_LUT4 communication_counter_1185_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n28485), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_11_lut (.I0(GND_net), .I1(n2450_adj_4946), .I2(VCC_net), 
            .I3(n28828), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1755_3_lut_3_lut (.I0(n2642), .I1(n6141), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13281_3_lut (.I0(encoder1_position[21]), .I1(n2947), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18010));   // quad.v(35[10] 41[6])
    defparam i13281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13280_3_lut (.I0(encoder1_position[20]), .I1(n2948), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18009));   // quad.v(35[10] 41[6])
    defparam i13280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13279_3_lut (.I0(encoder1_position[19]), .I1(n2949), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18008));   // quad.v(35[10] 41[6])
    defparam i13279_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1185_add_4_13 (.CI(n28485), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n28486));
    SB_LUT4 i13278_3_lut (.I0(encoder1_position[18]), .I1(n2950), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18007));   // quad.v(35[10] 41[6])
    defparam i13278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_825_i34_4_lut (.I0(n655), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34_adj_4967));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_i1756_3_lut_3_lut (.I0(n2642), .I1(n6142), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35236_3_lut (.I0(n34_adj_4967), .I1(n95), .I2(n41_adj_4971), 
            .I3(GND_net), .O(n42068));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35236_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35237_3_lut (.I0(n42068), .I1(n94), .I2(n43_adj_4972), .I3(GND_net), 
            .O(n42069));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35237_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13277_3_lut (.I0(encoder1_position[17]), .I1(n2951), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18006));   // quad.v(35[10] 41[6])
    defparam i13277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n27881), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1185_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n28484), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_12 (.CI(n28484), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n28485));
    SB_LUT4 i34203_4_lut (.I0(n43_adj_4972), .I1(n41_adj_4971), .I2(n39_adj_4970), 
            .I3(n40330), .O(n41035));
    defparam i34203_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_825_i38_3_lut (.I0(n36_adj_4968), .I1(n96), 
            .I2(n39_adj_4970), .I3(GND_net), .O(n38_adj_4969));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13276_3_lut (.I0(encoder1_position[16]), .I1(n2952), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18005));   // quad.v(35[10] 41[6])
    defparam i13276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1757_3_lut_3_lut (.I0(n2642), .I1(n6143), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35094_3_lut (.I0(n42069), .I1(n93), .I2(n45_adj_4974), .I3(GND_net), 
            .O(n44_adj_4973));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35094_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34831_4_lut (.I0(n44_adj_4973), .I1(n38_adj_4969), .I2(n45_adj_4974), 
            .I3(n41035), .O(n41663));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34831_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n41663), .I1(n15797), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'hceef;
    SB_LUT4 i36279_4_lut (.I0(r_SM_Main[2]), .I1(n40217), .I2(n40218), 
            .I3(r_SM_Main[1]), .O(n24450));
    defparam i36279_4_lut.LUT_INIT = 16'h0511;
    SB_CARRY rem_4_add_1653_11 (.CI(n28828), .I0(n2450_adj_4946), .I1(VCC_net), 
            .CO(n28829));
    SB_LUT4 div_46_LessThan_742_i41_2_lut (.I0(n1172_adj_4751), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4966));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1653_10_lut (.I0(GND_net), .I1(n2451_adj_4945), .I2(VCC_net), 
            .I3(n28827), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13291_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n35976), 
            .I3(GND_net), .O(n18020));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13291_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_1185_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n28483), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_11 (.CI(n28483), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n28484));
    SB_LUT4 div_46_i1758_3_lut_3_lut (.I0(n2642), .I1(n6144), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4718), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n654));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1761_3_lut_3_lut (.I0(n2642), .I1(n6147), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut_adj_1752 (.I0(n2742), .I1(n2743), .I2(n2747), .I3(n2750), 
            .O(n33_adj_4801));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1752.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_1185_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n28482), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_742_i36_4_lut (.I0(n654), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36_adj_4963));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_742_i40_3_lut (.I0(n38_adj_4964), .I1(n96), 
            .I2(n41_adj_4966), .I3(GND_net), .O(n40_adj_4965));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13302_3_lut (.I0(color[4]), .I1(n17111), .I2(n15_adj_4714), 
            .I3(GND_net), .O(n18031));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i13302_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35435_4_lut (.I0(n40_adj_4965), .I1(n36_adj_4963), .I2(n41_adj_4966), 
            .I3(n40390), .O(n42267));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35435_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13301_3_lut (.I0(color[3]), .I1(n17111), .I2(n15_adj_4714), 
            .I3(GND_net), .O(n18030));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i13301_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35436_3_lut (.I0(n42267), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n42268));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35436_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13300_3_lut (.I0(color[2]), .I1(n17111), .I2(n15_adj_4714), 
            .I3(GND_net), .O(n18029));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i13300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1762_3_lut_3_lut (.I0(n2642), .I1(n6148), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35354_3_lut (.I0(n42268), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n42186));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35354_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i19_4_lut_adj_1753 (.I0(n33_adj_4801), .I1(n35), .I2(n34_adj_4800), 
            .I3(n36_adj_4799), .O(n2768));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n42186), .I1(n15851), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823), .I2(n2768), .I3(GND_net), 
            .O(n2855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13232_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17961));   // verilog/coms.v(126[12] 292[6])
    defparam i13232_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1185_add_4_10 (.CI(n28482), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n28483));
    SB_CARRY rem_4_add_1653_10 (.CI(n28827), .I0(n2451_adj_4945), .I1(VCC_net), 
            .CO(n28828));
    SB_LUT4 div_46_i1759_3_lut_3_lut (.I0(n2642), .I1(n6145), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1760_3_lut_3_lut (.I0(n2642), .I1(n6146), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1185_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n28481), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_3 (.CI(n27881), .I0(n1457), .I1(VCC_net), .CO(n27882));
    SB_LUT4 rem_4_add_1653_9_lut (.I0(GND_net), .I1(n2452_adj_4944), .I2(VCC_net), 
            .I3(n28826), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_9 (.CI(n28826), .I0(n2452_adj_4944), .I1(VCC_net), 
            .CO(n28827));
    SB_LUT4 rem_4_add_1653_8_lut (.I0(GND_net), .I1(n2453_adj_4943), .I2(VCC_net), 
            .I3(n28825), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4961));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1775_3_lut_3_lut (.I0(n2642), .I1(n6161), .I2(n668), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1764_3_lut_3_lut (.I0(n2642), .I1(n6150), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_9 (.CI(n28481), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n28482));
    SB_LUT4 div_46_i1396_3_lut_3_lut (.I0(n2093), .I1(n6019), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4719), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n653));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_8 (.CI(n28825), .I0(n2453_adj_4943), .I1(VCC_net), 
            .CO(n28826));
    SB_LUT4 rem_4_add_983_2_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(VCC_net), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13231_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17960));   // verilog/coms.v(126[12] 292[6])
    defparam i13231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1395_3_lut_3_lut (.I0(n2093), .I1(n6018), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1185_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n28480), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1765_3_lut_3_lut (.I0(n2642), .I1(n6151), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1766_3_lut_3_lut (.I0(n2642), .I1(n6152), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_8 (.CI(n28480), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n28481));
    SB_LUT4 div_46_i1767_3_lut_3_lut (.I0(n2642), .I1(n6153), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1185_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n28479), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_7 (.CI(n28479), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n28480));
    SB_LUT4 communication_counter_1185_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n28478), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27_3_lut (.I0(n1166), .I1(n35327), .I2(state[0]), .I3(GND_net), 
            .O(n19_adj_5255));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4929));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2002_3_lut (.I0(n2945_adj_4815), .I1(n3012_adj_4785), 
            .I2(n2966_adj_4798), .I3(GND_net), .O(n3044));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2001_3_lut (.I0(n2944), .I1(n3011_adj_4786), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3043));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1773_3_lut_3_lut (.I0(n2642), .I1(n6159), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_657_i38_4_lut (.I0(n653), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4958));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_657_i42_3_lut (.I0(n40_adj_4959), .I1(n96), 
            .I2(n43_adj_4961), .I3(GND_net), .O(n42_adj_4960));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY communication_counter_1185_add_4_6 (.CI(n28478), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n28479));
    SB_LUT4 i24_3_lut_adj_1755 (.I0(n40225), .I1(bit_ctr[8]), .I2(n4442), 
            .I3(GND_net), .O(n33433));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1755.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1756 (.I0(bit_ctr[15]), .I1(n40236), .I2(n4442), 
            .I3(GND_net), .O(n33461));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1756.LUT_INIT = 16'hacac;
    SB_LUT4 i35240_4_lut (.I0(n42_adj_4960), .I1(n38_adj_4958), .I2(n43_adj_4961), 
            .I3(n40401), .O(n42072));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35240_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 communication_counter_1185_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n28477), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1774_3_lut_3_lut (.I0(n2642), .I1(n6160), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1770_3_lut_3_lut (.I0(n2642), .I1(n6156), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_5 (.CI(n28477), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n28478));
    SB_LUT4 div_46_i1771_3_lut_3_lut (.I0(n2642), .I1(n6157), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35241_3_lut (.I0(n42072), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n42073));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35241_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i1772_3_lut_3_lut (.I0(n2642), .I1(n6158), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n42073), .I1(n15794), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'hceef;
    SB_LUT4 communication_counter_1185_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n28476), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13307_3_lut (.I0(quadA_debounced_adj_4699), .I1(reg_B_adj_5390[1]), 
            .I2(n35775), .I3(GND_net), .O(n18036));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13307_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1458), .I1(GND_net), 
            .CO(n27881));
    SB_LUT4 div_46_i1768_3_lut_3_lut (.I0(n2642), .I1(n6154), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1763_3_lut_3_lut (.I0(n2642), .I1(n6149), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1185_add_4_4 (.CI(n28476), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n28477));
    SB_LUT4 i13310_3_lut (.I0(setpoint[2]), .I1(n4351), .I2(n36881), .I3(GND_net), 
            .O(n18039));   // verilog/coms.v(126[12] 292[6])
    defparam i13310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22717_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4688), .I3(GND_net), 
            .O(n8_adj_4687));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22717_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 communication_counter_1185_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n28475), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1185_add_4_3 (.CI(n28475), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n28476));
    SB_LUT4 rem_4_add_1653_7_lut (.I0(GND_net), .I1(n2454_adj_4942), .I2(GND_net), 
            .I3(n28824), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_7 (.CI(n28824), .I0(n2454_adj_4942), .I1(GND_net), 
            .CO(n28825));
    SB_LUT4 communication_counter_1185_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1185_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13309_3_lut (.I0(setpoint[1]), .I1(n4350), .I2(n36881), .I3(GND_net), 
            .O(n18038));   // verilog/coms.v(126[12] 292[6])
    defparam i13309_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1185_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n28475));
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n43086), .I1(n2_adj_5272), .I2(n3452), 
            .I3(n28474), .O(color_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i22709_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4689), .I3(GND_net), 
            .O(n6_adj_4688));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22709_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_i1398_3_lut_3_lut (.I0(n2093), .I1(n6021), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n43090), .I1(n2_adj_5272), .I2(n3453), 
            .I3(n28473), .O(color_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13312_3_lut (.I0(setpoint[4]), .I1(n4353), .I2(n36881), .I3(GND_net), 
            .O(n18041));   // verilog/coms.v(126[12] 292[6])
    defparam i13312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13311_3_lut (.I0(setpoint[3]), .I1(n4352), .I2(n36881), .I3(GND_net), 
            .O(n18040));   // verilog/coms.v(126[12] 292[6])
    defparam i13311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4720), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2298_8 (.CI(n28473), .I0(n2_adj_5272), .I1(n3453), 
            .CO(n28474));
    SB_LUT4 i13251_3_lut (.I0(encoder0_position[15]), .I1(n3003), .I2(count_enable), 
            .I3(GND_net), .O(n17980));   // quad.v(35[10] 41[6])
    defparam i13251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13250_3_lut (.I0(encoder0_position[14]), .I1(n3004), .I2(count_enable), 
            .I3(GND_net), .O(n17979));   // quad.v(35[10] 41[6])
    defparam i13250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13249_3_lut (.I0(encoder0_position[13]), .I1(n3005), .I2(count_enable), 
            .I3(GND_net), .O(n17978));   // quad.v(35[10] 41[6])
    defparam i13249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13248_3_lut (.I0(encoder0_position[12]), .I1(n3006), .I2(count_enable), 
            .I3(GND_net), .O(n17977));   // quad.v(35[10] 41[6])
    defparam i13248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n43093), .I1(n2_adj_5272), .I2(n3454), 
            .I3(n28472), .O(color_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i22693_2_lut (.I0(n651), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5263));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22693_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_2298_7 (.CI(n28472), .I0(n2_adj_5272), .I1(n3454), 
            .CO(n28473));
    SB_LUT4 i13247_3_lut (.I0(encoder0_position[11]), .I1(n3007), .I2(count_enable), 
            .I3(GND_net), .O(n17976));   // quad.v(35[10] 41[6])
    defparam i13247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13246_3_lut (.I0(encoder0_position[10]), .I1(n3008), .I2(count_enable), 
            .I3(GND_net), .O(n17975));   // quad.v(35[10] 41[6])
    defparam i13246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13316_3_lut (.I0(setpoint[8]), .I1(n4357), .I2(n36881), .I3(GND_net), 
            .O(n18045));   // verilog/coms.v(126[12] 292[6])
    defparam i13316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13315_3_lut (.I0(setpoint[7]), .I1(n4356), .I2(n36881), .I3(GND_net), 
            .O(n18044));   // verilog/coms.v(126[12] 292[6])
    defparam i13315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n43096), .I1(n2_adj_5272), .I2(n3455), 
            .I3(n28471), .O(color_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13314_3_lut (.I0(setpoint[6]), .I1(n4355), .I2(n36881), .I3(GND_net), 
            .O(n18043));   // verilog/coms.v(126[12] 292[6])
    defparam i13314_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2298_6 (.CI(n28471), .I0(n2_adj_5272), .I1(n3455), 
            .CO(n28472));
    SB_LUT4 div_46_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n43099), .I1(n2_adj_5272), .I2(n3456), 
            .I3(n28470), .O(color_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13313_3_lut (.I0(setpoint[5]), .I1(n4354), .I2(n36881), .I3(GND_net), 
            .O(n18042));   // verilog/coms.v(126[12] 292[6])
    defparam i13313_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2298_5 (.CI(n28470), .I0(n2_adj_5272), .I1(n3456), 
            .CO(n28471));
    SB_LUT4 div_46_LessThan_570_i40_4_lut (.I0(n652), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4955));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_570_i44_3_lut (.I0(n42_adj_4956), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4957));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n43102), .I1(n2_adj_5272), .I2(n3457), 
            .I3(n28469), .O(color_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i34825_4_lut (.I0(n44_adj_4957), .I1(n40_adj_4955), .I2(n45), 
            .I3(n40409), .O(n41657));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34825_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_2298_4 (.CI(n28469), .I0(n2_adj_5272), .I1(n3457), 
            .CO(n28470));
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n41657), .I1(n15791), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_5272), 
            .I2(n3458), .I3(n28468), .O(color_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_3 (.CI(n28468), .I0(n2_adj_5272), .I1(n3458), 
            .CO(n28469));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_5272), 
            .I2(n3360), .I3(VCC_net), .O(color_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_5272), .I1(n3360), 
            .CO(n28468));
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5531_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n28467), 
            .O(n10194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1394_3_lut_3_lut (.I0(n2093), .I1(n6017), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4928));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(\FRAME_MATCHER.state_31__N_2661 [2]), .I1(n7_adj_4818), 
            .I2(\FRAME_MATCHER.i_31__N_2625 ), .I3(n2957_adj_4678), .O(n6_adj_4679));   // verilog/coms.v(126[12] 292[6])
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfcec;
    SB_LUT4 i3_4_lut_adj_1760 (.I0(\FRAME_MATCHER.i_31__N_2621 ), .I1(n6_adj_4679), 
            .I2(n9001), .I3(n122), .O(n8));   // verilog/coms.v(126[12] 292[6])
    defparam i3_4_lut_adj_1760.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1761 (.I0(\FRAME_MATCHER.state_31__N_2661 [2]), .I1(n8), 
            .I2(n63), .I3(n5_adj_5312), .O(n43329));   // verilog/coms.v(126[12] 292[6])
    defparam i4_4_lut_adj_1761.LUT_INIT = 16'hefcf;
    SB_LUT4 add_5531_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n28466), 
            .O(n10195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22677_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_5306), .I3(GND_net), 
            .O(n6_adj_5305));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22677_3_lut.LUT_INIT = 16'he8e8;
    SB_CARRY add_5531_6 (.CI(n28466), .I0(n3354), .I1(GND_net), .CO(n28467));
    SB_LUT4 add_5531_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n28465), 
            .O(n10196)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22661_2_lut (.I0(n650), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5308));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22661_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_5531_5 (.CI(n28465), .I0(n3355), .I1(GND_net), .CO(n28466));
    SB_LUT4 add_5531_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n28464), 
            .O(n10197)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4715), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n651));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i483_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5531_4 (.CI(n28464), .I0(n3356), .I1(VCC_net), .CO(n28465));
    SB_LUT4 add_5531_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n28463), 
            .O(n10198)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5531_3 (.CI(n28463), .I0(n3357), .I1(VCC_net), .CO(n28464));
    SB_LUT4 div_46_LessThan_481_i42_4_lut (.I0(n651), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4951));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35242_3_lut (.I0(n42_adj_4951), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n42074));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35242_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13259_3_lut (.I0(encoder0_position[23]), .I1(n2995), .I2(count_enable), 
            .I3(GND_net), .O(n17988));   // quad.v(35[10] 41[6])
    defparam i13259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35243_3_lut (.I0(n42074), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n42075));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35243_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n42075), .I1(n15788), .I2(n96), .I3(n35299), 
            .O(n806));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hefce;
    SB_LUT4 i13258_3_lut (.I0(encoder0_position[22]), .I1(n2996), .I2(count_enable), 
            .I3(GND_net), .O(n17987));   // quad.v(35[10] 41[6])
    defparam i13258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22637_2_lut (.I0(n511), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5307));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22637_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_5531_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10199)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5531_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5531_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n28463));
    SB_LUT4 div_46_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4716), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n650));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2314_25_lut (.I0(n249), .I1(n43152), .I2(n248), .I3(n28462), 
            .O(displacement_23__N_229[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1596_3_lut_3_lut (.I0(n2381), .I1(n6087), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_390_i44_4_lut (.I0(n650), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44_adj_4950));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34821_3_lut (.I0(n44_adj_4950), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n41653));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34821_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n41653), .I1(n15785), .I2(n97), .I3(n35295), 
            .O(n671));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hefce;
    SB_LUT4 i22613_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22613_2_lut.LUT_INIT = 16'heeee;
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4717), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_297_i46_4_lut (.I0(n511), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n46), .I1(n15774), .I2(n98), .I3(n35278), 
            .O(n533));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hefce;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n224), .I1(n99), .I2(n15845), .I3(n558), 
            .O(n5_adj_5257));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'h555d;
    SB_LUT4 div_46_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4702), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33684_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n40177));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33684_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n40177), .I1(n15845), .I2(n99), .I3(n5_adj_5257), 
            .O(n392));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n15817));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1767 (.I0(n81), .I1(n15866), .I2(GND_net), .I3(GND_net), 
            .O(n15883));
    defparam i1_2_lut_adj_1767.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_2314_24_lut (.I0(n393), .I1(n43152), .I2(n392), .I3(n28461), 
            .O(displacement_23__N_229[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1768 (.I0(n84), .I1(n15812), .I2(GND_net), .I3(GND_net), 
            .O(n15863));
    defparam i1_2_lut_adj_1768.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4927));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1260_rep_43_3_lut (.I0(n1851), .I1(n1918), .I2(n1877), 
            .I3(GND_net), .O(n1950));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1260_rep_43_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1259_3_lut (.I0(n1850), .I1(n1917), .I2(n1877), .I3(GND_net), 
            .O(n1949));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1258_3_lut (.I0(n1849), .I1(n1916), .I2(n1877), .I3(GND_net), 
            .O(n1948));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1263_3_lut (.I0(n1854), .I1(n1921), .I2(n1877), .I3(GND_net), 
            .O(n1953));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1262_rep_44_3_lut (.I0(n1853), .I1(n1920), .I2(n1877), 
            .I3(GND_net), .O(n1952));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1262_rep_44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1256_3_lut (.I0(n1847), .I1(n1914), .I2(n1877), .I3(GND_net), 
            .O(n1946));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_2314_24 (.CI(n28461), .I0(n43152), .I1(n392), .CO(n28462));
    SB_LUT4 div_46_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1769 (.I0(n87), .I1(n15808), .I2(GND_net), .I3(GND_net), 
            .O(n15857));
    defparam i1_2_lut_adj_1769.LUT_INIT = 16'hdddd;
    SB_LUT4 rem_4_i1255_3_lut (.I0(n1846), .I1(n1913), .I2(n1877), .I3(GND_net), 
            .O(n1945));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1254_3_lut (.I0(n1845), .I1(n1912), .I2(n1877), .I3(GND_net), 
            .O(n1944));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1265_3_lut (.I0(n1856), .I1(n1923), .I2(n1877), .I3(GND_net), 
            .O(n1955));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1261_rep_45_3_lut (.I0(n1852), .I1(n1919), .I2(n1877), 
            .I3(GND_net), .O(n1951));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1261_rep_45_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1264_3_lut (.I0(n1855), .I1(n1922), .I2(n1877), .I3(GND_net), 
            .O(n1954));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34863_3_lut (.I0(n1653_adj_4847), .I1(n1720), .I2(n1679), 
            .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34864_3_lut (.I0(n1752), .I1(n1819), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1194_3_lut (.I0(n1753), .I1(n1820), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1195_3_lut (.I0(n1754_adj_4834), .I1(n1821), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1192_3_lut (.I0(n1751), .I1(n1818), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651_adj_4845), .I1(n1718), .I2(n1679), 
            .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63_adj_4690), 
            .I2(gearBoxRatio[23]), .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13257_3_lut (.I0(encoder0_position[21]), .I1(n2997), .I2(count_enable), 
            .I3(GND_net), .O(n17986));   // quad.v(35[10] 41[6])
    defparam i13257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i1127_rep_47_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), 
            .I3(GND_net), .O(n1753));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1127_rep_47_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34865_3_lut (.I0(n1553_adj_4849), .I1(n1620), .I2(n1580), 
            .I3(GND_net), .O(n1652_adj_4846));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34866_3_lut (.I0(n1652_adj_4846), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755_adj_4835));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650_adj_4844), .I1(n1717), .I2(n1679), 
            .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754_adj_4834));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757_adj_4837));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756_adj_4836));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650_adj_4844));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648_adj_4841));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4780), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1062_rep_50_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), 
            .I3(GND_net), .O(n1656));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1062_rep_50_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647_adj_4840));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1770 (.I0(n90), .I1(n15854), .I2(GND_net), .I3(GND_net), 
            .O(n15801));
    defparam i1_2_lut_adj_1770.LUT_INIT = 16'hdddd;
    SB_LUT4 add_2314_23_lut (.I0(n534), .I1(n43152), .I2(n533), .I3(n28460), 
            .O(displacement_23__N_229[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i991_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), .I3(GND_net), 
            .O(n1553_adj_4849));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4781), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i994_rep_56_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), 
            .I3(GND_net), .O(n1556));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i994_rep_56_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418), .I2(n1382), .I3(GND_net), 
            .O(n1450));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419), .I2(n1382), .I3(GND_net), 
            .O(n1451));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4825), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420), .I2(n1382), .I3(GND_net), 
            .O(n1452));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4826), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13256_3_lut (.I0(encoder0_position[20]), .I1(n2998), .I2(count_enable), 
            .I3(GND_net), .O(n17985));   // quad.v(35[10] 41[6])
    defparam i13256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_2314_23 (.CI(n28460), .I0(n43152), .I1(n533), .CO(n28461));
    SB_LUT4 i1_2_lut_adj_1771 (.I0(n93), .I1(n15851), .I2(GND_net), .I3(GND_net), 
            .O(n15794));
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_rep_58_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), 
            .I3(GND_net), .O(n1356));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i858_rep_58_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4824), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4827), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4782), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4831), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4832), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i584_3_lut (.I0(n852), .I1(n6_adj_5304), .I2(n884), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i584_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4828), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i722_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), .I3(GND_net), 
            .O(n1156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2314_22_lut (.I0(n672), .I1(n43152), .I2(n671), .I3(n28459), 
            .O(displacement_23__N_229[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4829), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4830), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19929_4_lut (.I0(n954), .I1(n953), .I2(n35529), .I3(n955), 
            .O(n986));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19929_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 rem_4_i586_3_lut (.I0(n749), .I1(n855), .I2(n884), .I3(GND_net), 
            .O(n956));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i586_3_lut.LUT_INIT = 16'h9a9a;
    SB_LUT4 i1_3_lut_adj_1772 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n35527));
    defparam i1_3_lut_adj_1772.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1773 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n37566));
    defparam i1_2_lut_adj_1773.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n1052), .I1(n37566), .I2(n1053), .I3(n35527), 
            .O(n1085));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfefa;
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1775 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n37570));
    defparam i1_2_lut_adj_1775.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n1154), .I1(n37570), .I2(n1155), .I3(n1157), 
            .O(n35523));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_1777 (.I0(n35523), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1778 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n35521));
    defparam i1_3_lut_adj_1778.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n1254), .I1(n1250), .I2(n35521), .I3(n1255), 
            .O(n6_adj_5251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1780 (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_5251), 
            .O(n1283));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1781 (.I0(n96), .I1(n15788), .I2(GND_net), .I3(GND_net), 
            .O(n15785));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'hdddd;
    SB_CARRY add_2314_22 (.CI(n28459), .I0(n43152), .I1(n671), .CO(n28460));
    SB_LUT4 div_46_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1782 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n35517));
    defparam i1_3_lut_adj_1782.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(n1351), .I1(n1354), .I2(n35517), .I3(n1355), 
            .O(n8_adj_4691));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i2_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1783 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4693));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1783.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1784 (.I0(n1352), .I1(n7_adj_4693), .I2(n1353), 
            .I3(n8_adj_4691), .O(n1382));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417), .I2(n1382), .I3(GND_net), 
            .O(n1449));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1785 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n37678));
    defparam i1_2_lut_adj_1785.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n1454), .I1(n37678), .I2(n1455), .I3(n1457), 
            .O(n35551));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1787 (.I0(n35551), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_5258));
    defparam i5_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1453), .I1(n12_adj_5258), .I2(n1449), .I3(n1448), 
            .O(n1481));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i926_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), .I3(GND_net), 
            .O(n1456));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554_adj_4850));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1788 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n35548));
    defparam i1_3_lut_adj_1788.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1789 (.I0(n558), .I1(n99), .I2(n224), .I3(n15845), 
            .O(n248));
    defparam i2_4_lut_adj_1789.LUT_INIT = 16'hff37;
    SB_LUT4 i36322_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n43152));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i36322_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2314_21_lut (.I0(n807), .I1(n43152), .I2(n806), .I3(n28458), 
            .O(displacement_23__N_229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12733_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n15626), 
            .I3(n4_adj_4713), .O(n17462));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12733_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3_4_lut_adj_1790 (.I0(n1554_adj_4850), .I1(n1551), .I2(n35548), 
            .I3(n1555), .O(n11_adj_5262));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1790.LUT_INIT = 16'heccc;
    SB_LUT4 i5_4_lut_adj_1791 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_5261));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1791.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1792 (.I0(n13_adj_5261), .I1(n11_adj_5262), .I2(n1553_adj_4849), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1792.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i990_rep_53_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), 
            .I3(GND_net), .O(n1552));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i990_rep_53_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651_adj_4845));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1059_3_lut (.I0(n1554_adj_4850), .I1(n1621), .I2(n1580), 
            .I3(GND_net), .O(n1653_adj_4847));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1793 (.I0(n1647_adj_4840), .I1(n1646_adj_4839), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4869));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1793.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1794 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n35565));
    defparam i1_3_lut_adj_1794.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1795 (.I0(n1653_adj_4847), .I1(n1652_adj_4846), 
            .I2(n1651_adj_4845), .I3(n10_adj_4869), .O(n16_adj_4858));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1796 (.I0(n1648_adj_4841), .I1(n1654), .I2(n35565), 
            .I3(n1655), .O(n11_adj_4868));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i2_4_lut_adj_1796.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut_adj_1797 (.I0(n11_adj_4868), .I1(n16_adj_4858), .I2(n1649_adj_4842), 
            .I3(n1650_adj_4844), .O(n1679));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649_adj_4842));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649_adj_4842), .I1(n1716), .I2(n1679), 
            .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648_adj_4841), .I1(n1715), .I2(n1679), 
            .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647_adj_4840), .I1(n1714), .I2(n1679), 
            .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1798 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16_adj_4759));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1799 (.I0(n1756_adj_4836), .I1(n1757_adj_4837), 
            .I2(n1758_adj_4838), .I3(GND_net), .O(n35557));
    defparam i1_3_lut_adj_1799.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1751), .I1(n16_adj_4759), .I2(n1753), .I3(GND_net), 
            .O(n18_adj_4758));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1800 (.I0(n1754_adj_4834), .I1(n1749), .I2(n35557), 
            .I3(n1755_adj_4835), .O(n13_adj_4760));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1800.LUT_INIT = 16'heccc;
    SB_LUT4 i9_4_lut_adj_1801 (.I0(n13_adj_4760), .I1(n18_adj_4758), .I2(n1752), 
            .I3(n1750), .O(n1778_adj_4833));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1801.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4779), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758_adj_4838));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12734_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n36115), .I3(GND_net), .O(n17463));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12735_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n36115), .I3(GND_net), .O(n17464));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12736_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n36115), .I3(GND_net), .O(n17465));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12737_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n36115), .I3(GND_net), .O(n17466));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758_adj_4838), .I1(n1825), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756_adj_4836), .I1(n1823), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755_adj_4835), .I1(n1822), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1198_rep_46_3_lut (.I0(n1757_adj_4837), .I1(n1824), .I2(n1778_adj_4833), 
            .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1198_rep_46_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1802 (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n37832));
    defparam i1_2_lut_adj_1802.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n1854), .I1(n37832), .I2(n1855), .I3(n1857), 
            .O(n35588));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'ha080;
    SB_LUT4 i7_4_lut_adj_1804 (.I0(n1847), .I1(n1846), .I2(n1850), .I3(n35588), 
            .O(n18_adj_4685));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1849), .I1(n1853), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4686));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1805 (.I0(n1851), .I1(n18_adj_4685), .I2(n1845), 
            .I3(n1844), .O(n20_adj_4684));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1806 (.I0(n1852), .I1(n20_adj_4684), .I2(n16_adj_4686), 
            .I3(n1848), .O(n1877));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4778), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4777), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1267_3_lut (.I0(n1858), .I1(n1925), .I2(n1877), .I3(GND_net), 
            .O(n1957));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1266_3_lut (.I0(n1857), .I1(n1924), .I2(n1877), .I3(GND_net), 
            .O(n1956));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1807 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n35573));
    defparam i1_3_lut_adj_1807.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1808 (.I0(n1954), .I1(n1951), .I2(n35573), .I3(n1955), 
            .O(n16_adj_4683));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1808.LUT_INIT = 16'heccc;
    SB_LUT4 i7_4_lut_adj_1809 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4681));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1809.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1952), .I1(n1953), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4682));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1810 (.I0(n19_adj_4681), .I1(n1947), .I2(n16_adj_4683), 
            .I3(n1948), .O(n22_adj_4680));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1811 (.I0(n1949), .I1(n22_adj_4680), .I2(n18_adj_4682), 
            .I3(n1950), .O(n1976_adj_5033));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1257_3_lut (.I0(n1848), .I1(n1915), .I2(n1877), .I3(GND_net), 
            .O(n1947));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976_adj_5033), 
            .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12738_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n36115), .I3(GND_net), .O(n17467));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12739_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n36115), .I3(GND_net), .O(n17468));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12739_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13255_3_lut (.I0(encoder0_position[19]), .I1(n2999), .I2(count_enable), 
            .I3(GND_net), .O(n17984));   // quad.v(35[10] 41[6])
    defparam i13255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12740_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n36115), .I3(GND_net), .O(n17469));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12740_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12741_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n36115), .I3(GND_net), .O(n17470));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12741_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12742_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n36115), .I3(GND_net), .O(n17471));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12742_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1405_3_lut_3_lut (.I0(n2093), .I1(n6028), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12743_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n36115), .I3(GND_net), .O(n17472));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12743_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12744_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n36115), .I3(GND_net), .O(n17473));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12744_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12745_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n36115), .I3(GND_net), .O(n17474));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12745_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12746_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n36115), .I3(GND_net), .O(n17475));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12746_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_3_lut (.I0(one_wire_N_513[5]), .I1(one_wire_N_513[9]), .I2(start), 
            .I3(GND_net), .O(n14_adj_5311));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1812 (.I0(one_wire_N_513[6]), .I1(one_wire_N_513[10]), 
            .I2(one_wire_N_513[8]), .I3(one_wire_N_513[11]), .O(n15_adj_5310));
    defparam i6_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1813 (.I0(n15_adj_5310), .I1(state[1]), .I2(n14_adj_5311), 
            .I3(one_wire_N_513[7]), .O(n35462));
    defparam i8_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1408_3_lut_3_lut (.I0(n2093), .I1(n6031), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12747_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n36115), .I3(GND_net), .O(n17476));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12747_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12748_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n36115), .I3(GND_net), .O(n17477));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12748_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2000_3_lut (.I0(n2943), .I1(n3010_adj_4787), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3042));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1999_3_lut (.I0(n2942), .I1(n3009_adj_4788), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3041));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4926));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1998_3_lut (.I0(n2941), .I1(n3008_adj_4789), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3040));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867), .I3(GND_net), 
            .O(n2950_adj_4810));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1943_rep_63_3_lut (.I0(n2854), .I1(n2921), .I2(n2867), 
            .I3(GND_net), .O(n2953_adj_4807));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1943_rep_63_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911), .I2(n2867), .I3(GND_net), 
            .O(n2943));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12749_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n36115), .I3(GND_net), .O(n17478));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12749_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1938_3_lut (.I0(n2849), .I1(n2916), .I2(n2867), .I3(GND_net), 
            .O(n2948_adj_4812));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839), .I1(n2906), .I2(n2867), .I3(GND_net), 
            .O(n2938));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907), .I2(n2867), .I3(GND_net), 
            .O(n2939));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838), .I1(n2905), .I2(n2867), .I3(GND_net), 
            .O(n2937));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912), .I2(n2867), .I3(GND_net), 
            .O(n2944));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1935_3_lut (.I0(n2846), .I1(n2913), .I2(n2867), .I3(GND_net), 
            .O(n2945_adj_4815));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1936_rep_64_3_lut (.I0(n2847), .I1(n2914), .I2(n2867), 
            .I3(GND_net), .O(n2946_adj_4814));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1936_rep_64_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1937_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), .I3(GND_net), 
            .O(n2947_adj_4813));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1942_rep_61_3_lut (.I0(n2853), .I1(n2920), .I2(n2867), 
            .I3(GND_net), .O(n2952_adj_4808));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1942_rep_61_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1941_3_lut (.I0(n2852), .I1(n2919), .I2(n2867), .I3(GND_net), 
            .O(n2951_adj_4809));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910), .I2(n2867), .I3(GND_net), 
            .O(n2942));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1939_rep_62_3_lut (.I0(n2850), .I1(n2917), .I2(n2867), 
            .I3(GND_net), .O(n2949_adj_4811));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1939_rep_62_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837), .I1(n2904), .I2(n2867), .I3(GND_net), 
            .O(n2936));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836), .I1(n2903), .I2(n2867), .I3(GND_net), 
            .O(n2935));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835), .I1(n2902), .I2(n2867), .I3(GND_net), 
            .O(n2934));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867), .I3(GND_net), 
            .O(n2955_adj_4805));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909), .I2(n2867), .I3(GND_net), 
            .O(n2941));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855), .I1(n2922), .I2(n2867), .I3(GND_net), 
            .O(n2954_adj_4806));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1868_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1873_3_lut (.I0(n2752), .I1(n2819), .I2(n2768), .I3(GND_net), 
            .O(n2851));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821), .I2(n2768), .I3(GND_net), 
            .O(n2853));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816), .I2(n2768), .I3(GND_net), 
            .O(n2848));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12750_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n36115), .I3(GND_net), .O(n17479));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12750_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2314_21 (.CI(n28458), .I0(n43152), .I1(n806), .CO(n28459));
    SB_LUT4 i12751_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n36115), .I3(GND_net), .O(n17480));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12751_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2314_20_lut (.I0(n939), .I1(n43152), .I2(n938), .I3(n28457), 
            .O(displacement_23__N_229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1653_6_lut (.I0(GND_net), .I1(n2455_adj_4941), .I2(GND_net), 
            .I3(n28823), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2314_20 (.CI(n28457), .I0(n43152), .I1(n938), .CO(n28458));
    SB_LUT4 i12752_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n36115), .I3(GND_net), .O(n17481));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12752_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12753_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n36115), .I3(GND_net), .O(n17482));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12753_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1653_6 (.CI(n28823), .I0(n2455_adj_4941), .I1(GND_net), 
            .CO(n28824));
    SB_LUT4 rem_4_add_1653_5_lut (.I0(GND_net), .I1(n2456_adj_4940), .I2(VCC_net), 
            .I3(n28822), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2314_19_lut (.I0(n1068), .I1(n43152), .I2(n1067), .I3(n28456), 
            .O(displacement_23__N_229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12754_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n36115), .I3(GND_net), .O(n17483));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12754_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2314_19 (.CI(n28456), .I0(n43152), .I1(n1067), .CO(n28457));
    SB_CARRY rem_4_add_1653_5 (.CI(n28822), .I0(n2456_adj_4940), .I1(VCC_net), 
            .CO(n28823));
    SB_LUT4 rem_4_add_1653_4_lut (.I0(GND_net), .I1(n2457_adj_4939), .I2(VCC_net), 
            .I3(n28821), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2314_18_lut (.I0(n1194), .I1(n43152), .I2(n1193), .I3(n28455), 
            .O(displacement_23__N_229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_18 (.CI(n28455), .I0(n43152), .I1(n1193), .CO(n28456));
    SB_LUT4 add_2314_17_lut (.I0(n1317), .I1(n43152), .I2(n1316), .I3(n28454), 
            .O(displacement_23__N_229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13254_3_lut (.I0(encoder0_position[18]), .I1(n3000), .I2(count_enable), 
            .I3(GND_net), .O(n17983));   // quad.v(35[10] 41[6])
    defparam i13254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1406_3_lut_3_lut (.I0(n2093), .I1(n6029), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13327_3_lut (.I0(setpoint[19]), .I1(n4368), .I2(n36881), 
            .I3(GND_net), .O(n18056));   // verilog/coms.v(126[12] 292[6])
    defparam i13327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12755_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n36115), .I3(GND_net), .O(n17484));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12755_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2314_17 (.CI(n28454), .I0(n43152), .I1(n1316), .CO(n28455));
    SB_LUT4 i12756_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n36115), .I3(GND_net), .O(n17485));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12756_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12757_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n36115), .I3(GND_net), .O(n17486));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12757_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12758_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n36115), .I3(GND_net), .O(n17487));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12758_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2314_16_lut (.I0(n1437), .I1(n43152), .I2(n1436), .I3(n28453), 
            .O(displacement_23__N_229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_16 (.CI(n28453), .I0(n43152), .I1(n1436), .CO(n28454));
    SB_LUT4 add_2314_15_lut (.I0(n1554), .I1(n43152), .I2(n1553), .I3(n28452), 
            .O(displacement_23__N_229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_15 (.CI(n28452), .I0(n43152), .I1(n1553), .CO(n28453));
    SB_LUT4 add_2314_14_lut (.I0(n1668), .I1(n43152), .I2(n1667), .I3(n28451), 
            .O(displacement_23__N_229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_14 (.CI(n28451), .I0(n43152), .I1(n1667), .CO(n28452));
    SB_LUT4 add_2314_13_lut (.I0(n1779), .I1(n43152), .I2(n1778), .I3(n28450), 
            .O(displacement_23__N_229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_13 (.CI(n28450), .I0(n43152), .I1(n1778), .CO(n28451));
    SB_LUT4 add_2314_12_lut (.I0(n1887), .I1(n43152), .I2(n1886), .I3(n28449), 
            .O(displacement_23__N_229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_12 (.CI(n28449), .I0(n43152), .I1(n1886), .CO(n28450));
    SB_LUT4 i13326_3_lut (.I0(setpoint[18]), .I1(n4367), .I2(n36881), 
            .I3(GND_net), .O(n18055));   // verilog/coms.v(126[12] 292[6])
    defparam i13326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2314_11_lut (.I0(n1992), .I1(n43152), .I2(n1991), .I3(n28448), 
            .O(displacement_23__N_229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_11 (.CI(n28448), .I0(n43152), .I1(n1991), .CO(n28449));
    SB_LUT4 add_2314_10_lut (.I0(n2094), .I1(n43152), .I2(n2093), .I3(n28447), 
            .O(displacement_23__N_229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12759_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n36115), .I3(GND_net), .O(n17488));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12759_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1598_3_lut_3_lut (.I0(n2381), .I1(n6089), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13325_3_lut (.I0(setpoint[17]), .I1(n4366), .I2(n36881), 
            .I3(GND_net), .O(n18054));   // verilog/coms.v(126[12] 292[6])
    defparam i13325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12760_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n36115), .I3(GND_net), .O(n17489));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12760_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12761_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n36115), .I3(GND_net), .O(n17490));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12761_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1653_4 (.CI(n28821), .I0(n2457_adj_4939), .I1(VCC_net), 
            .CO(n28822));
    SB_LUT4 rem_4_add_1653_3_lut (.I0(GND_net), .I1(n2458_adj_4938), .I2(GND_net), 
            .I3(n28820), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_3 (.CI(n28820), .I0(n2458_adj_4938), .I1(GND_net), 
            .CO(n28821));
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4870), .I1(VCC_net), 
            .CO(n28820));
    SB_LUT4 rem_4_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4887), .I2(VCC_net), 
            .I3(n28819), .O(n2636_adj_4857)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2314_10 (.CI(n28447), .I0(n43152), .I1(n2093), .CO(n28448));
    SB_LUT4 rem_4_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4886), .I2(VCC_net), 
            .I3(n28818), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_23 (.CI(n28818), .I0(n2538_adj_4886), .I1(VCC_net), 
            .CO(n28819));
    SB_LUT4 add_2314_9_lut (.I0(n2193), .I1(n43152), .I2(n2192), .I3(n28446), 
            .O(displacement_23__N_229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_9 (.CI(n28446), .I0(n43152), .I1(n2192), .CO(n28447));
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4885), .I2(VCC_net), 
            .I3(n28817), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2314_8_lut (.I0(n2289), .I1(n43152), .I2(n2288), .I3(n28445), 
            .O(displacement_23__N_229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1720_22 (.CI(n28817), .I0(n2539_adj_4885), .I1(VCC_net), 
            .CO(n28818));
    SB_CARRY add_2314_8 (.CI(n28445), .I0(n43152), .I1(n2288), .CO(n28446));
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4884), .I2(VCC_net), 
            .I3(n28816), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2314_7_lut (.I0(n2382), .I1(n43152), .I2(n2381), .I3(n28444), 
            .O(displacement_23__N_229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1720_21 (.CI(n28816), .I0(n2540_adj_4884), .I1(VCC_net), 
            .CO(n28817));
    SB_CARRY add_2314_7 (.CI(n28444), .I0(n43152), .I1(n2381), .CO(n28445));
    SB_LUT4 add_2314_6_lut (.I0(n2472), .I1(n43152), .I2(n2471), .I3(n28443), 
            .O(displacement_23__N_229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_6 (.CI(n28443), .I0(n43152), .I1(n2471), .CO(n28444));
    SB_LUT4 add_2314_5_lut (.I0(n2559), .I1(n43152), .I2(n2558), .I3(n28442), 
            .O(displacement_23__N_229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4883), .I2(VCC_net), 
            .I3(n28815), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2314_5 (.CI(n28442), .I0(n43152), .I1(n2558), .CO(n28443));
    SB_CARRY rem_4_add_1720_20 (.CI(n28815), .I0(n2541_adj_4883), .I1(VCC_net), 
            .CO(n28816));
    SB_LUT4 add_2314_4_lut (.I0(n2643), .I1(n43152), .I2(n2642), .I3(n28441), 
            .O(displacement_23__N_229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4882), .I2(VCC_net), 
            .I3(n28814), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2314_4 (.CI(n28441), .I0(n43152), .I1(n2642), .CO(n28442));
    SB_CARRY rem_4_add_1720_19 (.CI(n28814), .I0(n2542_adj_4882), .I1(VCC_net), 
            .CO(n28815));
    SB_LUT4 add_2314_3_lut (.I0(n2724), .I1(n43152), .I2(n2723), .I3(n28440), 
            .O(displacement_23__N_229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2314_3 (.CI(n28440), .I0(n43152), .I1(n2723), .CO(n28441));
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4881), .I2(VCC_net), 
            .I3(n28813), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_18 (.CI(n28813), .I0(n2543_adj_4881), .I1(VCC_net), 
            .CO(n28814));
    SB_LUT4 add_2314_2_lut (.I0(n2802), .I1(n43152), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2314_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4880), .I2(VCC_net), 
            .I3(n28812), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2314_2 (.CI(VCC_net), .I0(n43152), .I1(n2801), .CO(n28440));
    SB_LUT4 add_2313_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n28439), 
            .O(n6164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n28438), 
            .O(n6165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_17 (.CI(n28812), .I0(n2544_adj_4880), .I1(VCC_net), 
            .CO(n28813));
    SB_CARRY add_2313_24 (.CI(n28438), .I0(n2700), .I1(n79), .CO(n28439));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4879), .I2(VCC_net), 
            .I3(n28811), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n28437), 
            .O(n6166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_23 (.CI(n28437), .I0(n2701), .I1(n80), .CO(n28438));
    SB_CARRY rem_4_add_1720_16 (.CI(n28811), .I0(n2545_adj_4879), .I1(VCC_net), 
            .CO(n28812));
    SB_LUT4 add_2313_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n28436), 
            .O(n6167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_22 (.CI(n28436), .I0(n2702), .I1(n81), .CO(n28437));
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4878), .I2(VCC_net), 
            .I3(n28810), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n28435), 
            .O(n6168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_21 (.CI(n28435), .I0(n2703), .I1(n82), .CO(n28436));
    SB_LUT4 add_2313_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n28434), 
            .O(n6169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13324_3_lut (.I0(setpoint[16]), .I1(n4365), .I2(n36881), 
            .I3(GND_net), .O(n18053));   // verilog/coms.v(126[12] 292[6])
    defparam i13324_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_20 (.CI(n28434), .I0(n2704), .I1(n83), .CO(n28435));
    SB_LUT4 add_2313_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n28433), 
            .O(n6170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_15 (.CI(n28810), .I0(n2546_adj_4878), .I1(VCC_net), 
            .CO(n28811));
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4877), .I2(VCC_net), 
            .I3(n28809), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_19 (.CI(n28433), .I0(n2705), .I1(n84), .CO(n28434));
    SB_CARRY rem_4_add_1720_14 (.CI(n28809), .I0(n2547_adj_4877), .I1(VCC_net), 
            .CO(n28810));
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4876), .I2(VCC_net), 
            .I3(n28808), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n28432), 
            .O(n6171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_13 (.CI(n28808), .I0(n2548_adj_4876), .I1(VCC_net), 
            .CO(n28809));
    SB_CARRY add_2313_18 (.CI(n28432), .I0(n2706), .I1(n85), .CO(n28433));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4875), .I2(VCC_net), 
            .I3(n28807), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n28431), 
            .O(n6172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_17 (.CI(n28431), .I0(n2707), .I1(n86), .CO(n28432));
    SB_CARRY rem_4_add_1720_12 (.CI(n28807), .I0(n2549_adj_4875), .I1(VCC_net), 
            .CO(n28808));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4874), .I2(VCC_net), 
            .I3(n28806), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n28430), 
            .O(n6173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12762_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n36115), .I3(GND_net), .O(n17491));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12762_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12763_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n36115), .I3(GND_net), .O(n17492));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12763_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13323_3_lut (.I0(setpoint[15]), .I1(n4364), .I2(n36881), 
            .I3(GND_net), .O(n18052));   // verilog/coms.v(126[12] 292[6])
    defparam i13323_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1720_11 (.CI(n28806), .I0(n2550_adj_4874), .I1(VCC_net), 
            .CO(n28807));
    SB_CARRY add_2313_16 (.CI(n28430), .I0(n2708), .I1(n87), .CO(n28431));
    SB_LUT4 add_2313_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n28429), 
            .O(n6174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4873), .I2(VCC_net), 
            .I3(n28805), .O(n2618_adj_4867)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_15 (.CI(n28429), .I0(n2709), .I1(n88), .CO(n28430));
    SB_LUT4 i13322_3_lut (.I0(setpoint[14]), .I1(n4363), .I2(n36881), 
            .I3(GND_net), .O(n18051));   // verilog/coms.v(126[12] 292[6])
    defparam i13322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12764_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n36115), .I3(GND_net), .O(n17493));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12764_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13321_3_lut (.I0(setpoint[13]), .I1(n4362), .I2(n36881), 
            .I3(GND_net), .O(n18050));   // verilog/coms.v(126[12] 292[6])
    defparam i13321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1407_3_lut_3_lut (.I0(n2093), .I1(n6030), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13320_3_lut (.I0(setpoint[12]), .I1(n4361), .I2(n36881), 
            .I3(GND_net), .O(n18049));   // verilog/coms.v(126[12] 292[6])
    defparam i13320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1403_3_lut_3_lut (.I0(n2093), .I1(n6026), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_3_lut_adj_1814 (.I0(n40227), .I1(bit_ctr[11]), .I2(n4442), 
            .I3(GND_net), .O(n33439));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1814.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1815 (.I0(bit_ctr[12]), .I1(n40228), .I2(n4442), 
            .I3(GND_net), .O(n33441));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1815.LUT_INIT = 16'hacac;
    SB_LUT4 i12723_3_lut (.I0(n17180), .I1(r_Bit_Index[0]), .I2(n17052), 
            .I3(GND_net), .O(n17452));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12723_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i12_3_lut_adj_1816 (.I0(n40276), .I1(byte_transmit_counter[0]), 
            .I2(n24391), .I3(GND_net), .O(n34173));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut_adj_1816.LUT_INIT = 16'hcaca;
    SB_LUT4 i12717_3_lut (.I0(n17189), .I1(r_Bit_Index_adj_5381[0]), .I2(n17058), 
            .I3(GND_net), .O(n17446));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12717_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i13319_3_lut (.I0(setpoint[11]), .I1(n4360), .I2(n36881), 
            .I3(GND_net), .O(n18048));   // verilog/coms.v(126[12] 292[6])
    defparam i13319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12772_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17501));   // verilog/coms.v(126[12] 292[6])
    defparam i12772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12773_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17502));   // verilog/coms.v(126[12] 292[6])
    defparam i12773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12774_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17503));   // verilog/coms.v(126[12] 292[6])
    defparam i12774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1871_3_lut (.I0(n2750), .I1(n2817), .I2(n2768), .I3(GND_net), 
            .O(n2849));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1874_3_lut (.I0(n2753), .I1(n2820), .I2(n2768), .I3(GND_net), 
            .O(n2852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12775_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17504));   // verilog/coms.v(126[12] 292[6])
    defparam i12775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1872_3_lut (.I0(n2751), .I1(n2818), .I2(n2768), .I3(GND_net), 
            .O(n2850));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1869_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), .I3(GND_net), 
            .O(n2847));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4769), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825), .I2(n2768), .I3(GND_net), 
            .O(n2857));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824), .I2(n2768), .I3(GND_net), 
            .O(n2856));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12776_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17505));   // verilog/coms.v(126[12] 292[6])
    defparam i12776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1817 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n35608));
    defparam i1_3_lut_adj_1817.LUT_INIT = 16'hfefe;
    SB_LUT4 i12777_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17506));   // verilog/coms.v(126[12] 292[6])
    defparam i12777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12778_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17507));   // verilog/coms.v(126[12] 292[6])
    defparam i12778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33_adj_4765), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3360));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12779_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17508));   // verilog/coms.v(126[12] 292[6])
    defparam i12779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12780_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17509));   // verilog/coms.v(126[12] 292[6])
    defparam i12780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12781_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17510));   // verilog/coms.v(126[12] 292[6])
    defparam i12781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12782_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17511));   // verilog/coms.v(126[12] 292[6])
    defparam i12782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36270_1_lut (.I0(n3457), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43102));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36270_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2287_3_lut (.I0(n3358), .I1(n10199), .I2(n3362), .I3(GND_net), 
            .O(n3457));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_2313_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n28428), 
            .O(n6175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_10 (.CI(n28805), .I0(n2551_adj_4873), .I1(VCC_net), 
            .CO(n28806));
    SB_CARRY add_2313_14 (.CI(n28428), .I0(n2710), .I1(n89), .CO(n28429));
    SB_LUT4 add_2313_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n28427), 
            .O(n6176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_13 (.CI(n28427), .I0(n2711), .I1(n90), .CO(n28428));
    SB_LUT4 i12783_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17512));   // verilog/coms.v(126[12] 292[6])
    defparam i12783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2313_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n28426), 
            .O(n6177)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12784_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17513));   // verilog/coms.v(126[12] 292[6])
    defparam i12784_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_12 (.CI(n28426), .I0(n2712), .I1(n91), .CO(n28427));
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4872), .I2(VCC_net), 
            .I3(n28804), .O(n2619_adj_4866)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n28425), 
            .O(n6178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12785_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17514));   // verilog/coms.v(126[12] 292[6])
    defparam i12785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12786_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17515));   // verilog/coms.v(126[12] 292[6])
    defparam i12786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13331_3_lut (.I0(setpoint[23]), .I1(n4372), .I2(n36881), 
            .I3(GND_net), .O(n18060));   // verilog/coms.v(126[12] 292[6])
    defparam i13331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12787_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17516));   // verilog/coms.v(126[12] 292[6])
    defparam i12787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12788_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17517));   // verilog/coms.v(126[12] 292[6])
    defparam i12788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12789_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17518));   // verilog/coms.v(126[12] 292[6])
    defparam i12789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36267_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43099));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36267_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1402_3_lut_3_lut (.I0(n2093), .I1(n6025), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n10198), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12790_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17519));   // verilog/coms.v(126[12] 292[6])
    defparam i12790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13330_3_lut (.I0(setpoint[22]), .I1(n4371), .I2(n36881), 
            .I3(GND_net), .O(n18059));   // verilog/coms.v(126[12] 292[6])
    defparam i13330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12791_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17520));   // verilog/coms.v(126[12] 292[6])
    defparam i12791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12792_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17521));   // verilog/coms.v(126[12] 292[6])
    defparam i12792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1409_3_lut_3_lut (.I0(n2093), .I1(n6032), .I2(n662), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36264_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43096));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36264_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n10197), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12793_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17522));   // verilog/coms.v(126[12] 292[6])
    defparam i12793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12794_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17523));   // verilog/coms.v(126[12] 292[6])
    defparam i12794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1818 (.I0(bit_ctr[2]), .I1(n40235), .I2(n4442), 
            .I3(GND_net), .O(n33459));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1818.LUT_INIT = 16'hacac;
    SB_LUT4 i12796_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[22] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17525));   // verilog/coms.v(126[12] 292[6])
    defparam i12796_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1720_9 (.CI(n28804), .I0(n2552_adj_4872), .I1(VCC_net), 
            .CO(n28805));
    SB_LUT4 i12797_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[22] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17526));   // verilog/coms.v(126[12] 292[6])
    defparam i12797_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_11 (.CI(n28425), .I0(n2713), .I1(n92), .CO(n28426));
    SB_LUT4 add_2313_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n28424), 
            .O(n6179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_10 (.CI(n28424), .I0(n2714), .I1(n93), .CO(n28425));
    SB_LUT4 i12798_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[22] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17527));   // verilog/coms.v(126[12] 292[6])
    defparam i12798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1400_3_lut_3_lut (.I0(n2093), .I1(n6023), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2313_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n28423), 
            .O(n6180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12799_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[22] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17528));   // verilog/coms.v(126[12] 292[6])
    defparam i12799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12800_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[22] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17529));   // verilog/coms.v(126[12] 292[6])
    defparam i12800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13329_3_lut (.I0(setpoint[21]), .I1(n4370), .I2(n36881), 
            .I3(GND_net), .O(n18058));   // verilog/coms.v(126[12] 292[6])
    defparam i13329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13328_3_lut (.I0(setpoint[20]), .I1(n4369), .I2(n36881), 
            .I3(GND_net), .O(n18057));   // verilog/coms.v(126[12] 292[6])
    defparam i13328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12801_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[22] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17530));   // verilog/coms.v(126[12] 292[6])
    defparam i12801_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12802_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[22] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17531));   // verilog/coms.v(126[12] 292[6])
    defparam i12802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1819 (.I0(bit_ctr[16]), .I1(n40237), .I2(n4442), 
            .I3(GND_net), .O(n33463));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1819.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_9 (.CI(n28423), .I0(n2715), .I1(n94), .CO(n28424));
    SB_LUT4 i13338_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1172), .I3(GND_net), .O(n18067));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4871), .I2(VCC_net), 
            .I3(n28803), .O(n2620_adj_4865)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n28647), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2313_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n28422), 
            .O(n6181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36261_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43093));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36261_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n10196), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12803_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[21] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17532));   // verilog/coms.v(126[12] 292[6])
    defparam i12803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12804_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[21] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17533));   // verilog/coms.v(126[12] 292[6])
    defparam i12804_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_8 (.CI(n28422), .I0(n2716), .I1(n95), .CO(n28423));
    SB_LUT4 add_2313_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n28421), 
            .O(n6182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12805_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[21] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17534));   // verilog/coms.v(126[12] 292[6])
    defparam i12805_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_7 (.CI(n28421), .I0(n2717), .I1(n96), .CO(n28422));
    SB_LUT4 add_2313_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n28420), 
            .O(n6183)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36258_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43090));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36258_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2313_6 (.CI(n28420), .I0(n2718), .I1(n97), .CO(n28421));
    SB_LUT4 add_2313_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n28419), 
            .O(n6184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n10195), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12806_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[21] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17535));   // verilog/coms.v(126[12] 292[6])
    defparam i12806_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2313_5 (.CI(n28419), .I0(n2719), .I1(n98), .CO(n28420));
    SB_LUT4 add_2313_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n28418), 
            .O(n6185)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_4 (.CI(n28418), .I0(n2720), .I1(n99), .CO(n28419));
    SB_LUT4 add_2313_3_lut (.I0(GND_net), .I1(n669), .I2(n558), .I3(n28417), 
            .O(n6186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2313_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2313_3 (.CI(n28417), .I0(n669), .I1(n558), .CO(n28418));
    SB_CARRY add_2313_2 (.CI(VCC_net), .I0(n670), .I1(VCC_net), .CO(n28417));
    SB_LUT4 add_2312_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n28416), 
            .O(n6140)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2312_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n28415), 
            .O(n6141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_14_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n28992), .O(n1646_adj_4839)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1720_8 (.CI(n28803), .I0(n2553_adj_4871), .I1(VCC_net), 
            .CO(n28804));
    SB_CARRY add_2312_22 (.CI(n28415), .I0(n2619), .I1(n80), .CO(n28416));
    SB_LUT4 i12807_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[21] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17536));   // verilog/coms.v(126[12] 292[6])
    defparam i12807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1820 (.I0(bit_ctr[24]), .I1(n40247), .I2(n4442), 
            .I3(GND_net), .O(n33483));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1820.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n28802), .O(n2621_adj_4864)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2312_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n28414), 
            .O(n6142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_21 (.CI(n28414), .I0(n2620), .I1(n81), .CO(n28415));
    SB_LUT4 add_2312_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n28413), 
            .O(n6143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_20 (.CI(n28413), .I0(n2621), .I1(n82), .CO(n28414));
    SB_LUT4 add_2312_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n28412), 
            .O(n6144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_13_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n28991), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_13 (.CI(n28991), .I0(n1548), .I1(VCC_net), 
            .CO(n28992));
    SB_CARRY add_2312_19 (.CI(n28412), .I0(n2622), .I1(n83), .CO(n28413));
    SB_LUT4 i12808_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[21] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17537));   // verilog/coms.v(126[12] 292[6])
    defparam i12808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12809_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[21] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17538));   // verilog/coms.v(126[12] 292[6])
    defparam i12809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1821 (.I0(n3341), .I1(n3348), .I2(n3351), .I3(n3350), 
            .O(n37660));
    defparam i1_4_lut_adj_1821.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2312_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n28411), 
            .O(n6145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(n3343), .I1(n3352), .I2(n3344), .I3(n3342), 
            .O(n37610));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1823 (.I0(n3338), .I1(n3339), .I2(n37660), .I3(GND_net), 
            .O(n37664));
    defparam i1_3_lut_adj_1823.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(n3347), .I1(n3353), .I2(n3346), .I3(n3349), 
            .O(n37684));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1825 (.I0(n3356), .I1(n3357), .I2(n3358), .I3(GND_net), 
            .O(n35641));
    defparam i1_3_lut_adj_1825.LUT_INIT = 16'hfefe;
    SB_CARRY add_2312_18 (.CI(n28411), .I0(n2623), .I1(n84), .CO(n28412));
    SB_LUT4 i1_3_lut_adj_1826 (.I0(n37610), .I1(n3340), .I2(n3345), .I3(GND_net), 
            .O(n37612));
    defparam i1_3_lut_adj_1826.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n28990), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_7 (.CI(n28802), .I0(n2554), .I1(GND_net), 
            .CO(n28803));
    SB_LUT4 add_2312_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n28410), 
            .O(n6146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_12 (.CI(n28990), .I0(n1549), .I1(VCC_net), 
            .CO(n28991));
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n28801), .O(n2622_adj_4863)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_17 (.CI(n28410), .I0(n2624), .I1(n85), .CO(n28411));
    SB_CARRY rem_4_add_1720_6 (.CI(n28801), .I0(n2555), .I1(GND_net), 
            .CO(n28802));
    SB_LUT4 add_2312_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n28409), 
            .O(n6147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n28989), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n28800), .O(n2623_adj_4862)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_16 (.CI(n28409), .I0(n2625), .I1(n86), .CO(n28410));
    SB_LUT4 add_2312_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n28408), 
            .O(n6148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_5 (.CI(n28800), .I0(n2556), .I1(VCC_net), 
            .CO(n28801));
    SB_CARRY rem_4_add_1050_11 (.CI(n28989), .I0(n1550), .I1(VCC_net), 
            .CO(n28990));
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n28799), .O(n2624_adj_4861)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_15 (.CI(n28408), .I0(n2626), .I1(n87), .CO(n28409));
    SB_LUT4 add_2312_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n28407), 
            .O(n6149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_4 (.CI(n28799), .I0(n2557), .I1(VCC_net), 
            .CO(n28800));
    SB_CARRY add_2312_14 (.CI(n28407), .I0(n2627), .I1(n88), .CO(n28408));
    SB_LUT4 add_2312_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n28406), 
            .O(n6150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n3354), .I1(n37612), .I2(n35641), .I3(n3355), 
            .O(n37614));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(n3335), .I1(n37684), .I2(n3334), .I3(n37664), 
            .O(n37686));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(n3336), .I1(n37686), .I2(n3332), .I3(n37614), 
            .O(n37688));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1830 (.I0(n3331), .I1(n3333), .I2(n3337), .I3(GND_net), 
            .O(n37474));
    defparam i1_3_lut_adj_1830.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n3329), .I1(n37474), .I2(n37688), .I3(n3330), 
            .O(n3362));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_LUT4 i36257_2_lut (.I0(n3362), .I1(n10194), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36257_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5272));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12810_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[21] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17539));   // verilog/coms.v(126[12] 292[6])
    defparam i12810_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12811_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[20] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17540));   // verilog/coms.v(126[12] 292[6])
    defparam i12811_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12812_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[20] [1]), 
            .I2(n30070), .I3(GND_net), .O(n17541));   // verilog/coms.v(126[12] 292[6])
    defparam i12812_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12813_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[20] [2]), 
            .I2(n30070), .I3(GND_net), .O(n17542));   // verilog/coms.v(126[12] 292[6])
    defparam i12813_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12814_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[20] [3]), 
            .I2(n30070), .I3(GND_net), .O(n17543));   // verilog/coms.v(126[12] 292[6])
    defparam i12814_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12815_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[20] [4]), 
            .I2(n30070), .I3(GND_net), .O(n17544));   // verilog/coms.v(126[12] 292[6])
    defparam i12815_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12816_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[20] [5]), 
            .I2(n30070), .I3(GND_net), .O(n17545));   // verilog/coms.v(126[12] 292[6])
    defparam i12816_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12817_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[20] [6]), 
            .I2(n30070), .I3(GND_net), .O(n17546));   // verilog/coms.v(126[12] 292[6])
    defparam i12817_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12818_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[20] [7]), 
            .I2(n30070), .I3(GND_net), .O(n17547));   // verilog/coms.v(126[12] 292[6])
    defparam i12818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12819_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n30070), 
            .I3(GND_net), .O(n17548));   // verilog/coms.v(126[12] 292[6])
    defparam i12819_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12820_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n30070), 
            .I3(GND_net), .O(n17549));   // verilog/coms.v(126[12] 292[6])
    defparam i12820_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12821_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n30070), 
            .I3(GND_net), .O(n17550));   // verilog/coms.v(126[12] 292[6])
    defparam i12821_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12822_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n30070), 
            .I3(GND_net), .O(n17551));   // verilog/coms.v(126[12] 292[6])
    defparam i12822_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2312_13 (.CI(n28406), .I0(n2628), .I1(n89), .CO(n28407));
    SB_LUT4 add_2312_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n28405), 
            .O(n6151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n28988), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4870), .I2(GND_net), 
            .I3(n28798), .O(n2625_adj_4860)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_12 (.CI(n28405), .I0(n2629), .I1(n90), .CO(n28406));
    SB_CARRY rem_4_add_1050_10 (.CI(n28988), .I0(n1551), .I1(VCC_net), 
            .CO(n28989));
    SB_CARRY rem_4_add_1720_3 (.CI(n28798), .I0(n2558_adj_4870), .I1(GND_net), 
            .CO(n28799));
    SB_LUT4 add_2312_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n28404), 
            .O(n6152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_11 (.CI(n28404), .I0(n2630), .I1(n91), .CO(n28405));
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n28987), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2312_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n28403), 
            .O(n6153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_10 (.CI(n28403), .I0(n2631), .I1(n92), .CO(n28404));
    SB_LUT4 add_2312_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n28402), 
            .O(n6154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_9 (.CI(n28402), .I0(n2632), .I1(n93), .CO(n28403));
    SB_LUT4 add_2312_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n28401), 
            .O(n6155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_8 (.CI(n28401), .I0(n2633), .I1(n94), .CO(n28402));
    SB_LUT4 add_2312_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n28400), 
            .O(n6156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_7 (.CI(n28400), .I0(n2634), .I1(n95), .CO(n28401));
    SB_LUT4 add_2312_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n28399), 
            .O(n6157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_6 (.CI(n28399), .I0(n2635), .I1(n96), .CO(n28400));
    SB_LUT4 add_2312_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n28398), 
            .O(n6158)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_5 (.CI(n28398), .I0(n2636), .I1(n97), .CO(n28399));
    SB_LUT4 add_2312_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n28397), 
            .O(n6159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_4 (.CI(n28397), .I0(n2637), .I1(n98), .CO(n28398));
    SB_LUT4 add_2312_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n28396), 
            .O(n6160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_3 (.CI(n28396), .I0(n2638), .I1(n99), .CO(n28397));
    SB_LUT4 add_2312_2_lut (.I0(GND_net), .I1(n668), .I2(n558), .I3(VCC_net), 
            .O(n6161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2312_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2312_2 (.CI(VCC_net), .I0(n668), .I1(n558), .CO(n28396));
    SB_LUT4 add_2311_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n28395), 
            .O(n6117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2311_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n28394), 
            .O(n6118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_21 (.CI(n28394), .I0(n2535), .I1(n81), .CO(n28395));
    SB_LUT4 add_2311_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n28393), 
            .O(n6119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_20 (.CI(n28393), .I0(n2536), .I1(n82), .CO(n28394));
    SB_LUT4 add_2311_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n28392), 
            .O(n6120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_19 (.CI(n28392), .I0(n2537), .I1(n83), .CO(n28393));
    SB_LUT4 add_2311_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n28391), 
            .O(n6121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_18 (.CI(n28391), .I0(n2538), .I1(n84), .CO(n28392));
    SB_LUT4 add_2311_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n28390), 
            .O(n6122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_17 (.CI(n28390), .I0(n2539), .I1(n85), .CO(n28391));
    SB_LUT4 add_2311_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n28389), 
            .O(n6123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1832 (.I0(bit_ctr[23]), .I1(n40246), .I2(n4442), 
            .I3(GND_net), .O(n33481));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1832.LUT_INIT = 16'hacac;
    SB_LUT4 i12823_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n30070), 
            .I3(GND_net), .O(n17552));   // verilog/coms.v(126[12] 292[6])
    defparam i12823_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822), .I2(n2768), .I3(GND_net), 
            .O(n2854));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1833 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4703));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1833.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1834 (.I0(n2856), .I1(n2857), .I2(n2858), .I3(GND_net), 
            .O(n35679));
    defparam i1_3_lut_adj_1834.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1835 (.I0(n2847), .I1(n2850), .I2(n2852), .I3(n2849), 
            .O(n36));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1836 (.I0(n2854), .I1(n2844), .I2(n35679), .I3(n2855), 
            .O(n27));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_4_lut_adj_1836.LUT_INIT = 16'heccc;
    SB_CARRY add_2311_16 (.CI(n28389), .I0(n2540), .I1(n86), .CO(n28390));
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2658), .I1(VCC_net), 
            .CO(n28798));
    SB_LUT4 i12824_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n30070), 
            .I3(GND_net), .O(n17553));   // verilog/coms.v(126[12] 292[6])
    defparam i12824_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2311_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n28388), 
            .O(n6124)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12825_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n30070), 
            .I3(GND_net), .O(n17554));   // verilog/coms.v(126[12] 292[6])
    defparam i12825_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2311_15 (.CI(n28388), .I0(n2541), .I1(n87), .CO(n28389));
    SB_LUT4 i12826_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n30070), 
            .I3(GND_net), .O(n17555));   // verilog/coms.v(126[12] 292[6])
    defparam i12826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2311_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n28387), 
            .O(n6125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_14 (.CI(n28387), .I0(n2542), .I1(n88), .CO(n28388));
    SB_LUT4 i22_3_lut_adj_1837 (.I0(bit_ctr[4]), .I1(n40245), .I2(n4442), 
            .I3(GND_net), .O(n33479));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1837.LUT_INIT = 16'hacac;
    SB_LUT4 i12828_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n30070), 
            .I3(GND_net), .O(n17557));   // verilog/coms.v(126[12] 292[6])
    defparam i12828_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13275_3_lut (.I0(encoder1_position[15]), .I1(n2953), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18004));   // quad.v(35[10] 41[6])
    defparam i13275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2311_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n28386), 
            .O(n6126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_13 (.CI(n28386), .I0(n2543), .I1(n89), .CO(n28387));
    SB_LUT4 i13274_3_lut (.I0(encoder1_position[14]), .I1(n2954), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n18003));   // quad.v(35[10] 41[6])
    defparam i13274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12829_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n30070), 
            .I3(GND_net), .O(n17558));   // verilog/coms.v(126[12] 292[6])
    defparam i12829_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12830_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n30070), 
            .I3(GND_net), .O(n17559));   // verilog/coms.v(126[12] 292[6])
    defparam i12830_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1838 (.I0(bit_ctr[26]), .I1(n40249), .I2(n4442), 
            .I3(GND_net), .O(n33487));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1838.LUT_INIT = 16'hacac;
    SB_LUT4 i12831_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n30070), 
            .I3(GND_net), .O(n17560));   // verilog/coms.v(126[12] 292[6])
    defparam i12831_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1839 (.I0(bit_ctr[25]), .I1(n40248), .I2(n4442), 
            .I3(GND_net), .O(n33485));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1839.LUT_INIT = 16'hacac;
    SB_LUT4 add_2311_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n28385), 
            .O(n6127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_9 (.CI(n28987), .I0(n1552), .I1(VCC_net), 
            .CO(n28988));
    SB_LUT4 i12832_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n30070), 
            .I3(GND_net), .O(n17561));   // verilog/coms.v(126[12] 292[6])
    defparam i12832_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12833_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n30070), 
            .I3(GND_net), .O(n17562));   // verilog/coms.v(126[12] 292[6])
    defparam i12833_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2311_12 (.CI(n28385), .I0(n2544), .I1(n90), .CO(n28386));
    SB_LUT4 i12834_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n30070), 
            .I3(GND_net), .O(n17563));   // verilog/coms.v(126[12] 292[6])
    defparam i12834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2311_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n28384), 
            .O(n6128)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_25_lut (.I0(n2636_adj_4857), .I1(n2636_adj_4857), 
            .I2(n2669), .I3(n28797), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2311_11 (.CI(n28384), .I0(n2545), .I1(n91), .CO(n28385));
    SB_LUT4 add_2311_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n28383), 
            .O(n6129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_10 (.CI(n28383), .I0(n2546), .I1(n92), .CO(n28384));
    SB_LUT4 add_2311_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n28382), 
            .O(n6130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_9 (.CI(n28382), .I0(n2547), .I1(n93), .CO(n28383));
    SB_LUT4 add_2311_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n28381), 
            .O(n6131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_8 (.CI(n28381), .I0(n2548), .I1(n94), .CO(n28382));
    SB_LUT4 add_2311_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n28380), 
            .O(n6132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_7 (.CI(n28380), .I0(n2549), .I1(n95), .CO(n28381));
    SB_LUT4 add_2311_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n28379), 
            .O(n6133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_6 (.CI(n28379), .I0(n2550), .I1(n96), .CO(n28380));
    SB_LUT4 add_2311_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n28378), 
            .O(n6134)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_5 (.CI(n28378), .I0(n2551), .I1(n97), .CO(n28379));
    SB_LUT4 add_2311_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n28377), 
            .O(n6135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_4 (.CI(n28377), .I0(n2552), .I1(n98), .CO(n28378));
    SB_LUT4 add_2311_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n28376), 
            .O(n6136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_3 (.CI(n28376), .I0(n2553), .I1(n99), .CO(n28377));
    SB_LUT4 add_2311_2_lut (.I0(GND_net), .I1(n667), .I2(n558), .I3(VCC_net), 
            .O(n6137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2311_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2311_2 (.CI(VCC_net), .I0(n667), .I1(n558), .CO(n28376));
    SB_LUT4 add_2310_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n28375), 
            .O(n6095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2310_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n28374), 
            .O(n6096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_20 (.CI(n28374), .I0(n2448), .I1(n82), .CO(n28375));
    SB_LUT4 add_2310_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n28373), 
            .O(n6097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_19 (.CI(n28373), .I0(n2449), .I1(n83), .CO(n28374));
    SB_LUT4 add_2310_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n28372), 
            .O(n6098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_18 (.CI(n28372), .I0(n2450), .I1(n84), .CO(n28373));
    SB_LUT4 add_2310_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n28371), 
            .O(n6099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_17 (.CI(n28371), .I0(n2451), .I1(n85), .CO(n28372));
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1553_adj_4849), .I2(VCC_net), 
            .I3(n28986), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_24_lut (.I0(n2637_adj_4856), .I1(n2637_adj_4856), 
            .I2(n2669), .I3(n28796), .O(n2736)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2310_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n28370), 
            .O(n6100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_16 (.CI(n28370), .I0(n2452), .I1(n86), .CO(n28371));
    SB_LUT4 add_2310_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n28369), 
            .O(n6101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_15 (.CI(n28369), .I0(n2453), .I1(n87), .CO(n28370));
    SB_LUT4 add_2310_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n28368), 
            .O(n6102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_14 (.CI(n28368), .I0(n2454), .I1(n88), .CO(n28369));
    SB_LUT4 add_2310_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n28367), 
            .O(n6103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_13 (.CI(n28367), .I0(n2455), .I1(n89), .CO(n28368));
    SB_LUT4 add_2310_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n28366), 
            .O(n6104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_12 (.CI(n28366), .I0(n2456), .I1(n90), .CO(n28367));
    SB_LUT4 add_2310_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n28365), 
            .O(n6105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_11 (.CI(n28365), .I0(n2457), .I1(n91), .CO(n28366));
    SB_LUT4 add_2310_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n28364), 
            .O(n6106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_10 (.CI(n28364), .I0(n2458), .I1(n92), .CO(n28365));
    SB_LUT4 add_2310_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n28363), 
            .O(n6107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_9 (.CI(n28363), .I0(n2459), .I1(n93), .CO(n28364));
    SB_LUT4 add_2310_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n28362), 
            .O(n6108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_8 (.CI(n28986), .I0(n1553_adj_4849), .I1(VCC_net), 
            .CO(n28987));
    SB_LUT4 i12835_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n30070), 
            .I3(GND_net), .O(n17564));   // verilog/coms.v(126[12] 292[6])
    defparam i12835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12836_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n30070), 
            .I3(GND_net), .O(n17565));   // verilog/coms.v(126[12] 292[6])
    defparam i12836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12837_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n30070), 
            .I3(GND_net), .O(n17566));   // verilog/coms.v(126[12] 292[6])
    defparam i12837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12838_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n30070), 
            .I3(GND_net), .O(n17567));   // verilog/coms.v(126[12] 292[6])
    defparam i12838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12839_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n30070), 
            .I3(GND_net), .O(n17568));   // verilog/coms.v(126[12] 292[6])
    defparam i12839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12840_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n30070), 
            .I3(GND_net), .O(n17569));   // verilog/coms.v(126[12] 292[6])
    defparam i12840_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2310_8 (.CI(n28362), .I0(n2460), .I1(n94), .CO(n28363));
    SB_LUT4 add_2310_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n28361), 
            .O(n6109)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_7 (.CI(n28361), .I0(n2461), .I1(n95), .CO(n28362));
    SB_LUT4 i12841_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n30070), 
            .I3(GND_net), .O(n17570));   // verilog/coms.v(126[12] 292[6])
    defparam i12841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13335_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1172), .I3(GND_net), .O(n18064));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12842_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n30070), 
            .I3(GND_net), .O(n17571));   // verilog/coms.v(126[12] 292[6])
    defparam i12842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12843_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n30070), 
            .I3(GND_net), .O(n17572));   // verilog/coms.v(126[12] 292[6])
    defparam i12843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12844_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n30070), 
            .I3(GND_net), .O(n17573));   // verilog/coms.v(126[12] 292[6])
    defparam i12844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2310_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n28360), 
            .O(n6110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_6 (.CI(n28360), .I0(n2462), .I1(n96), .CO(n28361));
    SB_CARRY rem_4_add_1787_24 (.CI(n28796), .I0(n2637_adj_4856), .I1(n2669), 
            .CO(n28797));
    SB_LUT4 add_2310_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n28359), 
            .O(n6111)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12845_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n30070), 
            .I3(GND_net), .O(n17574));   // verilog/coms.v(126[12] 292[6])
    defparam i12845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12846_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n30070), 
            .I3(GND_net), .O(n17575));   // verilog/coms.v(126[12] 292[6])
    defparam i12846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12847_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n30070), 
            .I3(GND_net), .O(n17576));   // verilog/coms.v(126[12] 292[6])
    defparam i12847_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2310_5 (.CI(n28359), .I0(n2463), .I1(n97), .CO(n28360));
    SB_LUT4 add_2310_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n28358), 
            .O(n6112)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12848_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n30070), 
            .I3(GND_net), .O(n17577));   // verilog/coms.v(126[12] 292[6])
    defparam i12848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12849_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17578));   // verilog/coms.v(126[12] 292[6])
    defparam i12849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1840 (.I0(bit_ctr[28]), .I1(n40251), .I2(n4442), 
            .I3(GND_net), .O(n33491));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1840.LUT_INIT = 16'hacac;
    SB_LUT4 i12850_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17579));   // verilog/coms.v(126[12] 292[6])
    defparam i12850_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2310_4 (.CI(n28358), .I0(n2464), .I1(n98), .CO(n28359));
    SB_LUT4 add_2310_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n28357), 
            .O(n6113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_3 (.CI(n28357), .I0(n2465), .I1(n99), .CO(n28358));
    SB_LUT4 add_2310_2_lut (.I0(GND_net), .I1(n666), .I2(n558), .I3(VCC_net), 
            .O(n6114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2310_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2310_2 (.CI(VCC_net), .I0(n666), .I1(n558), .CO(n28357));
    SB_LUT4 add_2309_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n28356), 
            .O(n6074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2309_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n28355), 
            .O(n6075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_19 (.CI(n28355), .I0(n2358), .I1(n83), .CO(n28356));
    SB_LUT4 add_2309_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n28354), 
            .O(n6076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_18 (.CI(n28354), .I0(n2359), .I1(n84), .CO(n28355));
    SB_LUT4 add_2309_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n28353), 
            .O(n6077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_17 (.CI(n28353), .I0(n2360), .I1(n85), .CO(n28354));
    SB_LUT4 add_2309_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n28352), 
            .O(n6078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_16 (.CI(n28352), .I0(n2361), .I1(n86), .CO(n28353));
    SB_LUT4 add_2309_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n28351), 
            .O(n6079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_15 (.CI(n28351), .I0(n2362), .I1(n87), .CO(n28352));
    SB_LUT4 add_2309_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n28350), 
            .O(n6080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_14 (.CI(n28350), .I0(n2363), .I1(n88), .CO(n28351));
    SB_LUT4 add_2309_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n28349), 
            .O(n6081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_13 (.CI(n28349), .I0(n2364), .I1(n89), .CO(n28350));
    SB_LUT4 add_2309_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n28348), 
            .O(n6082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_12 (.CI(n28348), .I0(n2365), .I1(n90), .CO(n28349));
    SB_LUT4 add_2309_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n28347), 
            .O(n6083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_11 (.CI(n28347), .I0(n2366), .I1(n91), .CO(n28348));
    SB_LUT4 add_2309_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n28346), 
            .O(n6084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_10 (.CI(n28346), .I0(n2367), .I1(n92), .CO(n28347));
    SB_LUT4 add_2309_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n28345), 
            .O(n6085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_9 (.CI(n28345), .I0(n2368), .I1(n93), .CO(n28346));
    SB_LUT4 add_2309_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n28344), 
            .O(n6086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_8 (.CI(n28344), .I0(n2369), .I1(n94), .CO(n28345));
    SB_LUT4 add_2309_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n28343), 
            .O(n6087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_7 (.CI(n28343), .I0(n2370), .I1(n95), .CO(n28344));
    SB_LUT4 add_2309_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n28342), 
            .O(n6088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_6 (.CI(n28342), .I0(n2371), .I1(n96), .CO(n28343));
    SB_LUT4 add_2309_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n28341), 
            .O(n6089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_5 (.CI(n28341), .I0(n2372), .I1(n97), .CO(n28342));
    SB_LUT4 add_2309_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n28340), 
            .O(n6090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_4 (.CI(n28340), .I0(n2373), .I1(n98), .CO(n28341));
    SB_LUT4 add_2309_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n28339), 
            .O(n6091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_3 (.CI(n28339), .I0(n2374), .I1(n99), .CO(n28340));
    SB_LUT4 add_2309_2_lut (.I0(GND_net), .I1(n665), .I2(n558), .I3(VCC_net), 
            .O(n6092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2309_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2309_2 (.CI(VCC_net), .I0(n665), .I1(n558), .CO(n28339));
    SB_LUT4 add_2308_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n28338), 
            .O(n6054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2308_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n28337), 
            .O(n6055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_18 (.CI(n28337), .I0(n2265), .I1(n84), .CO(n28338));
    SB_LUT4 add_2308_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n28336), 
            .O(n6056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_17 (.CI(n28336), .I0(n2266), .I1(n85), .CO(n28337));
    SB_LUT4 add_2308_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n28335), 
            .O(n6057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_16 (.CI(n28335), .I0(n2267), .I1(n86), .CO(n28336));
    SB_LUT4 add_2308_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n28334), 
            .O(n6058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_15 (.CI(n28334), .I0(n2268), .I1(n87), .CO(n28335));
    SB_LUT4 add_2308_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n28333), 
            .O(n6059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_14 (.CI(n28333), .I0(n2269), .I1(n88), .CO(n28334));
    SB_LUT4 add_2308_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n28332), 
            .O(n6060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_13 (.CI(n28332), .I0(n2270), .I1(n89), .CO(n28333));
    SB_LUT4 add_2308_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n28331), 
            .O(n6061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_12 (.CI(n28331), .I0(n2271), .I1(n90), .CO(n28332));
    SB_LUT4 add_2308_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n28330), 
            .O(n6062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_11 (.CI(n28330), .I0(n2272), .I1(n91), .CO(n28331));
    SB_LUT4 add_2308_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n28329), 
            .O(n6063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_10 (.CI(n28329), .I0(n2273), .I1(n92), .CO(n28330));
    SB_LUT4 add_2308_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n28328), 
            .O(n6064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_9 (.CI(n28328), .I0(n2274), .I1(n93), .CO(n28329));
    SB_LUT4 add_2308_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n28327), 
            .O(n6065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_8 (.CI(n28327), .I0(n2275), .I1(n94), .CO(n28328));
    SB_LUT4 add_2308_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n28326), 
            .O(n6066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_7 (.CI(n28326), .I0(n2276), .I1(n95), .CO(n28327));
    SB_LUT4 add_2308_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n28325), 
            .O(n6067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_6 (.CI(n28325), .I0(n2277), .I1(n96), .CO(n28326));
    SB_LUT4 add_2308_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n28324), 
            .O(n6068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_5 (.CI(n28324), .I0(n2278), .I1(n97), .CO(n28325));
    SB_LUT4 add_2308_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n28323), 
            .O(n6069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_4 (.CI(n28323), .I0(n2279), .I1(n98), .CO(n28324));
    SB_LUT4 add_2308_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n28322), 
            .O(n6070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_3 (.CI(n28322), .I0(n2280), .I1(n99), .CO(n28323));
    SB_LUT4 add_2308_2_lut (.I0(GND_net), .I1(n664), .I2(n558), .I3(VCC_net), 
            .O(n6071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2308_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2308_2 (.CI(VCC_net), .I0(n664), .I1(n558), .CO(n28322));
    SB_LUT4 add_2307_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n28321), 
            .O(n6035)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2307_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n28320), 
            .O(n6036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_17 (.CI(n28320), .I0(n2169), .I1(n85), .CO(n28321));
    SB_LUT4 add_2307_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n28319), 
            .O(n6037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_16 (.CI(n28319), .I0(n2170), .I1(n86), .CO(n28320));
    SB_LUT4 add_2307_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n28318), 
            .O(n6038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_15 (.CI(n28318), .I0(n2171), .I1(n87), .CO(n28319));
    SB_LUT4 add_2307_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n28317), 
            .O(n6039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_14 (.CI(n28317), .I0(n2172), .I1(n88), .CO(n28318));
    SB_LUT4 add_2307_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n28316), 
            .O(n6040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_13 (.CI(n28316), .I0(n2173), .I1(n89), .CO(n28317));
    SB_LUT4 add_2307_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n28315), 
            .O(n6041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_12 (.CI(n28315), .I0(n2174), .I1(n90), .CO(n28316));
    SB_LUT4 add_2307_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n28314), 
            .O(n6042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_11 (.CI(n28314), .I0(n2175), .I1(n91), .CO(n28315));
    SB_LUT4 i33830_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24520), .I3(start), .O(n40256));
    defparam i33830_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 i12851_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17580));   // verilog/coms.v(126[12] 292[6])
    defparam i12851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12852_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17581));   // verilog/coms.v(126[12] 292[6])
    defparam i12852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12853_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17582));   // verilog/coms.v(126[12] 292[6])
    defparam i12853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12854_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17583));   // verilog/coms.v(126[12] 292[6])
    defparam i12854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12855_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17584));   // verilog/coms.v(126[12] 292[6])
    defparam i12855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24520), .I3(state[1]), .O(n36877));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i12856_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17585));   // verilog/coms.v(126[12] 292[6])
    defparam i12856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12857_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17586));   // verilog/coms.v(126[12] 292[6])
    defparam i12857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12858_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17587));   // verilog/coms.v(126[12] 292[6])
    defparam i12858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12859_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17588));   // verilog/coms.v(126[12] 292[6])
    defparam i12859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12860_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17589));   // verilog/coms.v(126[12] 292[6])
    defparam i12860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12861_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17590));   // verilog/coms.v(126[12] 292[6])
    defparam i12861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1841 (.I0(bit_ctr[27]), .I1(n40250), .I2(n4442), 
            .I3(GND_net), .O(n33489));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1841.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_1842 (.I0(n2840), .I1(n2842), .I2(n2841), .I3(n2843), 
            .O(n34));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_LUT4 i12862_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17591));   // verilog/coms.v(126[12] 292[6])
    defparam i12862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12863_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17592));   // verilog/coms.v(126[12] 292[6])
    defparam i12863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1843 (.I0(bit_ctr[30]), .I1(n40253), .I2(n4442), 
            .I3(GND_net), .O(n33495));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1843.LUT_INIT = 16'hacac;
    SB_LUT4 i12864_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17593));   // verilog/coms.v(126[12] 292[6])
    defparam i12864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12865_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17594));   // verilog/coms.v(126[12] 292[6])
    defparam i12865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2307_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n28313), 
            .O(n6043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_10 (.CI(n28313), .I0(n2176), .I1(n92), .CO(n28314));
    SB_LUT4 add_2307_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n28312), 
            .O(n6044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_9 (.CI(n28312), .I0(n2177), .I1(n93), .CO(n28313));
    SB_LUT4 add_2307_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n28311), 
            .O(n6045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_8 (.CI(n28311), .I0(n2178), .I1(n94), .CO(n28312));
    SB_LUT4 add_2307_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n28310), 
            .O(n6046)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_7 (.CI(n28310), .I0(n2179), .I1(n95), .CO(n28311));
    SB_LUT4 add_2307_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n28309), 
            .O(n6047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_6 (.CI(n28309), .I0(n2180), .I1(n96), .CO(n28310));
    SB_LUT4 add_2307_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n28308), 
            .O(n6048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_5 (.CI(n28308), .I0(n2181), .I1(n97), .CO(n28309));
    SB_LUT4 add_2307_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n28307), 
            .O(n6049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_4 (.CI(n28307), .I0(n2182), .I1(n98), .CO(n28308));
    SB_LUT4 add_2307_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n28306), 
            .O(n6050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_3 (.CI(n28306), .I0(n2183), .I1(n99), .CO(n28307));
    SB_LUT4 add_2307_2_lut (.I0(GND_net), .I1(n663), .I2(n558), .I3(VCC_net), 
            .O(n6051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2307_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2307_2 (.CI(VCC_net), .I0(n663), .I1(n558), .CO(n28306));
    SB_LUT4 add_2306_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n28305), 
            .O(n6017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2306_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n28304), 
            .O(n6018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_16 (.CI(n28304), .I0(n2070), .I1(n86), .CO(n28305));
    SB_LUT4 add_2306_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n28303), 
            .O(n6019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_15 (.CI(n28303), .I0(n2071), .I1(n87), .CO(n28304));
    SB_LUT4 add_2306_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n28302), 
            .O(n6020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_14 (.CI(n28302), .I0(n2072), .I1(n88), .CO(n28303));
    SB_LUT4 add_2306_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n28301), 
            .O(n6021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_13 (.CI(n28301), .I0(n2073), .I1(n89), .CO(n28302));
    SB_LUT4 add_2306_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n28300), 
            .O(n6022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_12 (.CI(n28300), .I0(n2074), .I1(n90), .CO(n28301));
    SB_LUT4 add_2306_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n28299), 
            .O(n6023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_11 (.CI(n28299), .I0(n2075), .I1(n91), .CO(n28300));
    SB_LUT4 add_2306_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n28298), 
            .O(n6024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_10 (.CI(n28298), .I0(n2076), .I1(n92), .CO(n28299));
    SB_LUT4 add_2306_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n28297), 
            .O(n6025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_9 (.CI(n28297), .I0(n2077), .I1(n93), .CO(n28298));
    SB_LUT4 add_2306_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n28296), 
            .O(n6026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_8 (.CI(n28296), .I0(n2078), .I1(n94), .CO(n28297));
    SB_LUT4 add_2306_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n28295), 
            .O(n6027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_7 (.CI(n28295), .I0(n2079), .I1(n95), .CO(n28296));
    SB_LUT4 add_2306_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n28294), 
            .O(n6028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_6 (.CI(n28294), .I0(n2080), .I1(n96), .CO(n28295));
    SB_LUT4 add_2306_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n28293), 
            .O(n6029)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_5 (.CI(n28293), .I0(n2081), .I1(n97), .CO(n28294));
    SB_LUT4 add_2306_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n28292), 
            .O(n6030)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_4 (.CI(n28292), .I0(n2082), .I1(n98), .CO(n28293));
    SB_LUT4 add_2306_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n28291), 
            .O(n6031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_3 (.CI(n28291), .I0(n2083), .I1(n99), .CO(n28292));
    SB_LUT4 add_2306_2_lut (.I0(GND_net), .I1(n662), .I2(n558), .I3(VCC_net), 
            .O(n6032)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2306_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2306_2 (.CI(VCC_net), .I0(n662), .I1(n558), .CO(n28291));
    SB_LUT4 add_2305_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n28290), 
            .O(n6000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2305_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n28289), 
            .O(n6001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_15 (.CI(n28289), .I0(n1968), .I1(n87), .CO(n28290));
    SB_LUT4 add_2305_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n28288), 
            .O(n6002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_14 (.CI(n28288), .I0(n1969), .I1(n88), .CO(n28289));
    SB_LUT4 i22_3_lut_adj_1844 (.I0(bit_ctr[29]), .I1(n40252), .I2(n4442), 
            .I3(GND_net), .O(n33493));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1844.LUT_INIT = 16'hacac;
    SB_LUT4 i12866_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17595));   // verilog/coms.v(126[12] 292[6])
    defparam i12866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12867_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17596));   // verilog/coms.v(126[12] 292[6])
    defparam i12867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1845 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1846 (.I0(n2848), .I1(n2853), .I2(n2851), .I3(n22_adj_4703), 
            .O(n37));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 i12868_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17597));   // verilog/coms.v(126[12] 292[6])
    defparam i12868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2305_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n28287), 
            .O(n6003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12869_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17598));   // verilog/coms.v(126[12] 292[6])
    defparam i12869_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF communication_counter_1185__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY add_2305_13 (.CI(n28287), .I0(n1970), .I1(n89), .CO(n28288));
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1554_adj_4850), .I2(GND_net), 
            .I3(n28985), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12870_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17599));   // verilog/coms.v(126[12] 292[6])
    defparam i12870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12871_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17600));   // verilog/coms.v(126[12] 292[6])
    defparam i12871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12872_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17601));   // verilog/coms.v(126[12] 292[6])
    defparam i12872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2305_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n28286), 
            .O(n6004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_12 (.CI(n28286), .I0(n1971), .I1(n90), .CO(n28287));
    SB_LUT4 add_2305_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n28285), 
            .O(n6005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_11 (.CI(n28285), .I0(n1972), .I1(n91), .CO(n28286));
    SB_LUT4 add_2305_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n28284), 
            .O(n6006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_10 (.CI(n28284), .I0(n1973), .I1(n92), .CO(n28285));
    SB_LUT4 add_2305_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n28283), 
            .O(n6007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_9 (.CI(n28283), .I0(n1974), .I1(n93), .CO(n28284));
    SB_LUT4 add_2305_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n28282), 
            .O(n6008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_8 (.CI(n28282), .I0(n1975), .I1(n94), .CO(n28283));
    SB_LUT4 add_2305_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n28281), 
            .O(n6009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_7 (.CI(n28281), .I0(n1976), .I1(n95), .CO(n28282));
    SB_LUT4 add_2305_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n28280), 
            .O(n6010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_6 (.CI(n28280), .I0(n1977), .I1(n96), .CO(n28281));
    SB_LUT4 add_2305_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n28279), 
            .O(n6011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_5 (.CI(n28279), .I0(n1978), .I1(n97), .CO(n28280));
    SB_LUT4 add_2305_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n28278), 
            .O(n6012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_4 (.CI(n28278), .I0(n1979), .I1(n98), .CO(n28279));
    SB_LUT4 add_2305_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n28277), 
            .O(n6013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_3 (.CI(n28277), .I0(n1980), .I1(n99), .CO(n28278));
    SB_LUT4 add_2305_2_lut (.I0(GND_net), .I1(n661), .I2(n558), .I3(VCC_net), 
            .O(n6014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2305_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2305_2 (.CI(VCC_net), .I0(n661), .I1(n558), .CO(n28277));
    SB_LUT4 add_2304_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n28276), 
            .O(n5984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2304_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n28275), 
            .O(n5985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_14 (.CI(n28275), .I0(n1863), .I1(n88), .CO(n28276));
    SB_LUT4 add_2304_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n28274), 
            .O(n5986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_13 (.CI(n28274), .I0(n1864), .I1(n89), .CO(n28275));
    SB_LUT4 add_2304_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n28273), 
            .O(n5987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_12 (.CI(n28273), .I0(n1865), .I1(n90), .CO(n28274));
    SB_LUT4 add_2304_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n28272), 
            .O(n5988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_11 (.CI(n28272), .I0(n1866), .I1(n91), .CO(n28273));
    SB_LUT4 add_2304_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n28271), 
            .O(n5989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_10 (.CI(n28271), .I0(n1867), .I1(n92), .CO(n28272));
    SB_LUT4 add_2304_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n28270), 
            .O(n5990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_9 (.CI(n28270), .I0(n1868), .I1(n93), .CO(n28271));
    SB_LUT4 add_2304_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n28269), 
            .O(n5991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_8 (.CI(n28269), .I0(n1869), .I1(n94), .CO(n28270));
    SB_LUT4 add_2304_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n28268), 
            .O(n5992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_7 (.CI(n28268), .I0(n1870), .I1(n95), .CO(n28269));
    SB_LUT4 add_2304_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n28267), 
            .O(n5993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_6 (.CI(n28267), .I0(n1871), .I1(n96), .CO(n28268));
    SB_LUT4 add_2304_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n28266), 
            .O(n5994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_5 (.CI(n28266), .I0(n1872), .I1(n97), .CO(n28267));
    SB_LUT4 add_2304_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n28265), 
            .O(n5995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_4 (.CI(n28265), .I0(n1873), .I1(n98), .CO(n28266));
    SB_LUT4 add_2304_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n28264), 
            .O(n5996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_3 (.CI(n28264), .I0(n1874), .I1(n99), .CO(n28265));
    SB_LUT4 add_2304_2_lut (.I0(GND_net), .I1(n660), .I2(n558), .I3(VCC_net), 
            .O(n5997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2304_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2304_2 (.CI(VCC_net), .I0(n660), .I1(n558), .CO(n28264));
    SB_LUT4 add_2303_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n28263), 
            .O(n5969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2303_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n28262), 
            .O(n5970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_13 (.CI(n28262), .I0(n1755), .I1(n89), .CO(n28263));
    SB_LUT4 add_2303_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n28261), 
            .O(n5971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_12 (.CI(n28261), .I0(n1756), .I1(n90), .CO(n28262));
    SB_LUT4 add_2303_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n28260), 
            .O(n5972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_11 (.CI(n28260), .I0(n1757), .I1(n91), .CO(n28261));
    SB_LUT4 add_2303_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n28259), 
            .O(n5973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_10 (.CI(n28259), .I0(n1758), .I1(n92), .CO(n28260));
    SB_LUT4 add_2303_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n28258), 
            .O(n5974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_9 (.CI(n28258), .I0(n1759), .I1(n93), .CO(n28259));
    SB_LUT4 add_2303_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n28257), 
            .O(n5975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_8 (.CI(n28257), .I0(n1760), .I1(n94), .CO(n28258));
    SB_LUT4 add_2303_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n28256), 
            .O(n5976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_7 (.CI(n28256), .I0(n1761), .I1(n95), .CO(n28257));
    SB_LUT4 add_2303_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n28255), 
            .O(n5977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_6 (.CI(n28255), .I0(n1762), .I1(n96), .CO(n28256));
    SB_LUT4 add_2303_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n28254), 
            .O(n5978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_5 (.CI(n28254), .I0(n1763), .I1(n97), .CO(n28255));
    SB_LUT4 add_2303_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n28253), 
            .O(n5979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_4 (.CI(n28253), .I0(n1764), .I1(n98), .CO(n28254));
    SB_LUT4 add_2303_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n28252), 
            .O(n5980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_3 (.CI(n28252), .I0(n1765), .I1(n99), .CO(n28253));
    SB_LUT4 add_2303_2_lut (.I0(GND_net), .I1(n659), .I2(n558), .I3(VCC_net), 
            .O(n5981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2303_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2303_2 (.CI(VCC_net), .I0(n659), .I1(n558), .CO(n28252));
    SB_LUT4 add_2302_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n28251), 
            .O(n5955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2302_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n28250), 
            .O(n5956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_12 (.CI(n28250), .I0(n1644), .I1(n90), .CO(n28251));
    SB_LUT4 add_2302_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n28249), 
            .O(n5957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12873_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17602));   // verilog/coms.v(126[12] 292[6])
    defparam i12873_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2302_11 (.CI(n28249), .I0(n1645), .I1(n91), .CO(n28250));
    SB_LUT4 add_2302_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n28248), 
            .O(n5958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_23_lut (.I0(n2638_adj_4855), .I1(n2638_adj_4855), 
            .I2(n2669), .I3(n28795), .O(n2737)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2302_10 (.CI(n28248), .I0(n1646), .I1(n92), .CO(n28249));
    SB_CARRY rem_4_add_1787_23 (.CI(n28795), .I0(n2638_adj_4855), .I1(n2669), 
            .CO(n28796));
    SB_LUT4 i12874_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17603));   // verilog/coms.v(126[12] 292[6])
    defparam i12874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2302_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n28247), 
            .O(n5959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12875_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17604));   // verilog/coms.v(126[12] 292[6])
    defparam i12875_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2302_9 (.CI(n28247), .I0(n1647), .I1(n93), .CO(n28248));
    SB_LUT4 i12612_4_lut (.I0(n17180), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n17052), .O(n17341));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12612_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 add_2302_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n28246), 
            .O(n5960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_8 (.CI(n28246), .I0(n1648), .I1(n94), .CO(n28247));
    SB_LUT4 add_2302_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n28245), 
            .O(n5961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_7 (.CI(n28245), .I0(n1649), .I1(n95), .CO(n28246));
    SB_LUT4 i22_3_lut_adj_1847 (.I0(bit_ctr[31]), .I1(n40254), .I2(n4442), 
            .I3(GND_net), .O(n33497));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1847.LUT_INIT = 16'hacac;
    SB_LUT4 add_2302_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n28244), 
            .O(n5962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_6 (.CI(n28244), .I0(n1650), .I1(n96), .CO(n28245));
    SB_LUT4 add_2302_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n28243), 
            .O(n5963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_5 (.CI(n28243), .I0(n1651), .I1(n97), .CO(n28244));
    SB_LUT4 div_46_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4924));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4923));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_3_lut_adj_1848 (.I0(n40277), .I1(byte_transmit_counter[1]), 
            .I2(n24391), .I3(GND_net), .O(n34177));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut_adj_1848.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4922));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1849 (.I0(n27), .I1(n36), .I2(n2845), .I3(n2846), 
            .O(n39));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i12609_4_lut (.I0(n17180), .I1(r_Bit_Index[2]), .I2(n4648), 
            .I3(n17052), .O(n17338));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12609_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i22_3_lut_adj_1850 (.I0(bit_ctr[14]), .I1(n40234), .I2(n4442), 
            .I3(GND_net), .O(n33457));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1850.LUT_INIT = 16'hacac;
    SB_LUT4 i20_4_lut_adj_1851 (.I0(n39), .I1(n37), .I2(n33), .I3(n34), 
            .O(n2867));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i20_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2302_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n28242), 
            .O(n5964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_4 (.CI(n28242), .I0(n1652), .I1(n98), .CO(n28243));
    SB_LUT4 add_2302_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n28241), 
            .O(n5965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_3 (.CI(n28241), .I0(n1653), .I1(n99), .CO(n28242));
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26_adj_4768), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2858));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2302_2_lut (.I0(GND_net), .I1(n658), .I2(n558), .I3(VCC_net), 
            .O(n5966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2302_2 (.CI(VCC_net), .I0(n658), .I1(n558), .CO(n28241));
    SB_LUT4 i22_3_lut_adj_1852 (.I0(bit_ctr[7]), .I1(n40233), .I2(n4442), 
            .I3(GND_net), .O(n33455));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1852.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4921));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1853 (.I0(blink), .I1(n15_adj_4714), .I2(GND_net), 
            .I3(GND_net), .O(blink_N_255));
    defparam i1_2_lut_adj_1853.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4920));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4919));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4918));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2301_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n28240), 
            .O(n5942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2301_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n28239), 
            .O(n5943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4917));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1050_7 (.CI(n28985), .I0(n1554_adj_4850), .I1(GND_net), 
            .CO(n28986));
    SB_LUT4 rem_4_add_1787_22_lut (.I0(n2639), .I1(n2639), .I2(n2669), 
            .I3(n28794), .O(n2738)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2301_11 (.CI(n28239), .I0(n1530), .I1(n91), .CO(n28240));
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4676));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4916));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4915));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2301_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n28238), 
            .O(n5944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_10 (.CI(n28238), .I0(n1531), .I1(n92), .CO(n28239));
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4675));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2301_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n28237), 
            .O(n5945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_9 (.CI(n28237), .I0(n1532), .I1(n93), .CO(n28238));
    SB_LUT4 add_2301_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n28236), 
            .O(n5946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2301_8 (.CI(n28236), .I0(n1533), .I1(n94), .CO(n28237));
    SB_LUT4 add_2301_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n28235), 
            .O(n5947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_7 (.CI(n28235), .I0(n1534), .I1(n95), .CO(n28236));
    SB_LUT4 div_46_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4914));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4674));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2301_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n28234), 
            .O(n5948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_6 (.CI(n28234), .I0(n1535), .I1(n96), .CO(n28235));
    SB_LUT4 div_46_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4913));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2301_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n28233), 
            .O(n5949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_5 (.CI(n28233), .I0(n1536), .I1(n97), .CO(n28234));
    SB_LUT4 add_2301_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n28232), 
            .O(n5950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2301_4 (.CI(n28232), .I0(n1537), .I1(n98), .CO(n28233));
    SB_LUT4 add_2301_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n28231), 
            .O(n5951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2301_3 (.CI(n28231), .I0(n1538), .I1(n99), .CO(n28232));
    SB_LUT4 add_2301_2_lut (.I0(GND_net), .I1(n657), .I2(n558), .I3(VCC_net), 
            .O(n5952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2301_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1185__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY add_2301_2 (.CI(VCC_net), .I0(n657), .I1(n558), .CO(n28231));
    SB_LUT4 add_2300_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n28230), 
            .O(n5930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n28984), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY rem_4_add_1787_22 (.CI(n28794), .I0(n2639), .I1(n2669), .CO(n28795));
    SB_LUT4 mux_70_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_106[0]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2300_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n28229), 
            .O(n5931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_21_lut (.I0(n2640), .I1(n2640), .I2(n2669), 
            .I3(n28793), .O(n2739)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mux_71_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_106[1]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut_adj_1854 (.I0(bit_ctr[6]), .I1(n40232), .I2(n4442), 
            .I3(GND_net), .O(n33453));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1854.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_106[2]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2300_10 (.CI(n28229), .I0(n1413), .I1(n92), .CO(n28230));
    SB_LUT4 add_2300_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n28228), 
            .O(n5932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2300_9 (.CI(n28228), .I0(n1414), .I1(n93), .CO(n28229));
    SB_LUT4 add_2300_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n28227), 
            .O(n5933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2300_8 (.CI(n28227), .I0(n1415), .I1(n94), .CO(n28228));
    SB_LUT4 add_2300_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n28226), 
            .O(n5934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_6 (.CI(n28984), .I0(n1555), .I1(GND_net), 
            .CO(n28985));
    SB_CARRY rem_4_add_1787_21 (.CI(n28793), .I0(n2640), .I1(n2669), .CO(n28794));
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n28983), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_20_lut (.I0(n2641), .I1(n2641), .I2(n2669), 
            .I3(n28792), .O(n2740)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2300_7 (.CI(n28226), .I0(n1416), .I1(n95), .CO(n28227));
    SB_CARRY rem_4_add_1050_5 (.CI(n28983), .I0(n1556), .I1(VCC_net), 
            .CO(n28984));
    SB_CARRY rem_4_add_1787_20 (.CI(n28792), .I0(n2641), .I1(n2669), .CO(n28793));
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n28982), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_19_lut (.I0(n2642_adj_4854), .I1(n2642_adj_4854), 
            .I2(n2669), .I3(n28791), .O(n2741)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2300_6_lut (.I0(GND_net), .I1(n1417_adj_4752), .I2(n96), 
            .I3(n28225), .O(n5935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2300_6 (.CI(n28225), .I0(n1417_adj_4752), .I1(n96), .CO(n28226));
    SB_CARRY rem_4_add_1050_4 (.CI(n28982), .I0(n1557), .I1(VCC_net), 
            .CO(n28983));
    SB_LUT4 add_2300_5_lut (.I0(GND_net), .I1(n1418_adj_4753), .I2(n97), 
            .I3(n28224), .O(n5936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_19 (.CI(n28791), .I0(n2642_adj_4854), .I1(n2669), 
            .CO(n28792));
    SB_LUT4 mux_71_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_2300_5 (.CI(n28224), .I0(n1418_adj_4753), .I1(n97), .CO(n28225));
    SB_LUT4 mux_70_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_106[3]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(n28981), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2300_4_lut (.I0(GND_net), .I1(n1419_adj_4754), .I2(n98), 
            .I3(n28223), .O(n5937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_18_lut (.I0(n2643_adj_4853), .I1(n2643_adj_4853), 
            .I2(n2669), .I3(n28790), .O(n2742)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2300_4 (.CI(n28223), .I0(n1419_adj_4754), .I1(n98), .CO(n28224));
    SB_LUT4 add_2300_3_lut (.I0(GND_net), .I1(n1420_adj_4755), .I2(n99), 
            .I3(n28222), .O(n5938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2300_3 (.CI(n28222), .I0(n1420_adj_4755), .I1(n99), .CO(n28223));
    SB_CARRY rem_4_add_1050_3 (.CI(n28981), .I0(n1558), .I1(GND_net), 
            .CO(n28982));
    SB_LUT4 mux_71_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY rem_4_add_1787_18 (.CI(n28790), .I0(n2643_adj_4853), .I1(n2669), 
            .CO(n28791));
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1658), .I1(VCC_net), 
            .CO(n28981));
    SB_LUT4 rem_4_add_1787_17_lut (.I0(n2644), .I1(n2644), .I2(n2669), 
            .I3(n28789), .O(n2743)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2300_2_lut (.I0(GND_net), .I1(n656), .I2(n558), .I3(VCC_net), 
            .O(n5939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2300_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_10_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n28980), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_70_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_106[4]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_17 (.CI(n28789), .I0(n2644), .I1(n2669), .CO(n28790));
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n28979), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_16_lut (.I0(n2645), .I1(n2645), .I2(n2669), 
            .I3(n28788), .O(n2744)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_2300_2 (.CI(VCC_net), .I0(n656), .I1(n558), .CO(n28222));
    SB_LUT4 add_2299_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n28221), 
            .O(n5919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2299_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n28220), 
            .O(n5920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_9 (.CI(n28220), .I0(n1293), .I1(n93), .CO(n28221));
    SB_CARRY rem_4_add_849_9 (.CI(n28979), .I0(n1251), .I1(VCC_net), .CO(n28980));
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n28978), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_16 (.CI(n28788), .I0(n2645), .I1(n2669), .CO(n28789));
    SB_LUT4 add_2299_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n28219), 
            .O(n5921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_8 (.CI(n28219), .I0(n1294), .I1(n94), .CO(n28220));
    SB_LUT4 add_2299_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n28218), 
            .O(n5922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_7 (.CI(n28218), .I0(n1295), .I1(n95), .CO(n28219));
    SB_LUT4 add_2299_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n28217), 
            .O(n5923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_15_lut (.I0(n2646), .I1(n2646), .I2(n2669), 
            .I3(n28787), .O(n2745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut (.I0(n852), .I1(n6_adj_5304), .I2(n746), .I3(GND_net), 
            .O(n884));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY add_2299_6 (.CI(n28217), .I0(n1296), .I1(n96), .CO(n28218));
    SB_LUT4 add_2299_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n28216), 
            .O(n5924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_5 (.CI(n28216), .I0(n1297), .I1(n97), .CO(n28217));
    SB_LUT4 add_2299_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n28215), 
            .O(n5925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_8 (.CI(n28978), .I0(n1252), .I1(VCC_net), .CO(n28979));
    SB_CARRY rem_4_add_1787_15 (.CI(n28787), .I0(n2646), .I1(n2669), .CO(n28788));
    SB_CARRY add_2299_4 (.CI(n28215), .I0(n1298), .I1(n98), .CO(n28216));
    SB_LUT4 rem_4_add_1787_14_lut (.I0(n2647), .I1(n2647), .I2(n2669), 
            .I3(n28786), .O(n2746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n28977), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_14 (.CI(n28786), .I0(n2647), .I1(n2669), .CO(n28787));
    SB_LUT4 rem_4_add_1787_13_lut (.I0(n2648), .I1(n2648), .I2(n2669), 
            .I3(n28785), .O(n2747)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_849_7 (.CI(n28977), .I0(n1253), .I1(VCC_net), .CO(n28978));
    SB_LUT4 i28526_2_lut_3_lut (.I0(n852), .I1(n6_adj_5304), .I2(n746), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i28526_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_CARRY rem_4_add_1787_13 (.CI(n28785), .I0(n2648), .I1(n2669), .CO(n28786));
    SB_LUT4 add_2299_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n28214), 
            .O(n5926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_3 (.CI(n28214), .I0(n1299), .I1(n99), .CO(n28215));
    SB_LUT4 add_2299_2_lut (.I0(GND_net), .I1(n655), .I2(n558), .I3(VCC_net), 
            .O(n5927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2299_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2299_2 (.CI(VCC_net), .I0(n655), .I1(n558), .CO(n28214));
    SB_LUT4 add_2298_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n28213), 
            .O(n5909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n28976), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_12_lut (.I0(n2649), .I1(n2649), .I2(n2669), 
            .I3(n28784), .O(n2748)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2298_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n28212), 
            .O(n5910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_12 (.CI(n28784), .I0(n2649), .I1(n2669), .CO(n28785));
    SB_CARRY add_2298_8 (.CI(n28212), .I0(n1170), .I1(n94), .CO(n28213));
    SB_LUT4 add_2298_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n28211), 
            .O(n5911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2298_7 (.CI(n28211), .I0(n1171), .I1(n95), .CO(n28212));
    SB_LUT4 add_2298_6_lut (.I0(GND_net), .I1(n1172_adj_4751), .I2(n96), 
            .I3(n28210), .O(n5912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2298_6 (.CI(n28210), .I0(n1172_adj_4751), .I1(n96), .CO(n28211));
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_5272), .I3(n29821), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_5273), .I3(n29820), .O(n3_adj_4832)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n29820), .I0(GND_net), .I1(n3_adj_5273), 
            .CO(n29821));
    SB_LUT4 add_2298_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n28209), 
            .O(n5913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_5274), .I3(n29819), .O(n4_adj_4831)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n29819), .I0(GND_net), .I1(n4_adj_5274), 
            .CO(n29820));
    SB_CARRY add_2298_5 (.CI(n28209), .I0(n1173), .I1(n97), .CO(n28210));
    SB_LUT4 add_2298_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n28208), 
            .O(n5914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_5275), .I3(n29818), .O(n5_adj_4830)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n29818), .I0(GND_net), .I1(n5_adj_5275), 
            .CO(n29819));
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_5276), .I3(n29817), .O(n6_adj_4829)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n29817), .I0(GND_net), .I1(n6_adj_5276), 
            .CO(n29818));
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_5277), .I3(n29816), .O(n7_adj_4828)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n29816), .I0(GND_net), .I1(n7_adj_5277), 
            .CO(n29817));
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_5278), .I3(n29815), .O(n8_adj_4827)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1185__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1185__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY add_2298_4 (.CI(n28208), .I0(n1174), .I1(n98), .CO(n28209));
    SB_LUT4 add_2298_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n28207), 
            .O(n5915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2298_3 (.CI(n28207), .I0(n1175), .I1(n99), .CO(n28208));
    SB_LUT4 add_2298_2_lut (.I0(GND_net), .I1(n654), .I2(n558), .I3(VCC_net), 
            .O(n5916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2298_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2298_2 (.CI(VCC_net), .I0(n654), .I1(n558), .CO(n28207));
    SB_LUT4 add_2297_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n28206), 
            .O(n5900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2297_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n28205), 
            .O(n5901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_7 (.CI(n28205), .I0(n1044), .I1(n95), .CO(n28206));
    SB_LUT4 add_2297_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n28204), 
            .O(n5902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_6 (.CI(n28204), .I0(n1045), .I1(n96), .CO(n28205));
    SB_LUT4 add_2297_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n28203), 
            .O(n5903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n29815), .I0(GND_net), .I1(n8_adj_5278), 
            .CO(n29816));
    SB_CARRY add_2297_5 (.CI(n28203), .I0(n1046), .I1(n97), .CO(n28204));
    SB_LUT4 add_2297_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n28202), 
            .O(n5904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_5279), .I3(n29814), .O(n9_adj_4826)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_4 (.CI(n28202), .I0(n1047), .I1(n98), .CO(n28203));
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n29814), .I0(GND_net), .I1(n9_adj_5279), 
            .CO(n29815));
    SB_CARRY rem_4_add_849_6 (.CI(n28976), .I0(n1254), .I1(GND_net), .CO(n28977));
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_5280), .I3(n29813), .O(n10_adj_4825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_11_lut (.I0(n2650), .I1(n2650), .I2(n2669), 
            .I3(n28783), .O(n2749)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_2297_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n28201), 
            .O(n5905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n29813), .I0(GND_net), .I1(n10_adj_5280), 
            .CO(n29814));
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_5281), .I3(n29812), .O(n11_adj_4824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2297_3 (.CI(n28201), .I0(n1048), .I1(n99), .CO(n28202));
    SB_LUT4 add_2297_2_lut (.I0(GND_net), .I1(n653), .I2(n558), .I3(VCC_net), 
            .O(n5906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2297_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n29812), .I0(GND_net), .I1(n11_adj_5281), 
            .CO(n29813));
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_5282), .I3(n29811), .O(n12_adj_4782)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n29811), .I0(GND_net), .I1(n12_adj_5282), 
            .CO(n29812));
    SB_CARRY add_2297_2 (.CI(VCC_net), .I0(n653), .I1(n558), .CO(n28201));
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n28975), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n28783), .I0(n2650), .I1(n2669), .CO(n28784));
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_5283), .I3(n29810), .O(n13_adj_4781)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n29810), .I0(GND_net), .I1(n13_adj_5283), 
            .CO(n29811));
    SB_LUT4 add_2296_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n28200), 
            .O(n5892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_5284), .I3(n29809), .O(n14_adj_4780)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n28199), 
            .O(n5893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_5 (.CI(n28975), .I0(n1255), .I1(GND_net), .CO(n28976));
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n29809), .I0(GND_net), .I1(n14_adj_5284), 
            .CO(n29810));
    SB_CARRY add_2296_6 (.CI(n28199), .I0(n915), .I1(n96), .CO(n28200));
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_5285), .I3(n29808), .O(n15_adj_4779)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n28198), 
            .O(n5894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2296_5 (.CI(n28198), .I0(n916), .I1(n97), .CO(n28199));
    SB_LUT4 add_2296_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n28197), 
            .O(n5895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n29808), .I0(GND_net), .I1(n15_adj_5285), 
            .CO(n29809));
    SB_CARRY add_2296_4 (.CI(n28197), .I0(n917), .I1(n98), .CO(n28198));
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_5286), .I3(n29807), .O(n16_adj_4778)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n29807), .I0(GND_net), .I1(n16_adj_5286), 
            .CO(n29808));
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_5287), .I3(n29806), .O(n17_adj_4777)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n28196), 
            .O(n5896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n29806), .I0(GND_net), .I1(n17_adj_5287), 
            .CO(n29807));
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_5288), .I3(n29805), .O(n18_adj_4776)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n29805), .I0(GND_net), .I1(n18_adj_5288), 
            .CO(n29806));
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_5289), .I3(n29804), .O(n19_adj_4775)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n29804), .I0(GND_net), .I1(n19_adj_5289), 
            .CO(n29805));
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_5290), .I3(n29803), .O(n20_adj_4774)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n29803), .I0(GND_net), .I1(n20_adj_5290), 
            .CO(n29804));
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_5291), .I3(n29802), .O(n21_adj_4773)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n29802), .I0(GND_net), .I1(n21_adj_5291), 
            .CO(n29803));
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_5292), .I3(n29801), .O(n22_adj_4772)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n29801), .I0(GND_net), .I1(n22_adj_5292), 
            .CO(n29802));
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_5293), .I3(n29800), .O(n23_adj_4771)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n29800), .I0(GND_net), .I1(n23_adj_5293), 
            .CO(n29801));
    SB_CARRY add_2296_3 (.CI(n28196), .I0(n918), .I1(n99), .CO(n28197));
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_5294), .I3(n29799), .O(n24_adj_4770)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n29799), .I0(GND_net), .I1(n24_adj_5294), 
            .CO(n29800));
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_5295), .I3(n29798), .O(n25_adj_4769)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2296_2_lut (.I0(GND_net), .I1(n652), .I2(n558), .I3(VCC_net), 
            .O(n5897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2296_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n29798), .I0(GND_net), .I1(n25_adj_5295), 
            .CO(n29799));
    SB_CARRY add_2296_2 (.CI(VCC_net), .I0(n652), .I1(n558), .CO(n28196));
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_5296), .I3(n29797), .O(n26_adj_4768)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n29797), .I0(GND_net), .I1(n26_adj_5296), 
            .CO(n29798));
    SB_LUT4 rem_4_add_1787_10_lut (.I0(n2651), .I1(n2651), .I2(n2669), 
            .I3(n28782), .O(n2750)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_5297), .I3(n29796), .O(n27_adj_4767)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n28974), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_4 (.CI(n28974), .I0(n1256), .I1(VCC_net), .CO(n28975));
    SB_CARRY rem_4_add_1787_10 (.CI(n28782), .I0(n2651), .I1(n2669), .CO(n28783));
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n29796), .I0(GND_net), .I1(n27_adj_5297), 
            .CO(n29797));
    SB_LUT4 rem_4_add_1787_9_lut (.I0(n2652), .I1(n2652), .I2(n2669), 
            .I3(n28781), .O(n2751)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_5298), .I3(n29795), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_9 (.CI(n28781), .I0(n2652), .I1(n2669), .CO(n28782));
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n29795), .I0(GND_net), .I1(n28_adj_5298), 
            .CO(n29796));
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n28973), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_8_lut (.I0(n2653), .I1(n2653), .I2(n2669), 
            .I3(n28780), .O(n2752)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_5299), .I3(n29794), .O(n29_adj_4766)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_8 (.CI(n28780), .I0(n2653), .I1(n2669), .CO(n28781));
    SB_CARRY rem_4_add_849_3 (.CI(n28973), .I0(n1257), .I1(VCC_net), .CO(n28974));
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n29794), .I0(GND_net), .I1(n29_adj_5299), 
            .CO(n29795));
    SB_LUT4 rem_4_add_849_2_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(VCC_net), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_7_lut (.I0(n2654), .I1(n2654), .I2(n43156), 
            .I3(n28779), .O(n2753)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_5300), .I3(n29793), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n29793), .I0(GND_net), .I1(n30_adj_5300), 
            .CO(n29794));
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1258), .I1(GND_net), 
            .CO(n28973));
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4839), .I2(VCC_net), 
            .I3(n28972), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_5301), .I3(n29792), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_7 (.CI(n28779), .I0(n2654), .I1(n43156), .CO(n28780));
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4840), .I2(VCC_net), 
            .I3(n28971), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n29792), .I0(GND_net), .I1(n31_adj_5301), 
            .CO(n29793));
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_5302), .I3(n29791), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n29791), .I0(GND_net), .I1(n32_adj_5302), 
            .CO(n29792));
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_5303), .I3(VCC_net), .O(n33_adj_4765)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_5303), 
            .CO(n29791));
    SB_CARRY rem_4_add_1117_14 (.CI(n28971), .I0(n1647_adj_4840), .I1(VCC_net), 
            .CO(n28972));
    SB_LUT4 rem_4_add_1787_6_lut (.I0(n2655), .I1(n2655), .I2(n43156), 
            .I3(n28778), .O(n2754)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1787_6 (.CI(n28778), .I0(n2655), .I1(n43156), .CO(n28779));
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4841), .I2(VCC_net), 
            .I3(n28970), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_5_lut (.I0(n2656), .I1(n2656), .I2(n2669), 
            .I3(n28777), .O(n2755)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1787_5 (.CI(n28777), .I0(n2656), .I1(n2669), .CO(n28778));
    SB_LUT4 rem_4_add_715_8_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n28190), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1117_13 (.CI(n28970), .I0(n1648_adj_4841), .I1(VCC_net), 
            .CO(n28971));
    SB_LUT4 rem_4_add_1787_4_lut (.I0(n2657), .I1(n2657), .I2(n2669), 
            .I3(n28776), .O(n2756)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4842), .I2(VCC_net), 
            .I3(n28969), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_23 (.CI(n28647), .I0(n3038), .I1(VCC_net), 
            .CO(n28648));
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n28189), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_7 (.CI(n28189), .I0(n1053), .I1(VCC_net), .CO(n28190));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n28188), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_4 (.CI(n28776), .I0(n2657), .I1(n2669), .CO(n28777));
    SB_CARRY rem_4_add_715_6 (.CI(n28188), .I0(n1054), .I1(GND_net), .CO(n28189));
    SB_CARRY rem_4_add_1117_12 (.CI(n28969), .I0(n1649_adj_4842), .I1(VCC_net), 
            .CO(n28970));
    SB_LUT4 rem_4_add_1787_3_lut (.I0(n2658), .I1(n2658), .I2(n43156), 
            .I3(n28775), .O(n2757)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n28187), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_3 (.CI(n28775), .I0(n2658), .I1(n43156), .CO(n28776));
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4844), .I2(VCC_net), 
            .I3(n28968), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_5 (.CI(n28187), .I0(n1055), .I1(GND_net), .CO(n28188));
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2758), .I1(VCC_net), 
            .CO(n28775));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n28774), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n28186), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_11 (.CI(n28968), .I0(n1650_adj_4844), .I1(VCC_net), 
            .CO(n28969));
    SB_CARRY rem_4_add_715_4 (.CI(n28186), .I0(n1056), .I1(VCC_net), .CO(n28187));
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n28185), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4845), .I2(VCC_net), 
            .I3(n28967), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_10 (.CI(n28967), .I0(n1651_adj_4845), .I1(VCC_net), 
            .CO(n28968));
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n28773), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_3 (.CI(n28185), .I0(n1057), .I1(VCC_net), .CO(n28186));
    SB_LUT4 rem_4_add_715_2_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(VCC_net), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1058), .I1(GND_net), 
            .CO(n28185));
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4846), .I2(VCC_net), 
            .I3(n28966), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_9 (.CI(n28966), .I0(n1652_adj_4846), .I1(VCC_net), 
            .CO(n28967));
    SB_CARRY rem_4_add_1854_25 (.CI(n28773), .I0(n2736), .I1(VCC_net), 
            .CO(n28774));
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4847), .I2(VCC_net), 
            .I3(n28965), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_8 (.CI(n28965), .I0(n1653_adj_4847), .I1(VCC_net), 
            .CO(n28966));
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n28772), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_24 (.CI(n28772), .I0(n2737), .I1(VCC_net), 
            .CO(n28773));
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n28964), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n28771), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_7 (.CI(n28964), .I0(n1654), .I1(GND_net), 
            .CO(n28965));
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n28963), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_23 (.CI(n28771), .I0(n2738), .I1(VCC_net), 
            .CO(n28772));
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n28770), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_22 (.CI(n28770), .I0(n2739), .I1(VCC_net), 
            .CO(n28771));
    SB_CARRY rem_4_add_1117_6 (.CI(n28963), .I0(n1655), .I1(GND_net), 
            .CO(n28964));
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n28769), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_21 (.CI(n28769), .I0(n2740), .I1(VCC_net), 
            .CO(n28770));
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n28962), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n28768), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_20 (.CI(n28768), .I0(n2741), .I1(VCC_net), 
            .CO(n28769));
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n28767), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_5 (.CI(n28962), .I0(n1656), .I1(VCC_net), 
            .CO(n28963));
    SB_CARRY rem_4_add_1854_19 (.CI(n28767), .I0(n2742), .I1(VCC_net), 
            .CO(n28768));
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n28961), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n28766), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_18 (.CI(n28766), .I0(n2743), .I1(VCC_net), 
            .CO(n28767));
    SB_CARRY rem_4_add_1117_4 (.CI(n28961), .I0(n1657), .I1(VCC_net), 
            .CO(n28962));
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n28765), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_17 (.CI(n28765), .I0(n2744), .I1(VCC_net), 
            .CO(n28766));
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n28960), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n28764), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_3 (.CI(n28960), .I0(n1658), .I1(GND_net), 
            .CO(n28961));
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4838), .I1(VCC_net), 
            .CO(n28960));
    SB_LUT4 rem_4_add_1184_16_lut (.I0(n1778_adj_4833), .I1(n1745), .I2(VCC_net), 
            .I3(n28959), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1854_16 (.CI(n28764), .I0(n2745), .I1(VCC_net), 
            .CO(n28765));
    SB_LUT4 rem_4_add_1184_15_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n28958), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n28763), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_15 (.CI(n28958), .I0(n1746), .I1(VCC_net), 
            .CO(n28959));
    SB_CARRY rem_4_add_1854_15 (.CI(n28763), .I0(n2746), .I1(VCC_net), 
            .CO(n28764));
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n28957), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n28762), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n28957), .I0(n1747), .I1(VCC_net), 
            .CO(n28958));
    SB_CARRY rem_4_add_1854_14 (.CI(n28762), .I0(n2747), .I1(VCC_net), 
            .CO(n28763));
    SB_LUT4 mux_71_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n28956), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n28761), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_13 (.CI(n28956), .I0(n1748), .I1(VCC_net), 
            .CO(n28957));
    SB_CARRY rem_4_add_1854_13 (.CI(n28761), .I0(n2748), .I1(VCC_net), 
            .CO(n28762));
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n28955), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n28760), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_12 (.CI(n28955), .I0(n1749), .I1(VCC_net), 
            .CO(n28956));
    SB_CARRY rem_4_add_1854_12 (.CI(n28760), .I0(n2749), .I1(VCC_net), 
            .CO(n28761));
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n28954), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n28759), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_11 (.CI(n28954), .I0(n1750), .I1(VCC_net), 
            .CO(n28955));
    SB_CARRY rem_4_add_1854_11 (.CI(n28759), .I0(n2750), .I1(VCC_net), 
            .CO(n28760));
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n28953), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n28758), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_10 (.CI(n28953), .I0(n1751), .I1(VCC_net), 
            .CO(n28954));
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n28952), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_10 (.CI(n28758), .I0(n2751), .I1(VCC_net), 
            .CO(n28759));
    SB_CARRY rem_4_add_1184_9 (.CI(n28952), .I0(n1752), .I1(VCC_net), 
            .CO(n28953));
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n28757), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n28951), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_9 (.CI(n28757), .I0(n2752), .I1(VCC_net), 
            .CO(n28758));
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n28756), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n28951), .I0(n1753), .I1(VCC_net), 
            .CO(n28952));
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1754_adj_4834), .I2(GND_net), 
            .I3(n28950), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_8 (.CI(n28756), .I0(n2753), .I1(VCC_net), 
            .CO(n28757));
    SB_LUT4 rem_4_add_782_9_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n28141), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n28140), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_8 (.CI(n28140), .I0(n1152), .I1(VCC_net), .CO(n28141));
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n28139), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_7 (.CI(n28950), .I0(n1754_adj_4834), .I1(GND_net), 
            .CO(n28951));
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n28755), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_7 (.CI(n28139), .I0(n1153), .I1(VCC_net), .CO(n28140));
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n28138), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_6 (.CI(n28138), .I0(n1154), .I1(GND_net), .CO(n28139));
    SB_CARRY rem_4_add_1854_7 (.CI(n28755), .I0(n2754), .I1(GND_net), 
            .CO(n28756));
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n28137), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1755_adj_4835), .I2(GND_net), 
            .I3(n28949), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n28754), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_6 (.CI(n28949), .I0(n1755_adj_4835), .I1(GND_net), 
            .CO(n28950));
    SB_CARRY rem_4_add_1854_6 (.CI(n28754), .I0(n2755), .I1(GND_net), 
            .CO(n28755));
    SB_CARRY rem_4_add_782_5 (.CI(n28137), .I0(n1155), .I1(GND_net), .CO(n28138));
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n28136), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_4 (.CI(n28136), .I0(n1156), .I1(VCC_net), .CO(n28137));
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n28135), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_3 (.CI(n28135), .I0(n1157), .I1(VCC_net), .CO(n28136));
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n28753), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_2_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(VCC_net), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1158), .I1(GND_net), 
            .CO(n28135));
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1756_adj_4836), .I2(VCC_net), 
            .I3(n28948), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_5 (.CI(n28753), .I0(n2756), .I1(VCC_net), 
            .CO(n28754));
    SB_CARRY rem_4_add_1184_5 (.CI(n28948), .I0(n1756_adj_4836), .I1(VCC_net), 
            .CO(n28949));
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n28752), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_4 (.CI(n28752), .I0(n2757), .I1(VCC_net), 
            .CO(n28753));
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1757_adj_4837), .I2(VCC_net), 
            .I3(n28947), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n28751), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_70_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_106[5]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_4 (.CI(n28947), .I0(n1757_adj_4837), .I1(VCC_net), 
            .CO(n28948));
    SB_CARRY rem_4_add_1854_3 (.CI(n28751), .I0(n2758), .I1(GND_net), 
            .CO(n28752));
    SB_LUT4 rem_4_add_648_7_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n27847), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n27846), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_6 (.CI(n27846), .I0(n954), .I1(GND_net), .CO(n27847));
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1758_adj_4838), .I2(GND_net), 
            .I3(n28946), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2858), .I1(VCC_net), 
            .CO(n28751));
    SB_LUT4 rem_4_add_1921_27_lut (.I0(n2867), .I1(n2834), .I2(VCC_net), 
            .I3(n28750), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_916_11_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n28125), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n28124), .O(n1417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n27845), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_10 (.CI(n28124), .I0(n1350), .I1(VCC_net), 
            .CO(n28125));
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n28123), .O(n1418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_9 (.CI(n28123), .I0(n1351), .I1(VCC_net), .CO(n28124));
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n28122), .O(n1419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_8 (.CI(n28122), .I0(n1352), .I1(VCC_net), .CO(n28123));
    SB_CARRY rem_4_add_1184_3 (.CI(n28946), .I0(n1758_adj_4838), .I1(GND_net), 
            .CO(n28947));
    SB_LUT4 rem_4_add_1921_26_lut (.I0(GND_net), .I1(n2835), .I2(VCC_net), 
            .I3(n28749), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_5 (.CI(n27845), .I0(n955), .I1(GND_net), .CO(n27846));
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n28121), .O(n1420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_7 (.CI(n28121), .I0(n1353), .I1(VCC_net), .CO(n28122));
    SB_LUT4 div_46_i1471_3_lut_3_lut (.I0(n2192), .I1(n6047), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n28120), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1855 (.I0(control_mode[0]), .I1(n15778), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4672));   // verilog/TinyFPGA_B.v(228[5:22])
    defparam i1_2_lut_3_lut_adj_1855.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n27844), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_6 (.CI(n28120), .I0(n1354), .I1(GND_net), .CO(n28121));
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n28119), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_5 (.CI(n28119), .I0(n1355), .I1(GND_net), .CO(n28120));
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n28118), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1856 (.I0(control_mode[0]), .I1(n15778), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(228[5:22])
    defparam i1_2_lut_3_lut_adj_1856.LUT_INIT = 16'hefef;
    SB_CARRY rem_4_add_916_4 (.CI(n28118), .I0(n1356), .I1(VCC_net), .CO(n28119));
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n28117), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_3 (.CI(n28117), .I0(n1357), .I1(VCC_net), .CO(n28118));
    SB_LUT4 rem_4_add_916_2_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(VCC_net), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1358), .I1(GND_net), 
            .CO(n28117));
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_229[23]), 
            .I2(n3_adj_4705), .I3(n28116), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_229[22]), 
            .I2(n3_adj_4705), .I3(n28115), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n28115), .I0(displacement_23__N_229[22]), 
            .I1(n3_adj_4705), .CO(n28116));
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1858), .I1(VCC_net), 
            .CO(n28946));
    SB_CARRY rem_4_add_1921_26 (.CI(n28749), .I0(n2835), .I1(VCC_net), 
            .CO(n28750));
    SB_CARRY rem_4_add_648_4 (.CI(n27844), .I0(n956), .I1(VCC_net), .CO(n27845));
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n27843), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_229[21]), 
            .I2(n3_adj_4705), .I3(n28114), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_17_lut (.I0(n1877), .I1(n1844), .I2(VCC_net), 
            .I3(n28945), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2836), .I2(VCC_net), 
            .I3(n28748), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n28114), .I0(displacement_23__N_229[21]), 
            .I1(n3_adj_4705), .CO(n28115));
    SB_LUT4 rem_4_add_1251_16_lut (.I0(GND_net), .I1(n1845), .I2(VCC_net), 
            .I3(n28944), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_229[20]), 
            .I2(n3_adj_4705), .I3(n28113), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n28113), .I0(displacement_23__N_229[20]), 
            .I1(n3_adj_4705), .CO(n28114));
    SB_CARRY rem_4_add_1921_25 (.CI(n28748), .I0(n2836), .I1(VCC_net), 
            .CO(n28749));
    SB_CARRY rem_4_add_648_3 (.CI(n27843), .I0(n957), .I1(VCC_net), .CO(n27844));
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2837), .I2(VCC_net), 
            .I3(n28747), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_16 (.CI(n28944), .I0(n1845), .I1(VCC_net), 
            .CO(n28945));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_229[19]), 
            .I2(n6_adj_4698), .I3(n28112), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_15_lut (.I0(GND_net), .I1(n1846), .I2(VCC_net), 
            .I3(n28943), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_24 (.CI(n28747), .I0(n2837), .I1(VCC_net), 
            .CO(n28748));
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n28112), .I0(displacement_23__N_229[19]), 
            .I1(n6_adj_4698), .CO(n28113));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_229[18]), 
            .I2(n7_adj_4697), .I3(n28111), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_2_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(VCC_net), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_15 (.CI(n28943), .I0(n1846), .I1(VCC_net), 
            .CO(n28944));
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2838), .I2(VCC_net), 
            .I3(n28746), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_14_lut (.I0(GND_net), .I1(n1847), .I2(VCC_net), 
            .I3(n28942), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_23 (.CI(n28746), .I0(n2838), .I1(VCC_net), 
            .CO(n28747));
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n28111), .I0(displacement_23__N_229[18]), 
            .I1(n7_adj_4697), .CO(n28112));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_229[17]), 
            .I2(n8_adj_4696), .I3(n28110), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n28110), .I0(displacement_23__N_229[17]), 
            .I1(n8_adj_4696), .CO(n28111));
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2839), .I2(VCC_net), 
            .I3(n28745), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_14 (.CI(n28942), .I0(n1847), .I1(VCC_net), 
            .CO(n28943));
    SB_CARRY rem_4_add_1921_22 (.CI(n28745), .I0(n2839), .I1(VCC_net), 
            .CO(n28746));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_229[16]), 
            .I2(n9_adj_4695), .I3(n28109), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n958), .I1(GND_net), .CO(n27843));
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n28109), .I0(displacement_23__N_229[16]), 
            .I1(n9_adj_4695), .CO(n28110));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_229[15]), 
            .I2(n10_adj_4694), .I3(n28108), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1459_3_lut_3_lut (.I0(n2192), .I1(n6035), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1251_13_lut (.I0(GND_net), .I1(n1848), .I2(VCC_net), 
            .I3(n28941), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n28744), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n28108), .I0(displacement_23__N_229[15]), 
            .I1(n10_adj_4694), .CO(n28109));
    SB_CARRY rem_4_add_1251_13 (.CI(n28941), .I0(n1848), .I1(VCC_net), 
            .CO(n28942));
    SB_LUT4 rem_4_add_1251_12_lut (.I0(GND_net), .I1(n1849), .I2(VCC_net), 
            .I3(n28940), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_21 (.CI(n28744), .I0(n2840), .I1(VCC_net), 
            .CO(n28745));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_229[14]), 
            .I2(n11_adj_4692), .I3(n28107), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n28107), .I0(displacement_23__N_229[14]), 
            .I1(n11_adj_4692), .CO(n28108));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_229[13]), 
            .I2(n12_adj_4737), .I3(n28106), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n28106), .I0(displacement_23__N_229[13]), 
            .I1(n12_adj_4737), .CO(n28107));
    SB_CARRY rem_4_add_1251_12 (.CI(n28940), .I0(n1849), .I1(VCC_net), 
            .CO(n28941));
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n28743), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_229[12]), 
            .I2(n13_adj_4738), .I3(n28105), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n28105), .I0(displacement_23__N_229[12]), 
            .I1(n13_adj_4738), .CO(n28106));
    SB_LUT4 rem_4_add_1251_11_lut (.I0(GND_net), .I1(n1850), .I2(VCC_net), 
            .I3(n28939), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_20 (.CI(n28743), .I0(n2841), .I1(VCC_net), 
            .CO(n28744));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_229[11]), 
            .I2(n14_adj_4739), .I3(n28104), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n28104), .I0(displacement_23__N_229[11]), 
            .I1(n14_adj_4739), .CO(n28105));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_229[10]), 
            .I2(n15_adj_4740), .I3(n28103), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n28742), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n28103), .I0(displacement_23__N_229[10]), 
            .I1(n15_adj_4740), .CO(n28104));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_229[9]), 
            .I2(n16_adj_4741), .I3(n28102), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n28102), .I0(displacement_23__N_229[9]), 
            .I1(n16_adj_4741), .CO(n28103));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_229[8]), 
            .I2(n17_adj_4742), .I3(n28101), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n28101), .I0(displacement_23__N_229[8]), 
            .I1(n17_adj_4742), .CO(n28102));
    SB_CARRY rem_4_add_1251_11 (.CI(n28939), .I0(n1850), .I1(VCC_net), 
            .CO(n28940));
    SB_CARRY rem_4_add_1921_19 (.CI(n28742), .I0(n2842), .I1(VCC_net), 
            .CO(n28743));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_229[7]), 
            .I2(n18_adj_4743), .I3(n28100), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n28100), .I0(displacement_23__N_229[7]), 
            .I1(n18_adj_4743), .CO(n28101));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_229[6]), 
            .I2(n19_adj_4744), .I3(n28099), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n28099), .I0(displacement_23__N_229[6]), 
            .I1(n19_adj_4744), .CO(n28100));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_229[5]), 
            .I2(n20_adj_4745), .I3(n28098), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27_adj_4767), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958_adj_4802));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n28098), .I0(displacement_23__N_229[5]), 
            .I1(n20_adj_4745), .CO(n28099));
    SB_LUT4 rem_4_add_1251_10_lut (.I0(GND_net), .I1(n1851), .I2(VCC_net), 
            .I3(n28938), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n28741), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_229[4]), 
            .I2(n21_adj_4746), .I3(n28097), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_10 (.CI(n28938), .I0(n1851), .I1(VCC_net), 
            .CO(n28939));
    SB_CARRY rem_4_add_1921_18 (.CI(n28741), .I0(n2843), .I1(VCC_net), 
            .CO(n28742));
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n28740), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n28097), .I0(displacement_23__N_229[4]), 
            .I1(n21_adj_4746), .CO(n28098));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_229[3]), 
            .I2(n22_adj_4747), .I3(n28096), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n28096), .I0(displacement_23__N_229[3]), 
            .I1(n22_adj_4747), .CO(n28097));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_229[2]), 
            .I2(n23_adj_4748), .I3(n28095), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n28095), .I0(displacement_23__N_229[2]), 
            .I1(n23_adj_4748), .CO(n28096));
    SB_LUT4 rem_4_add_1251_9_lut (.I0(GND_net), .I1(n1852), .I2(VCC_net), 
            .I3(n28937), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_17 (.CI(n28740), .I0(n2844), .I1(VCC_net), 
            .CO(n28741));
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_229[1]), 
            .I2(n24_adj_4749), .I3(n28094), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n28094), .I0(displacement_23__N_229[1]), 
            .I1(n24_adj_4749), .CO(n28095));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_229[0]), 
            .I2(n25_adj_4750), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_229[0]), 
            .I1(n25_adj_4750), .CO(n28094));
    SB_CARRY rem_4_add_1251_9 (.CI(n28937), .I0(n1852), .I1(VCC_net), 
            .CO(n28938));
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n28739), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_8_lut (.I0(GND_net), .I1(n1853), .I2(VCC_net), 
            .I3(n28936), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_16 (.CI(n28739), .I0(n2845), .I1(VCC_net), 
            .CO(n28740));
    SB_CARRY rem_4_add_1251_8 (.CI(n28936), .I0(n1853), .I1(VCC_net), 
            .CO(n28937));
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n28738), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_15 (.CI(n28738), .I0(n2846), .I1(VCC_net), 
            .CO(n28739));
    SB_LUT4 rem_4_add_1251_7_lut (.I0(GND_net), .I1(n1854), .I2(GND_net), 
            .I3(n28935), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n28737), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_7 (.CI(n28935), .I0(n1854), .I1(GND_net), 
            .CO(n28936));
    SB_CARRY rem_4_add_1921_14 (.CI(n28737), .I0(n2847), .I1(VCC_net), 
            .CO(n28738));
    SB_LUT4 rem_4_add_1251_6_lut (.I0(GND_net), .I1(n1855), .I2(GND_net), 
            .I3(n28934), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n28736), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1857 (.I0(bit_ctr[5]), .I1(n40231), .I2(n4442), 
            .I3(GND_net), .O(n33451));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1857.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1251_6 (.CI(n28934), .I0(n1855), .I1(GND_net), 
            .CO(n28935));
    SB_CARRY rem_4_add_1921_13 (.CI(n28736), .I0(n2848), .I1(VCC_net), 
            .CO(n28737));
    SB_LUT4 rem_4_add_1251_5_lut (.I0(GND_net), .I1(n1856), .I2(VCC_net), 
            .I3(n28933), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n28735), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_5 (.CI(n28933), .I0(n1856), .I1(VCC_net), 
            .CO(n28934));
    SB_CARRY rem_4_add_1921_12 (.CI(n28735), .I0(n2849), .I1(VCC_net), 
            .CO(n28736));
    SB_LUT4 mux_71_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 rem_4_add_1251_4_lut (.I0(GND_net), .I1(n1857), .I2(VCC_net), 
            .I3(n28932), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_4 (.CI(n28932), .I0(n1857), .I1(VCC_net), 
            .CO(n28933));
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n28734), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_11 (.CI(n28734), .I0(n2850), .I1(VCC_net), 
            .CO(n28735));
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n28733), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_3_lut (.I0(GND_net), .I1(n1858), .I2(GND_net), 
            .I3(n28931), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_10 (.CI(n28733), .I0(n2851), .I1(VCC_net), 
            .CO(n28734));
    SB_CARRY rem_4_add_1251_3 (.CI(n28931), .I0(n1858), .I1(GND_net), 
            .CO(n28932));
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n28732), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1958), .I1(VCC_net), 
            .CO(n28931));
    SB_LUT4 rem_4_add_1318_18_lut (.I0(n1976_adj_5033), .I1(n1943), .I2(VCC_net), 
            .I3(n28930), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1318_17_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n28929), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_17 (.CI(n28929), .I0(n1944), .I1(VCC_net), 
            .CO(n28930));
    SB_CARRY rem_4_add_1921_9 (.CI(n28732), .I0(n2852), .I1(VCC_net), 
            .CO(n28733));
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n28731), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY rem_4_add_1921_8 (.CI(n28731), .I0(n2853), .I1(VCC_net), 
            .CO(n28732));
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n28928), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n28730), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n28928), .I0(n1945), .I1(VCC_net), 
            .CO(n28929));
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n28927), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_7 (.CI(n28730), .I0(n2854), .I1(GND_net), 
            .CO(n28731));
    SB_CARRY rem_4_add_1318_15 (.CI(n28927), .I0(n1946), .I1(VCC_net), 
            .CO(n28928));
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n28926), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2855), .I2(GND_net), 
            .I3(n28729), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_14 (.CI(n28926), .I0(n1947), .I1(VCC_net), 
            .CO(n28927));
    SB_CARRY rem_4_add_1921_6 (.CI(n28729), .I0(n2855), .I1(GND_net), 
            .CO(n28730));
    SB_LUT4 i22_3_lut_adj_1858 (.I0(bit_ctr[13]), .I1(n40230), .I2(n4442), 
            .I3(GND_net), .O(n33445));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1858.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n28728), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_5 (.CI(n28728), .I0(n2856), .I1(VCC_net), 
            .CO(n28729));
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n28925), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2857), .I2(VCC_net), 
            .I3(n28727), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_4 (.CI(n28727), .I0(n2857), .I1(VCC_net), 
            .CO(n28728));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2858), .I2(GND_net), 
            .I3(n28726), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_3 (.CI(n28726), .I0(n2858), .I1(GND_net), 
            .CO(n28727));
    SB_LUT4 mux_70_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_106[6]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1859 (.I0(bit_ctr[0]), .I1(n40229), .I2(n4442), 
            .I3(GND_net), .O(n33443));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1859.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1318_13 (.CI(n28925), .I0(n1948), .I1(VCC_net), 
            .CO(n28926));
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n28924), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2958_adj_4802), .I1(VCC_net), 
            .CO(n28726));
    SB_CARRY rem_4_add_1318_12 (.CI(n28924), .I0(n1949), .I1(VCC_net), 
            .CO(n28925));
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n28923), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_11 (.CI(n28923), .I0(n1950), .I1(VCC_net), 
            .CO(n28924));
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n28922), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_24_lut (.I0(duty[22]), .I1(n43164), .I2(n3), .I3(n28060), 
            .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1318_10 (.CI(n28922), .I0(n1951), .I1(VCC_net), 
            .CO(n28923));
    SB_LUT4 add_565_23_lut (.I0(duty[21]), .I1(n43164), .I2(n4), .I3(n28059), 
            .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n28921), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4913), .I3(n28725), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_565_23 (.CI(n28059), .I0(n43164), .I1(n4), .CO(n28060));
    SB_LUT4 add_565_22_lut (.I0(duty[20]), .I1(n43164), .I2(n5), .I3(n28058), 
            .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_22 (.CI(n28058), .I0(n43164), .I1(n5), .CO(n28059));
    SB_LUT4 mux_71_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_565_21_lut (.I0(duty[19]), .I1(n43164), .I2(n6), .I3(n28057), 
            .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_21 (.CI(n28057), .I0(n43164), .I1(n6), .CO(n28058));
    SB_LUT4 add_565_20_lut (.I0(duty[18]), .I1(n43164), .I2(n7), .I3(n28056), 
            .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_20 (.CI(n28056), .I0(n43164), .I1(n7), .CO(n28057));
    SB_LUT4 add_565_19_lut (.I0(duty[17]), .I1(n43164), .I2(n8_adj_4674), 
            .I3(n28055), .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_19 (.CI(n28055), .I0(n43164), .I1(n8_adj_4674), .CO(n28056));
    SB_CARRY rem_4_add_1318_9 (.CI(n28921), .I0(n1952), .I1(VCC_net), 
            .CO(n28922));
    SB_LUT4 div_46_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4914), .I3(n28724), .O(n3_adj_4702)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_18_lut (.I0(duty[16]), .I1(n43164), .I2(n9), .I3(n28054), 
            .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_18 (.CI(n28054), .I0(n43164), .I1(n9), .CO(n28055));
    SB_CARRY div_46_unary_minus_2_add_3_24 (.CI(n28724), .I0(GND_net), .I1(n3_adj_4914), 
            .CO(n28725));
    SB_LUT4 add_565_17_lut (.I0(duty[15]), .I1(n43164), .I2(n10_adj_4675), 
            .I3(n28053), .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_17 (.CI(n28053), .I0(n43164), .I1(n10_adj_4675), 
            .CO(n28054));
    SB_LUT4 div_46_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4915), .I3(n28723), .O(n4_adj_4717)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_16_lut (.I0(duty[14]), .I1(n43164), .I2(n11), .I3(n28052), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_16 (.CI(n28052), .I0(n43164), .I1(n11), .CO(n28053));
    SB_LUT4 add_565_15_lut (.I0(duty[13]), .I1(n43164), .I2(n12), .I3(n28051), 
            .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_46_unary_minus_2_add_3_23 (.CI(n28723), .I0(GND_net), .I1(n4_adj_4915), 
            .CO(n28724));
    SB_CARRY add_565_15 (.CI(n28051), .I0(n43164), .I1(n12), .CO(n28052));
    SB_LUT4 div_46_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4916), .I3(n28722), .O(n5_adj_4716)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_14_lut (.I0(duty[12]), .I1(n43164), .I2(n13), .I3(n28050), 
            .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_14 (.CI(n28050), .I0(n43164), .I1(n13), .CO(n28051));
    SB_LUT4 add_565_13_lut (.I0(duty[11]), .I1(n43164), .I2(n14), .I3(n28049), 
            .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_13 (.CI(n28049), .I0(n43164), .I1(n14), .CO(n28050));
    SB_LUT4 add_565_12_lut (.I0(duty[10]), .I1(n43164), .I2(n15_adj_4676), 
            .I3(n28048), .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n28920), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_565_12 (.CI(n28048), .I0(n43164), .I1(n15_adj_4676), 
            .CO(n28049));
    SB_CARRY rem_4_add_1318_8 (.CI(n28920), .I0(n1953), .I1(VCC_net), 
            .CO(n28921));
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n28919), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_22 (.CI(n28722), .I0(GND_net), .I1(n5_adj_4916), 
            .CO(n28723));
    SB_LUT4 add_565_11_lut (.I0(duty[9]), .I1(n43164), .I2(n16), .I3(n28047), 
            .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_11 (.CI(n28047), .I0(n43164), .I1(n16), .CO(n28048));
    SB_LUT4 add_565_10_lut (.I0(duty[8]), .I1(n43164), .I2(n17), .I3(n28046), 
            .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1318_7 (.CI(n28919), .I0(n1954), .I1(GND_net), 
            .CO(n28920));
    SB_CARRY add_565_10 (.CI(n28046), .I0(n43164), .I1(n17), .CO(n28047));
    SB_LUT4 div_46_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4917), .I3(n28721), .O(n6_adj_4715)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_9_lut (.I0(duty[7]), .I1(n43164), .I2(n18), .I3(n28045), 
            .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_9 (.CI(n28045), .I0(n43164), .I1(n18), .CO(n28046));
    SB_LUT4 add_565_8_lut (.I0(duty[6]), .I1(n43164), .I2(n19), .I3(n28044), 
            .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_8 (.CI(n28044), .I0(n43164), .I1(n19), .CO(n28045));
    SB_LUT4 add_565_7_lut (.I0(duty[5]), .I1(n43164), .I2(n20), .I3(n28043), 
            .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n28918), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_21 (.CI(n28721), .I0(GND_net), .I1(n6_adj_4917), 
            .CO(n28722));
    SB_CARRY add_565_7 (.CI(n28043), .I0(n43164), .I1(n20), .CO(n28044));
    SB_LUT4 div_46_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4918), .I3(n28720), .O(n7_adj_4720)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_565_6_lut (.I0(duty[4]), .I1(n43164), .I2(n21), .I3(n28042), 
            .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_46_unary_minus_2_add_3_20 (.CI(n28720), .I0(GND_net), .I1(n7_adj_4918), 
            .CO(n28721));
    SB_CARRY add_565_6 (.CI(n28042), .I0(n43164), .I1(n21), .CO(n28043));
    SB_LUT4 add_565_5_lut (.I0(duty[3]), .I1(n43164), .I2(n22), .I3(n28041), 
            .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_70_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_106[7]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_6 (.CI(n28918), .I0(n1955), .I1(GND_net), 
            .CO(n28919));
    SB_LUT4 div_46_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4919), .I3(n28719), .O(n8_adj_4719)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_565_5 (.CI(n28041), .I0(n43164), .I1(n22), .CO(n28042));
    SB_LUT4 add_565_4_lut (.I0(duty[2]), .I1(n43164), .I2(n23), .I3(n28040), 
            .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_4 (.CI(n28040), .I0(n43164), .I1(n23), .CO(n28041));
    SB_LUT4 add_565_3_lut (.I0(duty[1]), .I1(n43164), .I2(n24), .I3(n28039), 
            .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_3 (.CI(n28039), .I0(n43164), .I1(n24), .CO(n28040));
    SB_LUT4 add_565_2_lut (.I0(duty[0]), .I1(n43164), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_565_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_565_2 (.CI(VCC_net), .I0(n43164), .I1(n25), .CO(n28039));
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n28917), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_5 (.CI(n28917), .I0(n1956), .I1(VCC_net), 
            .CO(n28918));
    SB_CARRY div_46_unary_minus_2_add_3_19 (.CI(n28719), .I0(GND_net), .I1(n8_adj_4919), 
            .CO(n28720));
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n28916), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4920), .I3(n28718), .O(n9_adj_4718)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_4 (.CI(n28916), .I0(n1957), .I1(VCC_net), 
            .CO(n28917));
    SB_CARRY div_46_unary_minus_2_add_3_18 (.CI(n28718), .I0(GND_net), .I1(n9_adj_4920), 
            .CO(n28719));
    SB_DFF blink_53 (.Q(blink), .C(LED_c), .D(blink_N_255));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(n28915), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4921), .I3(n28717), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_3 (.CI(n28915), .I0(n1958), .I1(GND_net), 
            .CO(n28916));
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n2058), .I1(VCC_net), 
            .CO(n28915));
    SB_LUT4 rem_4_add_1385_19_lut (.I0(n2075_adj_4994), .I1(n2042), .I2(VCC_net), 
            .I3(n28914), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY div_46_unary_minus_2_add_3_17 (.CI(n28717), .I0(GND_net), .I1(n10_adj_4921), 
            .CO(n28718));
    SB_LUT4 div_46_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4922), .I3(n28716), .O(n11_adj_4725)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_18_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n28913), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_18 (.CI(n28913), .I0(n2043), .I1(VCC_net), 
            .CO(n28914));
    SB_LUT4 mux_71_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY div_46_unary_minus_2_add_3_16 (.CI(n28716), .I0(GND_net), .I1(n11_adj_4922), 
            .CO(n28717));
    SB_LUT4 div_46_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4923), .I3(n28715), .O(n12_adj_4724)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n28912), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_15 (.CI(n28715), .I0(GND_net), .I1(n12_adj_4923), 
            .CO(n28716));
    SB_LUT4 div_46_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4924), .I3(n28714), .O(n13_adj_4723)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_14 (.CI(n28714), .I0(GND_net), .I1(n13_adj_4924), 
            .CO(n28715));
    SB_CARRY rem_4_add_1385_17 (.CI(n28912), .I0(n2044), .I1(VCC_net), 
            .CO(n28913));
    SB_LUT4 div_46_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4925), .I3(n28713), .O(n14_adj_4722)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n28911), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24_3_lut_adj_1860 (.I0(n40224), .I1(bit_ctr[9]), .I2(n4442), 
            .I3(GND_net), .O(n33431));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1860.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_106[8]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_16 (.CI(n28911), .I0(n2045), .I1(VCC_net), 
            .CO(n28912));
    SB_LUT4 div_46_i1470_3_lut_3_lut (.I0(n2192), .I1(n6046), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n28910), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12876_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17605));   // verilog/coms.v(126[12] 292[6])
    defparam i12876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12877_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17606));   // verilog/coms.v(126[12] 292[6])
    defparam i12877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12878_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17607));   // verilog/coms.v(126[12] 292[6])
    defparam i12878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12879_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17608));   // verilog/coms.v(126[12] 292[6])
    defparam i12879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12880_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13263), .I3(GND_net), .O(n17609));   // verilog/coms.v(126[12] 292[6])
    defparam i12880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12881_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13263), .I3(GND_net), .O(n17610));   // verilog/coms.v(126[12] 292[6])
    defparam i12881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12882_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13263), .I3(GND_net), .O(n17611));   // verilog/coms.v(126[12] 292[6])
    defparam i12882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12883_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13263), .I3(GND_net), .O(n17612));   // verilog/coms.v(126[12] 292[6])
    defparam i12883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12884_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13263), .I3(GND_net), .O(n17613));   // verilog/coms.v(126[12] 292[6])
    defparam i12884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12885_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13263), .I3(GND_net), .O(n17614));   // verilog/coms.v(126[12] 292[6])
    defparam i12885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12886_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13263), .I3(GND_net), .O(n17615));   // verilog/coms.v(126[12] 292[6])
    defparam i12886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12887_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13263), .I3(GND_net), .O(n17616));   // verilog/coms.v(126[12] 292[6])
    defparam i12887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12888_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13263), .I3(GND_net), .O(n17617));   // verilog/coms.v(126[12] 292[6])
    defparam i12888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12889_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13263), .I3(GND_net), .O(n17618));   // verilog/coms.v(126[12] 292[6])
    defparam i12889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12890_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13263), .I3(GND_net), .O(n17619));   // verilog/coms.v(126[12] 292[6])
    defparam i12890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12891_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13263), .I3(GND_net), .O(n17620));   // verilog/coms.v(126[12] 292[6])
    defparam i12891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12892_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13263), .I3(GND_net), .O(n17621));   // verilog/coms.v(126[12] 292[6])
    defparam i12892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12893_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13263), .I3(GND_net), .O(n17622));   // verilog/coms.v(126[12] 292[6])
    defparam i12893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12894_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13263), .I3(GND_net), .O(n17623));   // verilog/coms.v(126[12] 292[6])
    defparam i12894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12895_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13263), .I3(GND_net), .O(n17624));   // verilog/coms.v(126[12] 292[6])
    defparam i12895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_106[9]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12896_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13263), .I3(GND_net), .O(n17625));   // verilog/coms.v(126[12] 292[6])
    defparam i12896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12897_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13263), .I3(GND_net), .O(n17626));   // verilog/coms.v(126[12] 292[6])
    defparam i12897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12898_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13263), .I3(GND_net), .O(n17627));   // verilog/coms.v(126[12] 292[6])
    defparam i12898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12899_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13263), .I3(GND_net), .O(n17628));   // verilog/coms.v(126[12] 292[6])
    defparam i12899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12900_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13263), .I3(GND_net), .O(n17629));   // verilog/coms.v(126[12] 292[6])
    defparam i12900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12901_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13263), .I3(GND_net), .O(n17630));   // verilog/coms.v(126[12] 292[6])
    defparam i12901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_106[10]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12902_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13263), .I3(GND_net), .O(n17631));   // verilog/coms.v(126[12] 292[6])
    defparam i12902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1861 (.I0(r_SM_Main_adj_5379[1]), .I1(r_SM_Main_adj_5379[0]), 
            .I2(r_SM_Main_adj_5379[2]), .I3(r_SM_Main_2__N_3579[1]), .O(n43694));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_adj_1861.LUT_INIT = 16'h0800;
    SB_LUT4 i12903_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13263), .I3(GND_net), .O(n17632));   // verilog/coms.v(126[12] 292[6])
    defparam i12903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12904_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13263), .I3(GND_net), .O(n17633));   // verilog/coms.v(126[12] 292[6])
    defparam i12904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12905_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13263), .I3(GND_net), .O(n17634));   // verilog/coms.v(126[12] 292[6])
    defparam i12905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_106[11]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1862 (.I0(n40223), .I1(bit_ctr[10]), .I2(n4442), 
            .I3(GND_net), .O(n33429));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1862.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_106[12]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12906_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13263), .I3(GND_net), .O(n17635));   // verilog/coms.v(126[12] 292[6])
    defparam i12906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12907_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13263), .I3(GND_net), .O(n17636));   // verilog/coms.v(126[12] 292[6])
    defparam i12907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12908_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13263), .I3(GND_net), .O(n17637));   // verilog/coms.v(126[12] 292[6])
    defparam i12908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_106[13]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12909_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13263), .I3(GND_net), .O(n17638));   // verilog/coms.v(126[12] 292[6])
    defparam i12909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12910_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13263), .I3(GND_net), .O(n17639));   // verilog/coms.v(126[12] 292[6])
    defparam i12910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12911_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13263), .I3(GND_net), .O(n17640));   // verilog/coms.v(126[12] 292[6])
    defparam i12911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12912_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13263), .I3(GND_net), .O(n17641));   // verilog/coms.v(126[12] 292[6])
    defparam i12912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12913_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13263), .I3(GND_net), .O(n17642));   // verilog/coms.v(126[12] 292[6])
    defparam i12913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_106[14]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12914_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13263), .I3(GND_net), .O(n17643));   // verilog/coms.v(126[12] 292[6])
    defparam i12914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut_adj_1863 (.I0(color_23__N_164[3]), .I1(color_23__N_164[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5260));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i3_2_lut_adj_1863.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(color_23__N_164[4]), .I1(color_23__N_164[6]), 
            .I2(color_23__N_164[2]), .I3(color_23__N_164[0]), .O(n13_adj_5259));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    SB_LUT4 i12915_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13263), .I3(GND_net), .O(n17644));   // verilog/coms.v(126[12] 292[6])
    defparam i12915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1865 (.I0(color_23__N_164[7]), .I1(n13_adj_5259), 
            .I2(n11_adj_5260), .I3(color_23__N_164[1]), .O(n15_adj_4714));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1865.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_71_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_106[15]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1467_3_lut_3_lut (.I0(n2192), .I1(n6043), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_adj_1866 (.I0(color_23__N_164[1]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n37586));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_2_lut_adj_1866.LUT_INIT = 16'heeee;
    SB_LUT4 mux_71_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_106[16]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12916_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13263), .I3(GND_net), .O(n17645));   // verilog/coms.v(126[12] 292[6])
    defparam i12916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12917_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13263), .I3(GND_net), .O(n17646));   // verilog/coms.v(126[12] 292[6])
    defparam i12917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12918_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13263), .I3(GND_net), .O(n17647));   // verilog/coms.v(126[12] 292[6])
    defparam i12918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12919_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13263), .I3(GND_net), .O(n17648));   // verilog/coms.v(126[12] 292[6])
    defparam i12919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12920_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13263), .I3(GND_net), .O(n17649));   // verilog/coms.v(126[12] 292[6])
    defparam i12920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12921_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13263), .I3(GND_net), .O(n17650));   // verilog/coms.v(126[12] 292[6])
    defparam i12921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12922_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13263), .I3(GND_net), .O(n17651));   // verilog/coms.v(126[12] 292[6])
    defparam i12922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12923_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13263), .I3(GND_net), .O(n17652));   // verilog/coms.v(126[12] 292[6])
    defparam i12923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12924_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13263), .I3(GND_net), .O(n17653));   // verilog/coms.v(126[12] 292[6])
    defparam i12924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12925_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13263), .I3(GND_net), .O(n17654));   // verilog/coms.v(126[12] 292[6])
    defparam i12925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12926_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13263), .I3(GND_net), .O(n17655));   // verilog/coms.v(126[12] 292[6])
    defparam i12926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12927_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13263), .I3(GND_net), .O(n17656));   // verilog/coms.v(126[12] 292[6])
    defparam i12927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12928_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13263), .I3(GND_net), .O(n17657));   // verilog/coms.v(126[12] 292[6])
    defparam i12928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_106[17]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(color_23__N_164[7]), .I1(n13_adj_5259), 
            .I2(n11_adj_5260), .I3(n37586), .O(n17111));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i13293_3_lut (.I0(color[1]), .I1(n17111), .I2(n15_adj_4714), 
            .I3(GND_net), .O(n18022));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i13293_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12929_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13263), .I3(GND_net), .O(n17658));   // verilog/coms.v(126[12] 292[6])
    defparam i12929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_106[18]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12930_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13263), .I3(GND_net), .O(n17659));   // verilog/coms.v(126[12] 292[6])
    defparam i12930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12931_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13263), .I3(GND_net), .O(n17660));   // verilog/coms.v(126[12] 292[6])
    defparam i12931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12932_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13263), .I3(GND_net), .O(n17661));   // verilog/coms.v(126[12] 292[6])
    defparam i12932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_106[19]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12933_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13263), .I3(GND_net), .O(n17662));   // verilog/coms.v(126[12] 292[6])
    defparam i12933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12934_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13263), .I3(GND_net), .O(n17663));   // verilog/coms.v(126[12] 292[6])
    defparam i12934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_106[20]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2858), .I1(n2925), .I2(n2867), .I3(GND_net), 
            .O(n2957_adj_4803));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12935_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13263), .I3(GND_net), .O(n17664));   // verilog/coms.v(126[12] 292[6])
    defparam i12935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12936_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13263), .I3(GND_net), .O(n17665));   // verilog/coms.v(126[12] 292[6])
    defparam i12936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12937_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13263), .I3(GND_net), .O(n17666));   // verilog/coms.v(126[12] 292[6])
    defparam i12937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_106[21]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12582_4_lut (.I0(n17189), .I1(r_Bit_Index_adj_5381[2]), .I2(n4670), 
            .I3(n17058), .O(n17311));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12582_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i12938_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13263), .I3(GND_net), .O(n17667));   // verilog/coms.v(126[12] 292[6])
    defparam i12938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12939_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13263), .I3(GND_net), .O(n17668));   // verilog/coms.v(126[12] 292[6])
    defparam i12939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1465_3_lut_3_lut (.I0(n2192), .I1(n6041), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12940_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13263), .I3(GND_net), .O(n17669));   // verilog/coms.v(126[12] 292[6])
    defparam i12940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12941_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13263), .I3(GND_net), .O(n17670));   // verilog/coms.v(126[12] 292[6])
    defparam i12941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_106[22]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12942_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13263), .I3(GND_net), .O(n17671));   // verilog/coms.v(126[12] 292[6])
    defparam i12942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12943_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13263), .I3(GND_net), .O(n17672));   // verilog/coms.v(126[12] 292[6])
    defparam i12943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1868 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5265));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i4_4_lut_adj_1868.LUT_INIT = 16'hfffe;
    SB_LUT4 i12944_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13263), .I3(GND_net), .O(n17673));   // verilog/coms.v(126[12] 292[6])
    defparam i12944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1869 (.I0(control_mode[6]), .I1(n10_adj_5265), 
            .I2(control_mode[2]), .I3(GND_net), .O(n15778));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i5_3_lut_adj_1869.LUT_INIT = 16'hfefe;
    SB_LUT4 i12945_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13263), .I3(GND_net), .O(n17674));   // verilog/coms.v(126[12] 292[6])
    defparam i12945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12946_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13263), .I3(GND_net), .O(n17675));   // verilog/coms.v(126[12] 292[6])
    defparam i12946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n15778), 
            .I3(GND_net), .O(n15_adj_4673));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i12947_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13263), .I3(GND_net), .O(n17676));   // verilog/coms.v(126[12] 292[6])
    defparam i12947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4673), .I3(n15), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12948_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13263), .I3(GND_net), .O(n17677));   // verilog/coms.v(126[12] 292[6])
    defparam i12948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_106[23]), 
            .I2(n15_adj_4672), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12949_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13263), .I3(GND_net), .O(n17678));   // verilog/coms.v(126[12] 292[6])
    defparam i12949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12950_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13263), .I3(GND_net), .O(n17679));   // verilog/coms.v(126[12] 292[6])
    defparam i12950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12951_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13263), .I3(GND_net), .O(n17680));   // verilog/coms.v(126[12] 292[6])
    defparam i12951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1475_3_lut_3_lut (.I0(n2192), .I1(n6051), .I2(n663), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12952_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13263), .I3(GND_net), .O(n17681));   // verilog/coms.v(126[12] 292[6])
    defparam i12952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12953_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13263), .I3(GND_net), .O(n17682));   // verilog/coms.v(126[12] 292[6])
    defparam i12953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12954_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13263), .I3(GND_net), .O(n17683));   // verilog/coms.v(126[12] 292[6])
    defparam i12954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12955_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13263), .I3(GND_net), .O(n17684));   // verilog/coms.v(126[12] 292[6])
    defparam i12955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12956_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13263), .I3(GND_net), .O(n17685));   // verilog/coms.v(126[12] 292[6])
    defparam i12956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12957_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13263), .I3(GND_net), .O(n17686));   // verilog/coms.v(126[12] 292[6])
    defparam i12957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12958_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13263), .I3(GND_net), .O(n17687));   // verilog/coms.v(126[12] 292[6])
    defparam i12958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12959_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13263), .I3(GND_net), .O(n17688));   // verilog/coms.v(126[12] 292[6])
    defparam i12959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12960_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13263), 
            .I3(GND_net), .O(n17689));   // verilog/coms.v(126[12] 292[6])
    defparam i12960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12961_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13263), 
            .I3(GND_net), .O(n17690));   // verilog/coms.v(126[12] 292[6])
    defparam i12961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12962_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13263), 
            .I3(GND_net), .O(n17691));   // verilog/coms.v(126[12] 292[6])
    defparam i12962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12963_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13263), 
            .I3(GND_net), .O(n17692));   // verilog/coms.v(126[12] 292[6])
    defparam i12963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12964_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13263), 
            .I3(GND_net), .O(n17693));   // verilog/coms.v(126[12] 292[6])
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12965_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13263), 
            .I3(GND_net), .O(n17694));   // verilog/coms.v(126[12] 292[6])
    defparam i12965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12966_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13263), 
            .I3(GND_net), .O(n17695));   // verilog/coms.v(126[12] 292[6])
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4750));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12967_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13263), 
            .I3(GND_net), .O(n17696));   // verilog/coms.v(126[12] 292[6])
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4749));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4748));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4747));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12968_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13263), 
            .I3(GND_net), .O(n17697));   // verilog/coms.v(126[12] 292[6])
    defparam i12968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12969_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13263), 
            .I3(GND_net), .O(n17698));   // verilog/coms.v(126[12] 292[6])
    defparam i12969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12970_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13263), 
            .I3(GND_net), .O(n17699));   // verilog/coms.v(126[12] 292[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4746));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4745));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12585_4_lut (.I0(n17189), .I1(r_Bit_Index_adj_5381[1]), .I2(r_Bit_Index_adj_5381[0]), 
            .I3(n17058), .O(n17314));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12585_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4744));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4743));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4742));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4741));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857), .I1(n2924), .I2(n2867), .I3(GND_net), 
            .O(n2956_adj_4804));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4740));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4739));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12971_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13263), 
            .I3(GND_net), .O(n17700));   // verilog/coms.v(126[12] 292[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4738));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4737));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4692));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1463_3_lut_3_lut (.I0(n2192), .I1(n6039), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2453_adj_4943));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1462_3_lut_3_lut (.I0(n2192), .I1(n6038), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1601_3_lut (.I0(n2352), .I1(n2419), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2451_adj_4945));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4694));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35010_3_lut (.I0(n2249), .I1(n2316), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34838_3_lut (.I0(n2348), .I1(n2415), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2447_adj_4949));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35012_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34836_3_lut (.I0(n2351), .I1(n2418), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2450_adj_4946));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4695));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4696));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1602_3_lut (.I0(n2353), .I1(n2420), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2452_adj_4944));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35103_3_lut (.I0(n38143), .I1(n2053), .I2(n41429), .I3(GND_net), 
            .O(n2350));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35104_3_lut (.I0(n2350), .I1(n2417), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2449_adj_4947));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1598_3_lut (.I0(n2349), .I1(n2416), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2448_adj_4948));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4697));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357_adj_4954), .I1(n2424), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2456_adj_4940));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1607_3_lut (.I0(n2358_adj_4953), .I1(n2425), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2457_adj_4939));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2455_adj_4941));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2454_adj_4942));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372_adj_4952), 
            .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1870 (.I0(n2439), .I1(n2438), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5317));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1870.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1871 (.I0(n2456_adj_4940), .I1(n2458_adj_4938), 
            .I2(GND_net), .I3(GND_net), .O(n37972));
    defparam i1_2_lut_adj_1871.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1872 (.I0(n2454_adj_4942), .I1(n37972), .I2(n2455_adj_4941), 
            .I3(n2457_adj_4939), .O(n35658));
    defparam i1_4_lut_adj_1872.LUT_INIT = 16'ha080;
    SB_LUT4 i13_4_lut_adj_1873 (.I0(n2448_adj_4948), .I1(n2449_adj_4947), 
            .I2(n2452_adj_4944), .I3(n18_adj_5317), .O(n30_adj_5313));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1874 (.I0(n2444), .I1(n2445), .I2(n35658), .I3(n2453_adj_4943), 
            .O(n28_adj_5315));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1874.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1875 (.I0(n2446), .I1(n2450_adj_4946), .I2(n2447_adj_4949), 
            .I3(n2451_adj_4945), .O(n29_adj_5314));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1876 (.I0(n2440), .I1(n2442), .I2(n2441), .I3(n2443), 
            .O(n27_adj_5316));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1876.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1877 (.I0(n27_adj_5316), .I1(n29_adj_5314), .I2(n28_adj_5315), 
            .I3(n30_adj_5313), .O(n2471_adj_4937));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1877.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4772), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458_adj_4938));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4698));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12972_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13263), 
            .I3(GND_net), .O(n17701));   // verilog/coms.v(126[12] 292[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36317_1_lut (.I0(n3263), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43147));
    defparam i36317_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12973_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13263), 
            .I3(GND_net), .O(n17702));   // verilog/coms.v(126[12] 292[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12974_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13263), 
            .I3(GND_net), .O(n17703));   // verilog/coms.v(126[12] 292[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1878 (.I0(n40273), .I1(byte_transmit_counter[5]), 
            .I2(n24391), .I3(GND_net), .O(n34001));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut_adj_1878.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1879 (.I0(n40274), .I1(byte_transmit_counter[4]), 
            .I2(n24391), .I3(GND_net), .O(n34037));   // verilog/coms.v(126[12] 292[6])
    defparam i12_3_lut_adj_1879.LUT_INIT = 16'hcaca;
    SB_LUT4 i22930_2_lut_3_lut (.I0(n749), .I1(n855), .I2(n748), .I3(GND_net), 
            .O(n6_adj_5304));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i22930_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4705));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1880 (.I0(n2956_adj_4804), .I1(n2957_adj_4803), 
            .I2(n2958_adj_4802), .I3(GND_net), .O(n35625));
    defparam i1_3_lut_adj_1880.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1881 (.I0(n2954_adj_4806), .I1(n2941), .I2(n35625), 
            .I3(n2955_adj_4805), .O(n27_adj_5331));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1881.LUT_INIT = 16'heccc;
    SB_LUT4 i13_4_lut_adj_1882 (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35_adj_5326));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1882.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n749), .I1(n855), .I2(n884), .I3(n748), 
            .O(n955));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hef10;
    SB_LUT4 i13333_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1172), .I3(GND_net), .O(n18062));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1461_3_lut_3_lut (.I0(n2192), .I1(n6037), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12975_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13263), 
            .I3(GND_net), .O(n17704));   // verilog/coms.v(126[12] 292[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12976_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13263), 
            .I3(GND_net), .O(n17705));   // verilog/coms.v(126[12] 292[6])
    defparam i12976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12977_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13263), 
            .I3(GND_net), .O(n17706));   // verilog/coms.v(126[12] 292[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164), .I3(GND_net), 
            .O(n3240));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164), .I3(GND_net), 
            .O(n3231));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215), .I2(n3164), .I3(GND_net), 
            .O(n3247));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209), .I2(n3164), .I3(GND_net), 
            .O(n3241));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214), .I2(n3164), .I3(GND_net), 
            .O(n3246));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1883 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_5327));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1883.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164), .I3(GND_net), 
            .O(n3235));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2138_3_lut (.I0(n3145), .I1(n3212), .I2(n3164), .I3(GND_net), 
            .O(n3244));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164), .I3(GND_net), 
            .O(n3236));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164), .I3(GND_net), 
            .O(n3233));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164), .I3(GND_net), 
            .O(n3234));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1884 (.I0(n35_adj_5326), .I1(n27_adj_5331), .I2(n2949_adj_4811), 
            .I3(n2942), .O(n40_adj_5318));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1884.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2142_3_lut (.I0(n3149), .I1(n3216), .I2(n3164), .I3(GND_net), 
            .O(n3248));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164), .I3(GND_net), 
            .O(n3239));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1885 (.I0(n2741), .I1(n2754), .I2(n35608), .I3(n2755), 
            .O(n24_adj_4817));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1885.LUT_INIT = 16'heaaa;
    SB_LUT4 i16_4_lut_adj_1886 (.I0(n2951_adj_4809), .I1(n2952_adj_4808), 
            .I2(n2947_adj_4813), .I3(n2946_adj_4814), .O(n38_adj_5320));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1886.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220), .I2(n3164), .I3(GND_net), 
            .O(n3252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164), .I3(GND_net), 
            .O(n3232));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211), .I2(n3164), .I3(GND_net), 
            .O(n3243));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2143_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221), .I2(n3164), .I3(GND_net), 
            .O(n3253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164), .I3(GND_net), 
            .O(n3238));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164), .I3(GND_net), 
            .O(n3237));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213), .I2(n3164), .I3(GND_net), 
            .O(n3245));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2144_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223), .I2(n3164), .I3(GND_net), 
            .O(n3255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210), .I2(n3164), .I3(GND_net), 
            .O(n3242));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222), .I2(n3164), .I3(GND_net), 
            .O(n3254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225), .I2(n3164), .I3(GND_net), 
            .O(n3257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224), .I2(n3164), .I3(GND_net), 
            .O(n3256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1887 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n35692));
    defparam i1_3_lut_adj_1887.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut_adj_1888 (.I0(n3254), .I1(n3242), .I2(n35692), .I3(n3255), 
            .O(n34_adj_5330));
    defparam i9_4_lut_adj_1888.LUT_INIT = 16'heccc;
    SB_LUT4 i16_4_lut_adj_1889 (.I0(n3250), .I1(n3245), .I2(n3237), .I3(n3238), 
            .O(n41_adj_5324));
    defparam i16_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n3253), .I1(n3249), .I2(n3243), .I3(GND_net), 
            .O(n38_adj_5329));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1890 (.I0(n3232), .I1(n3252), .I2(n3239), .I3(n3248), 
            .O(n43_adj_5323));
    defparam i18_4_lut_adj_1890.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1891 (.I0(n3234), .I1(n3230), .I2(n3233), .I3(n3236), 
            .O(n40_adj_5325));
    defparam i15_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n41_adj_5324), .I1(n3244), .I2(n34_adj_5330), 
            .I3(n3235), .O(n46_adj_5321));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1892 (.I0(n3246), .I1(n3241), .I2(n3251), .I3(n3247), 
            .O(n39_adj_5328));
    defparam i14_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1893 (.I0(n43_adj_5323), .I1(n3231), .I2(n38_adj_5329), 
            .I3(n3240), .O(n47));
    defparam i22_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_5328), .I2(n46_adj_5321), 
            .I3(n40_adj_5325), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1464_3_lut_3_lut (.I0(n2192), .I1(n6040), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12978_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13263), 
            .I3(GND_net), .O(n17707));   // verilog/coms.v(126[12] 292[6])
    defparam i12978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12979_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13263), 
            .I3(GND_net), .O(n17708));   // verilog/coms.v(126[12] 292[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12980_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13263), 
            .I3(GND_net), .O(n17709));   // verilog/coms.v(126[12] 292[6])
    defparam i12980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1460_3_lut_3_lut (.I0(n2192), .I1(n6036), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34841_3_lut (.I0(n2153), .I1(n2220), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34845_3_lut (.I0(n2149), .I1(n2216), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34846_3_lut (.I0(n2248), .I1(n2315), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34843_3_lut (.I0(n2150), .I1(n2217), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2346));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1474_3_lut_3_lut (.I0(n2192), .I1(n6050), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34597_3_lut (.I0(n2273_adj_4962), .I1(n2174_adj_4975), .I2(n2075_adj_4994), 
            .I3(GND_net), .O(n41429));
    defparam i34597_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1398_rep_25_3_lut (.I0(n2120), .I1(n2219), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n38149));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1398_rep_25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1465_rep_19_3_lut (.I0(n38149), .I1(n2318), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n38143));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1465_rep_19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1535_3_lut (.I0(n2254), .I1(n2321), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1531_3_lut (.I0(n2250), .I1(n2317), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1534_3_lut (.I0(n2253), .I1(n2320), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2357_adj_4954));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273_adj_4962), 
            .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1894 (.I0(n2356), .I1(n2358_adj_4953), .I2(GND_net), 
            .I3(GND_net), .O(n37728));
    defparam i1_2_lut_adj_1894.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n2354), .I1(n37728), .I2(n2355), .I3(n2357_adj_4954), 
            .O(n35590));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'ha080;
    SB_LUT4 i12_4_lut_adj_1896 (.I0(n2352), .I1(n2349), .I2(n2353), .I3(n2350), 
            .O(n28_adj_4843));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1896.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1897 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n35590), 
            .O(n26_adj_4859));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1897.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1898 (.I0(n2346), .I1(n2348), .I2(n2347), .I3(n2351), 
            .O(n27_adj_4851));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1899 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_4888));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1899.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1900 (.I0(n25_adj_4888), .I1(n27_adj_4851), .I2(n26_adj_4859), 
            .I3(n28_adj_4843), .O(n2372_adj_4952));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4773), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358_adj_4953));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12981_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13263), 
            .I3(GND_net), .O(n17710));   // verilog/coms.v(126[12] 292[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13318_3_lut (.I0(setpoint[10]), .I1(n4359), .I2(n36881), 
            .I3(GND_net), .O(n18047));   // verilog/coms.v(126[12] 292[6])
    defparam i13318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12982_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13263), 
            .I3(GND_net), .O(n17711));   // verilog/coms.v(126[12] 292[6])
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4912));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4911));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4910));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4909));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1467_3_lut (.I0(n2154), .I1(n2221), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1472_3_lut_3_lut (.I0(n2192), .I1(n6048), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35115_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1464_3_lut (.I0(n2151), .I1(n2218), .I2(n2174_adj_4975), 
            .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1901 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n35653));
    defparam i1_3_lut_adj_1901.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1902 (.I0(n2250), .I1(n2252), .I2(n2251), .I3(n2253), 
            .O(n26_adj_5333));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1903 (.I0(n2254), .I1(n2246), .I2(n35653), .I3(n2255), 
            .O(n19_adj_5335));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1903.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_1904 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5336));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1904.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1905 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_5334));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1906 (.I0(n19_adj_5335), .I1(n26_adj_5333), .I2(n2249), 
            .I3(n2247), .O(n28_adj_5332));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1906.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1907 (.I0(n2248), .I1(n28_adj_5332), .I2(n24_adj_5334), 
            .I3(n16_adj_5336), .O(n2273_adj_4962));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4774), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12983_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13263), 
            .I3(GND_net), .O(n17712));   // verilog/coms.v(126[12] 292[6])
    defparam i12983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1473_3_lut_3_lut (.I0(n2192), .I1(n6049), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1469_3_lut_3_lut (.I0(n2192), .I1(n6045), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4908));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12984_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13263), .I3(GND_net), .O(n17713));   // verilog/coms.v(126[12] 292[6])
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12985_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13263), .I3(GND_net), .O(n17714));   // verilog/coms.v(126[12] 292[6])
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4907));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4906));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12987_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13263), .I3(GND_net), .O(n17716));   // verilog/coms.v(126[12] 292[6])
    defparam i12987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_3_lut (.I0(n2945_adj_4815), .I1(n34_adj_5327), .I2(n2944), 
            .I3(GND_net), .O(n39_adj_5319));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_i1468_3_lut_3_lut (.I0(n2192), .I1(n6044), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i15_4_lut_adj_1908 (.I0(n2948_adj_4812), .I1(n2943), .I2(n2953_adj_4807), 
            .I3(n2950_adj_4810), .O(n37_adj_5322));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1908.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1909 (.I0(n37_adj_5322), .I1(n39_adj_5319), .I2(n38_adj_5320), 
            .I3(n40_adj_5318), .O(n2966_adj_4798));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i21_4_lut_adj_1909.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908), .I2(n2867), .I3(GND_net), 
            .O(n2940));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1997_3_lut (.I0(n2940), .I1(n3007_adj_4790), .I2(n2966_adj_4798), 
            .I3(GND_net), .O(n3039));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1466_3_lut_3_lut (.I0(n2192), .I1(n6042), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5303));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5302));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5301));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5300));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36326_1_lut (.I0(n2669), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43156));
    defparam i36326_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5299));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1594_3_lut_3_lut (.I0(n2381), .I1(n6085), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1599_3_lut_3_lut (.I0(n2381), .I1(n6090), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5298));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5297));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5296));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5295));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5294));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5293));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5292));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5291));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5290));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5289));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5288));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5287));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5286));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5285));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5284));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5283));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5282));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5281));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5280));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5279));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .GND_net(GND_net), .n34179(n34179), .byte_transmit_counter({Open_0, 
         Open_1, byte_transmit_counter[5:2], Open_2, Open_3}), .n34135(n34135), 
         .n18046(n18046), .setpoint({setpoint}), .n18047(n18047), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n34037(n34037), .n34001(n34001), .n34177(n34177), .\byte_transmit_counter[1] (byte_transmit_counter[1]), 
         .n18057(n18057), .n18058(n18058), .n18059(n18059), .n18060(n18060), 
         .n18048(n18048), .n18049(n18049), .n18050(n18050), .n18051(n18051), 
         .n18052(n18052), .n18053(n18053), .n18054(n18054), .n18055(n18055), 
         .n18056(n18056), .n43329(n43329), .n18042(n18042), .n18043(n18043), 
         .n18044(n18044), .n18045(n18045), .n18040(n18040), .n18041(n18041), 
         .n18038(n18038), .n18039(n18039), .n17960(n17960), .PWMLimit({PWMLimit}), 
         .n17961(n17961), .n17936(n17936), .\data_in_frame[24] ({\data_in_frame[24] }), 
         .n17937(n17937), .n17938(n17938), .n17939(n17939), .n17940(n17940), 
         .n17941(n17941), .n17942(n17942), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .n17962(n17962), .n17963(n17963), .n17964(n17964), .n17965(n17965), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .n17956(n17956), .n17957(n17957), 
         .n17958(n17958), .n17959(n17959), .n17954(n17954), .n17955(n17955), 
         .n17952(n17952), .n17953(n17953), .n17950(n17950), .n17951(n17951), 
         .n17948(n17948), .n17949(n17949), .n17946(n17946), .n17947(n17947), 
         .n17943(n17943), .n17944(n17944), .n17945(n17945), .n17935(n17935), 
         .\data_in_frame[22] ({\data_in_frame[22] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_in_frame[2] ({\data_in_frame[2] [7:3], Open_4, Open_5, 
         Open_6}), .\FRAME_MATCHER.state[1] (\FRAME_MATCHER.state [1]), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .rx_data({rx_data}), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[2][0] (\data_in_frame[2] [0]), .\data_in_frame[2][2] (\data_in_frame[2] [2]), 
         .n17743(n17743), .control_mode({control_mode}), .n17742(n17742), 
         .n17741(n17741), .n17740(n17740), .n17739(n17739), .n17738(n17738), 
         .n17737(n17737), .n17736(n17736), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n17735(n17735), .\data_in_frame[10] ({\data_in_frame[10] }), .n17734(n17734), 
         .rx_data_ready(rx_data_ready), .n17733(n17733), .n17732(n17732), 
         .tx_active(tx_active), .n63(n63), .n17731(n17731), .n17730(n17730), 
         .n17729(n17729), .n17728(n17728), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n17727(n17727), .n17726(n17726), .n17725(n17725), .n17724(n17724), 
         .n17723(n17723), .n17722(n17722), .n17721(n17721), .n17720(n17720), 
         .\data_out_frame[18] ({\data_out_frame[18] [7:3], Open_7, Open_8, 
         Open_9}), .n17719(n17719), .n17718(n17718), .n17717(n17717), 
         .n17716(n17716), .n17714(n17714), .\data_out_frame[18][1] (\data_out_frame[18] [1]), 
         .n17713(n17713), .\data_out_frame[18][0] (\data_out_frame[18] [0]), 
         .n17712(n17712), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n17711(n17711), .n17710(n17710), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .n17709(n17709), .n17708(n17708), .n17707(n17707), .n17706(n17706), 
         .n17705(n17705), .n17704(n17704), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n17703(n17703), .n17702(n17702), .n17701(n17701), .n17700(n17700), 
         .n17699(n17699), .n17698(n17698), .n17697(n17697), .n17696(n17696), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .n17695(n17695), 
         .n17694(n17694), .n17693(n17693), .n17692(n17692), .n17691(n17691), 
         .n17690(n17690), .n17689(n17689), .n17688(n17688), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n17687(n17687), .n17686(n17686), .n17685(n17685), .n17684(n17684), 
         .n17683(n17683), .n17682(n17682), .n17681(n17681), .n17680(n17680), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n17679(n17679), 
         .n17678(n17678), .n17677(n17677), .n17676(n17676), .n17675(n17675), 
         .n17674(n17674), .n17673(n17673), .n17672(n17672), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n17671(n17671), .n17670(n17670), .n17669(n17669), .n17668(n17668), 
         .n17667(n17667), .n17666(n17666), .n17665(n17665), .n17664(n17664), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n17663(n17663), 
         .n17662(n17662), .n17661(n17661), .n17660(n17660), .n17659(n17659), 
         .n17658(n17658), .n17657(n17657), .n17656(n17656), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n17655(n17655), .n17654(n17654), .n17653(n17653), .n17652(n17652), 
         .n17651(n17651), .n17650(n17650), .n17649(n17649), .n17648(n17648), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .n17647(n17647), .n17646(n17646), 
         .n17645(n17645), .n17644(n17644), .n17643(n17643), .n17642(n17642), 
         .n17641(n17641), .n17640(n17640), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .n17639(n17639), .n17638(n17638), .n17637(n17637), .n17636(n17636), 
         .n17635(n17635), .n17634(n17634), .n17633(n17633), .n17632(n17632), 
         .n17631(n17631), .n17630(n17630), .n17629(n17629), .n17628(n17628), 
         .n17627(n17627), .n17626(n17626), .n17625(n17625), .n17624(n17624), 
         .n17623(n17623), .n17622(n17622), .n17621(n17621), .n17620(n17620), 
         .n17619(n17619), .n17618(n17618), .n17617(n17617), .n17616(n17616), 
         .n17615(n17615), .n17614(n17614), .n17613(n17613), .n17612(n17612), 
         .n17611(n17611), .n17610(n17610), .n17609(n17609), .n17608(n17608), 
         .\data_in[3] ({\data_in[3] }), .n17607(n17607), .n17606(n17606), 
         .n17605(n17605), .n17604(n17604), .n17603(n17603), .n17602(n17602), 
         .n17601(n17601), .n17600(n17600), .\data_in[2] ({\data_in[2] }), 
         .n17599(n17599), .n17598(n17598), .n17597(n17597), .n17596(n17596), 
         .n17595(n17595), .n17594(n17594), .n17593(n17593), .n17592(n17592), 
         .\data_in[1] ({\data_in[1] }), .n17591(n17591), .n17590(n17590), 
         .n17589(n17589), .n17588(n17588), .n17587(n17587), .n17586(n17586), 
         .n17585(n17585), .n17584(n17584), .\data_in[0] ({\data_in[0] }), 
         .n17583(n17583), .n17582(n17582), .n17581(n17581), .n17580(n17580), 
         .n17579(n17579), .n17578(n17578), .n17577(n17577), .\Ki[15] (Ki[15]), 
         .n17576(n17576), .\Ki[14] (Ki[14]), .n17575(n17575), .\Ki[13] (Ki[13]), 
         .n17574(n17574), .\Ki[12] (Ki[12]), .n17573(n17573), .\Ki[11] (Ki[11]), 
         .n17572(n17572), .\Ki[10] (Ki[10]), .n30070(n30070), .n17571(n17571), 
         .\Ki[9] (Ki[9]), .n17570(n17570), .\Ki[8] (Ki[8]), .n17569(n17569), 
         .\Ki[7] (Ki[7]), .n17568(n17568), .\Ki[6] (Ki[6]), .n17567(n17567), 
         .\Ki[5] (Ki[5]), .n17566(n17566), .\Ki[4] (Ki[4]), .n17565(n17565), 
         .\Ki[3] (Ki[3]), .n17564(n17564), .\Ki[2] (Ki[2]), .n17563(n17563), 
         .\Ki[1] (Ki[1]), .n17562(n17562), .\Kp[15] (Kp[15]), .n17561(n17561), 
         .\Kp[14] (Kp[14]), .n17560(n17560), .\Kp[13] (Kp[13]), .n17559(n17559), 
         .\Kp[12] (Kp[12]), .n17558(n17558), .\Kp[11] (Kp[11]), .n17557(n17557), 
         .\Kp[10] (Kp[10]), .\Kp[9] (Kp[9]), .n17555(n17555), .\Kp[8] (Kp[8]), 
         .n17554(n17554), .\Kp[7] (Kp[7]), .n17553(n17553), .\Kp[6] (Kp[6]), 
         .n17552(n17552), .\Kp[5] (Kp[5]), .n17551(n17551), .\Kp[4] (Kp[4]), 
         .n17550(n17550), .\Kp[3] (Kp[3]), .n17549(n17549), .\Kp[2] (Kp[2]), 
         .n17548(n17548), .\Kp[1] (Kp[1]), .n17547(n17547), .gearBoxRatio({gearBoxRatio}), 
         .n4351(n4351), .n17546(n17546), .n17545(n17545), .n17544(n17544), 
         .n17543(n17543), .n17542(n17542), .n4350(n4350), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n17541(n17541), .n17540(n17540), .n17539(n17539), .n17538(n17538), 
         .n17537(n17537), .n17536(n17536), .n17535(n17535), .n4353(n4353), 
         .n17534(n17534), .n17533(n17533), .n4352(n4352), .n17532(n17532), 
         .n17531(n17531), .n17530(n17530), .n17529(n17529), .n17528(n17528), 
         .n17527(n17527), .n4357(n4357), .n17526(n17526), .n17525(n17525), 
         .n17523(n17523), .IntegralLimit({IntegralLimit}), .n17522(n17522), 
         .n4356(n4356), .n4355(n4355), .n4354(n4354), .n17521(n17521), 
         .n17520(n17520), .n17519(n17519), .n788(n788), .n17518(n17518), 
         .n17517(n17517), .n17516(n17516), .n17515(n17515), .n17514(n17514), 
         .n17513(n17513), .n17512(n17512), .n17511(n17511), .n17510(n17510), 
         .n17509(n17509), .n17508(n17508), .n122(n122), .n9001(n9001), 
         .n34675(n34675), .\FRAME_MATCHER.i_31__N_2621 (\FRAME_MATCHER.i_31__N_2621 ), 
         .n17507(n17507), .n17506(n17506), .n3894(n3894), .n17505(n17505), 
         .n5(n5_adj_5312), .n17504(n17504), .n17503(n17503), .n17502(n17502), 
         .n17501(n17501), .n34173(n34173), .n4368(n4368), .n4367(n4367), 
         .n4366(n4366), .n4365(n4365), .n4364(n4364), .n4363(n4363), 
         .n4362(n4362), .n4361(n4361), .n4360(n4360), .n17417(n17417), 
         .n4372(n4372), .n4371(n4371), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n4370(n4370), .LED_c(LED_c), .n4369(n4369), .n34067(n34067), 
         .n17398(n17398), .n17396(n17396), .n17395(n17395), .n17394(n17394), 
         .\Ki[0] (Ki[0]), .n17393(n17393), .\Kp[0] (Kp[0]), .n17392(n17392), 
         .\FRAME_MATCHER.i_31__N_2625 (\FRAME_MATCHER.i_31__N_2625 ), .n17249(n17249), 
         .n40273(n40273), .n40274(n40274), .n40275(n40275), .n40278(n40278), 
         .n40277(n40277), .n40276(n40276), .n36887(n36887), .n24391(n24391), 
         .n4359(n4359), .\displacement[18] (displacement[18]), .n13263(n13263), 
         .\FRAME_MATCHER.state_31__N_2661[2] (\FRAME_MATCHER.state_31__N_2661 [2]), 
         .n7(n7_adj_4818), .\FRAME_MATCHER.state_31__N_2661[0] (\FRAME_MATCHER.state_31__N_2661 [0]), 
         .n4349(n4349), .n2957(n2957_adj_4678), .n36881(n36881), .n4358(n4358), 
         .n17314(n17314), .r_Bit_Index({r_Bit_Index_adj_5381}), .n17311(n17311), 
         .r_SM_Main({r_SM_Main_adj_5379}), .n17446(n17446), .n17412(n17412), 
         .n17411(n17411), .n17410(n17410), .tx_o(tx_o), .VCC_net(VCC_net), 
         .\r_SM_Main_2__N_3579[1] (r_SM_Main_2__N_3579[1]), .n17058(n17058), 
         .n43694(n43694), .n4670(n4670), .n17189(n17189), .n4(n4_adj_4677), 
         .n3(n3_adj_5264), .n8936(n8936), .n10627(n10627), .tx_enable(tx_enable), 
         .n17338(n17338), .r_Bit_Index_adj_11({r_Bit_Index}), .n17341(n17341), 
         .n24450(n24450), .\r_SM_Main[1]_adj_6 (r_SM_Main[1]), .r_Rx_Data(r_Rx_Data), 
         .PIN_13_N_105(PIN_13_N_105), .\r_SM_Main[2]_adj_7 (r_SM_Main[2]), 
         .n40218(n40218), .n40217(n40217), .n17452(n17452), .n17462(n17462), 
         .n4_adj_8(n4_adj_4713), .n17429(n17429), .n17428(n17428), .n17427(n17427), 
         .n17426(n17426), .n17425(n17425), .n17403(n17403), .n17052(n17052), 
         .n17180(n17180), .n4648(n4648), .n17343(n17343), .n17342(n17342), 
         .n43211(n43211), .n15734(n15734), .n15626(n15626), .n23653(n23653), 
         .n4_adj_9(n4_adj_4736), .n4_adj_10(n4_adj_4704)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(202[8] 223[4])
    SB_LUT4 i12613_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n23653), 
            .I3(n15734), .O(n17342));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12613_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12614_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n15626), 
            .I3(n23653), .O(n17343));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12614_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 i12519_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n36115), .I3(GND_net), .O(n17248));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12520_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17249));   // verilog/coms.v(126[12] 292[6])
    defparam i12520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34037_2_lut (.I0(n35424), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n40258));   // verilog/neopixel.v(35[12] 117[6])
    defparam i34037_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31_4_lut (.I0(n40258), .I1(n40256), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n33499));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5278));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5277));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5276));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5275));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5274));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5273));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23068_2_lut (.I0(n855), .I1(n884), .I2(GND_net), .I3(GND_net), 
            .O(n957));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i23068_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25_4_lut (.I0(n15744), .I1(n35327), .I2(state[0]), .I3(n24628), 
            .O(n11_adj_5256));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i12663_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[22] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17392));   // verilog/coms.v(126[12] 292[6])
    defparam i12663_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12664_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n30070), 
            .I3(GND_net), .O(n17393));   // verilog/coms.v(126[12] 292[6])
    defparam i12664_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12665_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n30070), 
            .I3(GND_net), .O(n17394));   // verilog/coms.v(126[12] 292[6])
    defparam i12665_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34094_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34094_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_46_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2), .I3(n5_adj_5257), 
            .O(n35278));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i12666_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17395));   // verilog/coms.v(126[12] 292[6])
    defparam i12666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12667_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17396));   // verilog/coms.v(126[12] 292[6])
    defparam i12667_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34065_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n511), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34065_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_46_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_5307), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_5309), 
            .I3(n35278), .O(n35295));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i34064_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n650), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34064_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_46_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_5305), 
            .I3(n35295), .O(n35299));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2_adj_5308), 
            .I3(n649), .O(n784));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_5306), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_5263), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4689), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i34061_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n651), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34061_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_46_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_4687), 
            .I3(n35299), .O(n914));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553_adj_4871), .I1(n2620_adj_4865), 
            .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542_adj_4882), .I1(n2609), .I2(n2570), 
            .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551_adj_4873), .I1(n2618_adj_4867), 
            .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4688), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552_adj_4872), .I1(n2619_adj_4866), 
            .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539_adj_4885), .I1(n2606), .I2(n2570), 
            .I3(GND_net), .O(n2638_adj_4855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538_adj_4886), .I1(n2605), .I2(n2570), 
            .I3(GND_net), .O(n2637_adj_4856));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544_adj_4880), .I1(n2611), .I2(n2570), 
            .I3(GND_net), .O(n2643_adj_4853));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550_adj_4874), .I1(n2617), .I2(n2570), 
            .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543_adj_4881), .I1(n2610), .I2(n2570), 
            .I3(GND_net), .O(n2642_adj_4854));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545_adj_4879), .I1(n2612), .I2(n2570), 
            .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547_adj_4877), .I1(n2614), .I2(n2570), 
            .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540_adj_4884), .I1(n2607), .I2(n2570), 
            .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546_adj_4878), .I1(n2613), .I2(n2570), 
            .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558_adj_4870), .I1(n2625_adj_4860), 
            .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4862), .I2(n2570), 
            .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4863), .I2(n2570), 
            .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548_adj_4876), .I1(n2615), .I2(n2570), 
            .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541_adj_4883), .I1(n2608), .I2(n2570), 
            .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1739_3_lut (.I0(n2554), .I1(n2621_adj_4864), .I2(n2570), 
            .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1734_3_lut (.I0(n2549_adj_4875), .I1(n2616), .I2(n2570), 
            .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4861), .I2(n2570), 
            .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1910 (.I0(n2648), .I1(n2653), .I2(n2640), .I3(n2647), 
            .O(n30_adj_4823));
    defparam i11_4_lut_adj_1910.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1911 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n37976));
    defparam i1_2_lut_adj_1911.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(n2654), .I1(n37976), .I2(n2655), .I3(n2657), 
            .O(n35671));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'ha080;
    SB_LUT4 i15_4_lut_adj_1913 (.I0(n2645), .I1(n30_adj_4823), .I2(n2639), 
            .I3(n2646), .O(n34_adj_4819));
    defparam i15_4_lut_adj_1913.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1914 (.I0(n2644), .I1(n2642_adj_4854), .I2(n2649), 
            .I3(n2643_adj_4853), .O(n32_adj_4821));
    defparam i13_4_lut_adj_1914.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1915 (.I0(n2637_adj_4856), .I1(n2636_adj_4857), 
            .I2(n2638_adj_4855), .I3(n2651), .O(n33_adj_4820));
    defparam i14_4_lut_adj_1915.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1916 (.I0(n2650), .I1(n2641), .I2(n35671), .I3(n2652), 
            .O(n31_adj_4822));
    defparam i12_4_lut_adj_1916.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1917 (.I0(n31_adj_4822), .I1(n33_adj_4820), .I2(n32_adj_4821), 
            .I3(n34_adj_4819), .O(n2669));
    defparam i18_4_lut_adj_1917.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1533_3_lut_3_lut (.I0(n2288), .I1(n6065), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12669_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n30070), .I3(GND_net), .O(n17398));   // verilog/coms.v(126[12] 292[6])
    defparam i12669_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1522_3_lut_3_lut (.I0(n2288), .I1(n6054), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12670_3_lut (.I0(encoder0_position[0]), .I1(n3018), .I2(count_enable), 
            .I3(GND_net), .O(n17399));   // quad.v(35[10] 41[6])
    defparam i12670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1918 (.I0(\FRAME_MATCHER.i_31__N_2621 ), .I1(\FRAME_MATCHER.i_31__N_2625 ), 
            .I2(n788), .I3(n2957_adj_4678), .O(n6_adj_4848));   // verilog/coms.v(126[12] 292[6])
    defparam i2_4_lut_adj_1918.LUT_INIT = 16'h0ace;
    SB_LUT4 div_46_i637_3_lut_3_lut (.I0(n938), .I1(n5895), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1919 (.I0(n63), .I1(\FRAME_MATCHER.state_31__N_2661 [0]), 
            .I2(n5_adj_4852), .I3(n6_adj_4848), .O(n34067));   // verilog/coms.v(126[12] 292[6])
    defparam i1_4_lut_adj_1919.LUT_INIT = 16'hddd5;
    SB_LUT4 i12672_3_lut (.I0(encoder1_position[0]), .I1(n2968), .I2(count_enable_adj_4701), 
            .I3(GND_net), .O(n17401));   // quad.v(35[10] 41[6])
    defparam i12672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12673_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n35976), 
            .I3(GND_net), .O(n17402));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12674_2_lut (.I0(r_SM_Main[2]), .I1(n43211), .I2(GND_net), 
            .I3(GND_net), .O(n17403));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12674_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_46_i1525_3_lut_3_lut (.I0(n2288), .I1(n6057), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4770), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i638_3_lut_3_lut (.I0(n938), .I1(n5896), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1523_3_lut_3_lut (.I0(n2288), .I1(n6055), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i639_3_lut_3_lut (.I0(n938), .I1(n5897), .I2(n652), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i636_3_lut_3_lut (.I0(n938), .I1(n5894), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1526_3_lut_3_lut (.I0(n2288), .I1(n6058), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i635_3_lut_3_lut (.I0(n938), .I1(n5893), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i634_3_lut_3_lut (.I0(n938), .I1(n5892), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4956));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33579_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n40409));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33579_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i723_3_lut_3_lut (.I0(n1067), .I1(n5904), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i724_3_lut_3_lut (.I0(n1067), .I1(n5905), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i725_3_lut_3_lut (.I0(n1067), .I1(n5906), .I2(n653), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i722_3_lut_3_lut (.I0(n1067), .I1(n5903), .I2(n1046), 
            .I3(GND_net), .O(n1172_adj_4751));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i721_3_lut_3_lut (.I0(n1067), .I1(n5902), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i720_3_lut_3_lut (.I0(n1067), .I1(n5901), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i719_3_lut_3_lut (.I0(n1067), .I1(n5900), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4959));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33571_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n40401));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33571_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1535_3_lut_3_lut (.I0(n2288), .I1(n6067), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i807_3_lut_3_lut (.I0(n1193), .I1(n5914), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i809_3_lut_3_lut (.I0(n1193), .I1(n5916), .I2(n654), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i808_3_lut_3_lut (.I0(n1193), .I1(n5915), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1593_3_lut_3_lut (.I0(n2381), .I1(n6084), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i805_3_lut_3_lut (.I0(n1193), .I1(n5912), .I2(n1172_adj_4751), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i803_3_lut_3_lut (.I0(n1193), .I1(n5910), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i804_3_lut_3_lut (.I0(n1193), .I1(n5911), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_5152));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12681_3_lut (.I0(tx_o), .I1(n3_adj_5264), .I2(r_SM_Main_adj_5379[2]), 
            .I3(GND_net), .O(n17410));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33476_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n40306));
    defparam i33476_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i806_3_lut_3_lut (.I0(n1193), .I1(n5913), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1532_3_lut_3_lut (.I0(n2288), .I1(n6064), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12682_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5379[1]), .I2(n8936), 
            .I3(n4_adj_4677), .O(n17411));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12682_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 div_46_i802_3_lut_3_lut (.I0(n1193), .I1(n5909), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12683_4_lut (.I0(r_SM_Main_adj_5379[2]), .I1(n10627), .I2(r_SM_Main_2__N_3579[1]), 
            .I3(r_SM_Main_adj_5379[0]), .O(n17412));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12683_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i12684_3_lut (.I0(quadB_debounced_adj_4700), .I1(reg_B_adj_5390[0]), 
            .I2(n35775), .I3(GND_net), .O(n17413));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12688_3_lut (.I0(setpoint[0]), .I1(n4349), .I2(n36881), .I3(GND_net), 
            .O(n17417));   // verilog/coms.v(126[12] 292[6])
    defparam i12688_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12695_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1172), .I3(GND_net), .O(n17424));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12696_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4736), 
            .I3(n15734), .O(n17425));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12696_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12697_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n15626), 
            .I3(n4_adj_4736), .O(n17426));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12697_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12698_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4704), 
            .I3(n15734), .O(n17427));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12698_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12699_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n15626), 
            .I3(n4_adj_4704), .O(n17428));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12699_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_5154));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12700_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4713), 
            .I3(n15734), .O(n17429));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12700_4_lut.LUT_INIT = 16'hccca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n18003(n18003), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n18004(n18004), .n18005(n18005), .n18006(n18006), 
            .n18007(n18007), .n18008(n18008), .n18009(n18009), .n18010(n18010), 
            .n18011(n18011), .n18012(n18012), .n18001(n18001), .n18002(n18002), 
            .n17999(n17999), .n18000(n18000), .n17997(n17997), .n17998(n17998), 
            .n17995(n17995), .n17996(n17996), .n17993(n17993), .n17994(n17994), 
            .n17990(n17990), .n17991(n17991), .n17992(n17992), .data_o({quadA_debounced_adj_4699, 
            quadB_debounced_adj_4700}), .GND_net(GND_net), .n2944({n2945, 
            n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
            n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
            n2962, n2963, n2964, n2965, n2966, n2967, n2968}), 
            .count_enable(count_enable_adj_4701), .n17401(n17401), .n18036(n18036), 
            .PIN_6_c_1(PIN_6_c_1), .reg_B({reg_B_adj_5390}), .n35775(n35775), 
            .n17413(n17413), .PIN_7_c_0(PIN_7_c_0)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(262[15] 267[4])
    SB_LUT4 i12702_4_lut (.I0(n35420), .I1(state[1]), .I2(state_3__N_362[1]), 
            .I3(n17008), .O(n17431));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12702_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 div_46_i1531_3_lut_3_lut (.I0(n2288), .I1(n6063), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4964));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_5156));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33455_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n40285));
    defparam i33455_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_5158));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_5176));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_5180));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34029_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n40861));
    defparam i34029_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_5182));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_5178));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33560_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n40390));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33560_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i34084_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n40916));
    defparam i34084_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1530_3_lut_3_lut (.I0(n2288), .I1(n6062), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_5198));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i890_3_lut_3_lut (.I0(n1316), .I1(n5926), .I2(n1299), 
            .I3(GND_net), .O(n1419_adj_4754));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_5202));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33911_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n40743));
    defparam i33911_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_5204));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_5200));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33952_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n40784));
    defparam i33952_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1529_3_lut_3_lut (.I0(n2288), .I1(n6061), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13317_3_lut (.I0(setpoint[9]), .I1(n4358), .I2(n36881), .I3(GND_net), 
            .O(n18046));   // verilog/coms.v(126[12] 292[6])
    defparam i13317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1528_3_lut_3_lut (.I0(n2288), .I1(n6060), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1524_3_lut_3_lut (.I0(n2288), .I1(n6056), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1539_3_lut_3_lut (.I0(n2288), .I1(n6071), .I2(n664), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i889_3_lut_3_lut (.I0(n1316), .I1(n5925), .I2(n1298), 
            .I3(GND_net), .O(n1418_adj_4753));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i891_3_lut_3_lut (.I0(n1316), .I1(n5927), .I2(n655), 
            .I3(GND_net), .O(n1420_adj_4755));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i887_3_lut_3_lut (.I0(n1316), .I1(n5923), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i886_3_lut_3_lut (.I0(n1316), .I1(n5922), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i888_3_lut_3_lut (.I0(n1316), .I1(n5924), .I2(n1297), 
            .I3(GND_net), .O(n1417_adj_4752));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i885_3_lut_3_lut (.I0(n1316), .I1(n5921), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i883_3_lut_3_lut (.I0(n1316), .I1(n5919), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i884_3_lut_3_lut (.I0(n1316), .I1(n5920), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1534_3_lut_3_lut (.I0(n2288), .I1(n6066), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33500_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n40330));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33500_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4968));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13337_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1172), .I3(GND_net), .O(n18066));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1527_3_lut_3_lut (.I0(n2288), .I1(n6059), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1538_3_lut_3_lut (.I0(n2288), .I1(n6070), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i970_3_lut_3_lut (.I0(n1436), .I1(n5938), .I2(n1420_adj_4755), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i964_3_lut_3_lut (.I0(n1436), .I1(n5932), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i968_3_lut_3_lut (.I0(n1436), .I1(n5936), .I2(n1418_adj_4753), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i969_3_lut_3_lut (.I0(n1436), .I1(n5937), .I2(n1419_adj_4754), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i967_3_lut_3_lut (.I0(n1436), .I1(n5935), .I2(n1417_adj_4752), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i963_3_lut_3_lut (.I0(n1436), .I1(n5931), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n34675), 
            .I2(n3894), .I3(n5_adj_5312), .O(n5_adj_4852));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff08;
    SB_LUT4 div_46_i971_3_lut_3_lut (.I0(n1436), .I1(n5939), .I2(n656), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1537_3_lut_3_lut (.I0(n2288), .I1(n6069), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i966_3_lut_3_lut (.I0(n1436), .I1(n5934), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1536_3_lut_3_lut (.I0(n2288), .I1(n6068), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i965_3_lut_3_lut (.I0(n1436), .I1(n5933), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i962_3_lut_3_lut (.I0(n1436), .I1(n5930), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33486_3_lut_4_lut (.I0(n1418_adj_4753), .I1(n97), .I2(n98), 
            .I3(n1419_adj_4754), .O(n40316));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33486_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_906_i34_3_lut_3_lut (.I0(n1418_adj_4753), .I1(n97), 
            .I2(n98), .I3(GND_net), .O(n34_adj_4977));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1047_3_lut_3_lut (.I0(n1553), .I1(n5950), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1045_3_lut_3_lut (.I0(n1553), .I1(n5948), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1048_3_lut_3_lut (.I0(n1553), .I1(n5951), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1042_3_lut_3_lut (.I0(n1553), .I1(n5945), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1049_3_lut_3_lut (.I0(n1553), .I1(n5952), .I2(n657), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1041_3_lut_3_lut (.I0(n1553), .I1(n5944), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1044_3_lut_3_lut (.I0(n1553), .I1(n5947), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1043_3_lut_3_lut (.I0(n1553), .I1(n5946), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1040_3_lut_3_lut (.I0(n1553), .I1(n5943), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1039_3_lut_3_lut (.I0(n1553), .I1(n5942), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1046_3_lut_3_lut (.I0(n1553), .I1(n5949), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36254_1_lut_2_lut (.I0(n3362), .I1(n10194), .I2(GND_net), 
            .I3(GND_net), .O(n43086));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36254_1_lut_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_46_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15845), 
            .O(n249));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1920 (.I0(n98), .I1(n97), .I2(n96), .I3(n15788), 
            .O(n15845));
    defparam i1_2_lut_4_lut_adj_1920.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1921 (.I0(n97), .I1(n96), .I2(n15788), 
            .I3(GND_net), .O(n15774));
    defparam i1_2_lut_3_lut_adj_1921.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_3_lut_4_lut (.I0(n855), .I1(n884), .I2(n956), .I3(n958), 
            .O(n35529));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1922 (.I0(n95), .I1(n94), .I2(n93), .I3(n15851), 
            .O(n15788));
    defparam i1_2_lut_4_lut_adj_1922.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1923 (.I0(n94), .I1(n93), .I2(n15851), 
            .I3(GND_net), .O(n15791));
    defparam i1_2_lut_3_lut_adj_1923.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4925));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1592_3_lut_3_lut (.I0(n2381), .I1(n6083), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1924 (.I0(n92), .I1(n91), .I2(n90), .I3(n15854), 
            .O(n15851));
    defparam i1_2_lut_4_lut_adj_1924.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1591_3_lut_3_lut (.I0(n2381), .I1(n6082), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1925 (.I0(n91), .I1(n90), .I2(n15854), 
            .I3(GND_net), .O(n15797));
    defparam i1_2_lut_3_lut_adj_1925.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1926 (.I0(n89), .I1(n88), .I2(n87), .I3(n15808), 
            .O(n15854));
    defparam i1_2_lut_4_lut_adj_1926.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1927 (.I0(n88), .I1(n87), .I2(n15808), 
            .I3(GND_net), .O(n15804));
    defparam i1_2_lut_3_lut_adj_1927.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1928 (.I0(n86), .I1(n85), .I2(n84), .I3(n15812), 
            .O(n15808));
    defparam i1_2_lut_4_lut_adj_1928.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6167), 
            .I3(n2724), .O(n41_adj_5244));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6168), 
            .I3(n2724), .O(n39_adj_5242));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4735), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n670));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6165), 
            .I3(n2724), .O(n45_adj_5246));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6166), 
            .I3(n2724), .O(n43_adj_5245));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6169), 
            .I3(n2724), .O(n37_adj_5241));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6173), 
            .I3(n2724), .O(n29_adj_5236));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6172), 
            .I3(n2724), .O(n31_adj_5238));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6177), 
            .I3(n2724), .O(n21_adj_5231));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6176), 
            .I3(n2724), .O(n23_adj_5232));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6175), 
            .I3(n2724), .O(n25_adj_5234));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6179), 
            .I3(n2724), .O(n17_adj_5229));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6178), 
            .I3(n2724), .O(n19_adj_5230));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6183), 
            .I3(n2724), .O(n9_adj_5222));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6170), 
            .I3(n2724), .O(n35_adj_5240));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6171), 
            .I3(n2724), .O(n33_adj_5239));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6184), 
            .I3(n2724), .O(n7_adj_5220));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6182), 
            .I3(n2724), .O(n11_adj_5224));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6181), 
            .I3(n2724), .O(n13_adj_5226));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6180), 
            .I3(n2724), .O(n15_adj_5227));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6174), 
            .I3(n2724), .O(n27_adj_5235));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33734_4_lut (.I0(n27_adj_5235), .I1(n15_adj_5227), .I2(n13_adj_5226), 
            .I3(n11_adj_5224), .O(n40564));
    defparam i33734_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_5239), 
            .I3(GND_net), .O(n12_adj_5225));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33659_2_lut (.I0(n33_adj_5239), .I1(n15_adj_5227), .I2(GND_net), 
            .I3(GND_net), .O(n40489));
    defparam i33659_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_5226), 
            .I3(GND_net), .O(n10_adj_5223));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i30_3_lut (.I0(n12_adj_5225), .I1(n83), 
            .I2(n35_adj_5240), .I3(GND_net), .O(n30_adj_5237));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1828_3_lut (.I0(n2720), .I1(n6185), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33836_3_lut (.I0(n7_adj_5220), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n40668));
    defparam i33836_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i34485_4_lut (.I0(n13_adj_5226), .I1(n11_adj_5224), .I2(n9_adj_5222), 
            .I3(n40668), .O(n41317));
    defparam i34485_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34475_4_lut (.I0(n19_adj_5230), .I1(n17_adj_5229), .I2(n15_adj_5227), 
            .I3(n41317), .O(n41307));
    defparam i34475_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35329_4_lut (.I0(n25_adj_5234), .I1(n23_adj_5232), .I2(n21_adj_5231), 
            .I3(n41307), .O(n42161));
    defparam i35329_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34829_4_lut (.I0(n31_adj_5238), .I1(n29_adj_5236), .I2(n27_adj_5235), 
            .I3(n42161), .O(n41661));
    defparam i34829_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35431_4_lut (.I0(n37_adj_5241), .I1(n35_adj_5240), .I2(n33_adj_5239), 
            .I3(n41661), .O(n42263));
    defparam i35431_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_5245), 
            .I3(GND_net), .O(n16_adj_5228));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_5220), 
            .I3(GND_net), .O(n6_adj_5219));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i35019_3_lut (.I0(n6_adj_5219), .I1(n90), .I2(n21_adj_5231), 
            .I3(GND_net), .O(n41851));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35019_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35020_3_lut (.I0(n41851), .I1(n89), .I2(n23_adj_5232), .I3(GND_net), 
            .O(n41852));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35020_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33765_4_lut (.I0(n21_adj_5231), .I1(n19_adj_5230), .I2(n17_adj_5229), 
            .I3(n9_adj_5222), .O(n40596));
    defparam i33765_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33621_2_lut (.I0(n43_adj_5245), .I1(n19_adj_5230), .I2(GND_net), 
            .I3(GND_net), .O(n40451));
    defparam i33621_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_5229), 
            .I3(GND_net), .O(n8_adj_5221));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i24_3_lut (.I0(n16_adj_5228), .I1(n78), 
            .I2(n45_adj_5246), .I3(GND_net), .O(n24_adj_5233));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33625_4_lut (.I0(n43_adj_5245), .I1(n25_adj_5234), .I2(n23_adj_5232), 
            .I3(n40596), .O(n40455));
    defparam i33625_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34859_4_lut (.I0(n24_adj_5233), .I1(n8_adj_5221), .I2(n45_adj_5246), 
            .I3(n40451), .O(n41691));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34859_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34440_3_lut (.I0(n41852), .I1(n88), .I2(n25_adj_5234), .I3(GND_net), 
            .O(n41272));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34440_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1829_3_lut (.I0(n669), .I1(n6186), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i4_4_lut (.I0(n670), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_5218));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35189_3_lut (.I0(n4_adj_5218), .I1(n87), .I2(n27_adj_5235), 
            .I3(GND_net), .O(n42021));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35189_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35190_3_lut (.I0(n42021), .I1(n86), .I2(n29_adj_5236), .I3(GND_net), 
            .O(n42022));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35190_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33699_4_lut (.I0(n33_adj_5239), .I1(n31_adj_5238), .I2(n29_adj_5236), 
            .I3(n40564), .O(n40529));
    defparam i33699_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35455_4_lut (.I0(n30_adj_5237), .I1(n10_adj_5223), .I2(n35_adj_5240), 
            .I3(n40489), .O(n42287));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35455_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35142_3_lut (.I0(n42022), .I1(n85), .I2(n31_adj_5238), .I3(GND_net), 
            .O(n41974));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35142_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35554_4_lut (.I0(n41974), .I1(n42287), .I2(n35_adj_5240), 
            .I3(n40529), .O(n42386));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35554_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35555_3_lut (.I0(n42386), .I1(n82), .I2(n37_adj_5241), .I3(GND_net), 
            .O(n42387));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35555_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35521_3_lut (.I0(n42387), .I1(n81), .I2(n39_adj_5242), .I3(GND_net), 
            .O(n42353));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35521_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33627_4_lut (.I0(n43_adj_5245), .I1(n41_adj_5244), .I2(n39_adj_5242), 
            .I3(n42263), .O(n40457));
    defparam i33627_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35323_4_lut (.I0(n41272), .I1(n41691), .I2(n45_adj_5246), 
            .I3(n40455), .O(n42155));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35323_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35502_3_lut (.I0(n42353), .I1(n80), .I2(n41_adj_5244), .I3(GND_net), 
            .O(n40_adj_5243));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35502_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1807_3_lut (.I0(n2699), .I1(n6164), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35325_4_lut (.I0(n40_adj_5243), .I1(n42155), .I2(n45_adj_5246), 
            .I3(n40457), .O(n42157));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35325_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35326_3_lut (.I0(n42157), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35326_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1929 (.I0(n85), .I1(n84), .I2(n15812), 
            .I3(GND_net), .O(n15860));
    defparam i1_2_lut_3_lut_adj_1929.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1930 (.I0(n83), .I1(n82), .I2(n81), .I3(n15866), 
            .O(n15812));
    defparam i1_2_lut_4_lut_adj_1930.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1931 (.I0(n82), .I1(n81), .I2(n15866), 
            .I3(GND_net), .O(n15880));
    defparam i1_2_lut_3_lut_adj_1931.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1932 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n15866));
    defparam i1_2_lut_4_lut_adj_1932.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1933 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n15871));
    defparam i1_2_lut_3_lut_adj_1933.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5215));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22645_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n511), .I3(n558), 
            .O(n4_adj_5309));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22645_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5213));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22669_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n650), .I3(n558), 
            .O(n4_adj_5306));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22669_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5217));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5216));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4728), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n669));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5210));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5211));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22701_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n651), .I3(n558), 
            .O(n4_adj_4689));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22701_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5208));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5209));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5199));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5201));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5207));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4984));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5203));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5205));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5206));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5212));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33932_4_lut (.I0(n29_adj_5212), .I1(n17_adj_5206), .I2(n15_adj_5205), 
            .I3(n13_adj_5203), .O(n40764));
    defparam i33932_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34603_4_lut (.I0(n11_adj_5201), .I1(n9_adj_5199), .I2(n2719), 
            .I3(n98), .O(n41435));
    defparam i34603_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34937_4_lut (.I0(n17_adj_5206), .I1(n15_adj_5205), .I2(n13_adj_5203), 
            .I3(n41435), .O(n41769));
    defparam i34937_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34925_4_lut (.I0(n23_adj_5209), .I1(n21_adj_5208), .I2(n19_adj_5207), 
            .I3(n41769), .O(n41757));
    defparam i34925_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33938_4_lut (.I0(n29_adj_5212), .I1(n27_adj_5211), .I2(n25_adj_5210), 
            .I3(n41757), .O(n40770));
    defparam i33938_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1777_i6_4_lut (.I0(n669), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_5197));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35023_3_lut (.I0(n6_adj_5197), .I1(n87), .I2(n29_adj_5212), 
            .I3(GND_net), .O(n41855));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35023_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1777_i32_3_lut (.I0(n14_adj_5204), .I1(n83), 
            .I2(n37_adj_5217), .I3(GND_net), .O(n32_adj_5214));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35024_3_lut (.I0(n41855), .I1(n86), .I2(n31_adj_5213), .I3(GND_net), 
            .O(n41856));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35024_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33916_4_lut (.I0(n35_adj_5216), .I1(n33_adj_5215), .I2(n31_adj_5213), 
            .I3(n40764), .O(n40748));
    defparam i33916_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35387_4_lut (.I0(n32_adj_5214), .I1(n12_adj_5202), .I2(n37_adj_5217), 
            .I3(n40743), .O(n42219));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35387_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34432_3_lut (.I0(n41856), .I1(n85), .I2(n33_adj_5215), .I3(GND_net), 
            .O(n41264));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34432_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35025_3_lut (.I0(n8_adj_5198), .I1(n90), .I2(n23_adj_5209), 
            .I3(GND_net), .O(n41857));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35025_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35026_3_lut (.I0(n41857), .I1(n89), .I2(n25_adj_5210), .I3(GND_net), 
            .O(n41858));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35026_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34563_4_lut (.I0(n25_adj_5210), .I1(n23_adj_5209), .I2(n21_adj_5208), 
            .I3(n40784), .O(n41395));
    defparam i34563_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34857_3_lut (.I0(n10_adj_5200), .I1(n91), .I2(n21_adj_5208), 
            .I3(GND_net), .O(n41689));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34857_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34430_3_lut (.I0(n41858), .I1(n88), .I2(n27_adj_5211), .I3(GND_net), 
            .O(n41262));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34430_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35163_4_lut (.I0(n35_adj_5216), .I1(n33_adj_5215), .I2(n31_adj_5213), 
            .I3(n40770), .O(n41995));
    defparam i35163_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35503_4_lut (.I0(n41264), .I1(n42219), .I2(n37_adj_5217), 
            .I3(n40748), .O(n42335));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35503_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35193_4_lut (.I0(n41262), .I1(n41689), .I2(n27_adj_5211), 
            .I3(n41395), .O(n42025));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35193_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_i1121_3_lut_3_lut (.I0(n1667), .I1(n5962), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35566_4_lut (.I0(n42025), .I1(n42335), .I2(n37_adj_5217), 
            .I3(n41995), .O(n42398));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35566_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35567_3_lut (.I0(n42398), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n42399));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35567_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35565_3_lut (.I0(n42399), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n42397));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35565_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35335_3_lut (.I0(n42397), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n42167));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35335_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i1123_3_lut_3_lut (.I0(n1667), .I1(n5964), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35336_3_lut (.I0(n42167), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n42168));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35336_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i2010_4_lut (.I0(n42168), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i2010_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1118_3_lut_3_lut (.I0(n1667), .I1(n5959), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1124_3_lut_3_lut (.I0(n1667), .I1(n5965), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34128_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n40960));
    defparam i34128_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1117_3_lut_3_lut (.I0(n1667), .I1(n5958), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4986));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4997));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1125_3_lut_3_lut (.I0(n1667), .I1(n5966), .I2(n658), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1120_3_lut_3_lut (.I0(n1667), .I1(n5961), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34099_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n40931));
    defparam i34099_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5194));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4999));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1119_3_lut_3_lut (.I0(n1667), .I1(n5960), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5196));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1116_3_lut_3_lut (.I0(n1667), .I1(n5957), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1115_3_lut_3_lut (.I0(n1667), .I1(n5956), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1114_3_lut_3_lut (.I0(n1667), .I1(n5955), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5192));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4729), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n668));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1590_3_lut_3_lut (.I0(n2381), .I1(n6081), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_5009));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5195));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34044_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n40876));
    defparam i34044_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_5011));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5189));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5190));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34020_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n40852));
    defparam i34020_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_5025));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5187));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5188));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_5021));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5177));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34009_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n40841));
    defparam i34009_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_5023));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5179));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5186));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_5036));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33954_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n40786));
    defparam i33954_2_lut_4_lut.LUT_INIT = 16'hf99f;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n17983(n17983), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n17984(n17984), .n17985(n17985), .n17986(n17986), 
            .n17987(n17987), .n17988(n17988), .n17975(n17975), .n17976(n17976), 
            .n17977(n17977), .n17978(n17978), .n17979(n17979), .n17980(n17980), 
            .n17981(n17981), .n17982(n17982), .n17971(n17971), .n17972(n17972), 
            .n17973(n17973), .n17974(n17974), .n17966(n17966), .n17967(n17967), 
            .n17968(n17968), .n17969(n17969), .n17970(n17970), .data_o({quadA_debounced, 
            quadB_debounced}), .count_enable(count_enable), .n17399(n17399), 
            .n2994({n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
            n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
            n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
            n3018}), .GND_net(GND_net), .n18020(n18020), .reg_B({reg_B}), 
            .n35976(n35976), .PIN_2_c_0(PIN_2_c_0), .n17402(n17402), .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(254[15] 259[4])
    SB_LUT4 div_46_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5181));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5184));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5191));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1122_3_lut_3_lut (.I0(n1667), .I1(n5963), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34047_4_lut (.I0(n31_adj_5191), .I1(n19_adj_5184), .I2(n17_adj_5183), 
            .I3(n15_adj_5181), .O(n40879));
    defparam i34047_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34691_4_lut (.I0(n13_adj_5179), .I1(n11_adj_5177), .I2(n2637), 
            .I3(n98), .O(n41523));
    defparam i34691_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34977_4_lut (.I0(n19_adj_5184), .I1(n17_adj_5183), .I2(n15_adj_5181), 
            .I3(n41523), .O(n41809));
    defparam i34977_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34975_4_lut (.I0(n25_adj_5188), .I1(n23_adj_5187), .I2(n21_adj_5186), 
            .I3(n41809), .O(n41807));
    defparam i34975_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34049_4_lut (.I0(n31_adj_5191), .I1(n29_adj_5190), .I2(n27_adj_5189), 
            .I3(n41807), .O(n40881));
    defparam i34049_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1722_i8_4_lut (.I0(n668), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_5175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35029_3_lut (.I0(n8_adj_5175), .I1(n87), .I2(n31_adj_5191), 
            .I3(GND_net), .O(n41861));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35029_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35030_3_lut (.I0(n41861), .I1(n86), .I2(n33_adj_5192), .I3(GND_net), 
            .O(n41862));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35030_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1722_i34_3_lut (.I0(n16_adj_5182), .I1(n83), 
            .I2(n39_adj_5196), .I3(GND_net), .O(n34_adj_5193));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34033_4_lut (.I0(n37_adj_5195), .I1(n35_adj_5194), .I2(n33_adj_5192), 
            .I3(n40879), .O(n40865));
    defparam i34033_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35385_4_lut (.I0(n34_adj_5193), .I1(n14_adj_5180), .I2(n39_adj_5196), 
            .I3(n40861), .O(n42217));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35385_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34422_3_lut (.I0(n41862), .I1(n85), .I2(n35_adj_5194), .I3(GND_net), 
            .O(n41254));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34422_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35031_3_lut (.I0(n10_adj_5176), .I1(n90), .I2(n25_adj_5188), 
            .I3(GND_net), .O(n41863));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35031_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35032_3_lut (.I0(n41863), .I1(n89), .I2(n27_adj_5189), .I3(GND_net), 
            .O(n41864));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35032_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34671_4_lut (.I0(n27_adj_5189), .I1(n25_adj_5188), .I2(n23_adj_5187), 
            .I3(n40916), .O(n41503));
    defparam i34671_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1722_i20_3_lut (.I0(n12_adj_5178), .I1(n91), 
            .I2(n23_adj_5187), .I3(GND_net), .O(n20_adj_5185));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34420_3_lut (.I0(n41864), .I1(n88), .I2(n29_adj_5190), .I3(GND_net), 
            .O(n41252));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34420_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35181_4_lut (.I0(n37_adj_5195), .I1(n35_adj_5194), .I2(n33_adj_5192), 
            .I3(n40881), .O(n42013));
    defparam i35181_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35536_4_lut (.I0(n41254), .I1(n42217), .I2(n39_adj_5196), 
            .I3(n40865), .O(n42368));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35536_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34855_4_lut (.I0(n41252), .I1(n20_adj_5185), .I2(n29_adj_5190), 
            .I3(n41503), .O(n41687));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34855_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35558_4_lut (.I0(n41687), .I1(n42368), .I2(n39_adj_5196), 
            .I3(n42013), .O(n42390));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35558_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35559_3_lut (.I0(n42390), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n42391));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35559_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35195_3_lut (.I0(n42391), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n42027));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35195_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35196_3_lut (.I0(n42027), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n42028));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35196_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1934 (.I0(n42028), .I1(n15817), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1934.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_5038));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33966_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n40798));
    defparam i33966_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_5040));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_5053));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33902_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n40734));
    defparam i33902_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_5055));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33914_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n40746));
    defparam i33914_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_5057));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4730), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n667));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_5070));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33797_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n40629));
    defparam i33797_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_5072));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1589_3_lut_3_lut (.I0(n2381), .I1(n6080), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5165));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5167));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_5074));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33822_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n40654));
    defparam i33822_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5153));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5155));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5162));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5163));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5164));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_5090));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5168));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33686_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n40516));
    defparam i33686_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_5092));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5157));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5159));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5160));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33466_4_lut (.I0(n33_adj_5168), .I1(n21_adj_5160), .I2(n19_adj_5159), 
            .I3(n17_adj_5157), .O(n40296));
    defparam i33466_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34197_4_lut (.I0(n15_adj_5155), .I1(n13_adj_5153), .I2(n2552), 
            .I3(n98), .O(n41029));
    defparam i34197_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34743_4_lut (.I0(n21_adj_5160), .I1(n19_adj_5159), .I2(n17_adj_5157), 
            .I3(n41029), .O(n41575));
    defparam i34743_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34741_4_lut (.I0(n27_adj_5164), .I1(n25_adj_5163), .I2(n23_adj_5162), 
            .I3(n41575), .O(n41573));
    defparam i34741_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33468_4_lut (.I0(n33_adj_5168), .I1(n31_adj_5167), .I2(n29_adj_5165), 
            .I3(n41573), .O(n40298));
    defparam i33468_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1665_i10_4_lut (.I0(n667), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_5151));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35197_3_lut (.I0(n10_adj_5151), .I1(n87), .I2(n33_adj_5168), 
            .I3(GND_net), .O(n42029));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35197_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35198_3_lut (.I0(n42029), .I1(n86), .I2(n35_adj_5170), .I3(GND_net), 
            .O(n42030));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35198_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i36_3_lut (.I0(n18_adj_5158), .I1(n83), 
            .I2(n41_adj_5174), .I3(GND_net), .O(n36_adj_5171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33460_4_lut (.I0(n39_adj_5173), .I1(n37_adj_5172), .I2(n35_adj_5170), 
            .I3(n40296), .O(n40290));
    defparam i33460_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35383_4_lut (.I0(n36_adj_5171), .I1(n16_adj_5156), .I2(n41_adj_5174), 
            .I3(n40285), .O(n42215));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35383_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35136_3_lut (.I0(n42030), .I1(n85), .I2(n37_adj_5172), .I3(GND_net), 
            .O(n34_adj_5169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35136_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i22_3_lut (.I0(n14_adj_5154), .I1(n91), 
            .I2(n25_adj_5163), .I3(GND_net), .O(n22_adj_5161));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35452_4_lut (.I0(n22_adj_5161), .I1(n12_adj_5152), .I2(n25_adj_5163), 
            .I3(n40306), .O(n42284));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35452_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35453_3_lut (.I0(n42284), .I1(n90), .I2(n27_adj_5164), .I3(GND_net), 
            .O(n42285));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35453_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35338_3_lut (.I0(n42285), .I1(n89), .I2(n29_adj_5165), .I3(GND_net), 
            .O(n42170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35338_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35001_4_lut (.I0(n39_adj_5173), .I1(n37_adj_5172), .I2(n35_adj_5170), 
            .I3(n40298), .O(n41833));
    defparam i35001_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35475_4_lut (.I0(n34_adj_5169), .I1(n42215), .I2(n41_adj_5174), 
            .I3(n40290), .O(n42307));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35475_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35318_3_lut (.I0(n42170), .I1(n88), .I2(n31_adj_5167), .I3(GND_net), 
            .O(n30_adj_5166));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35318_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35562_4_lut (.I0(n30_adj_5166), .I1(n42307), .I2(n41_adj_5174), 
            .I3(n41833), .O(n42394));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35562_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35563_3_lut (.I0(n42394), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n42395));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35563_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35561_3_lut (.I0(n42395), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n42393));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35561_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1935 (.I0(n42393), .I1(n15871), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1935.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1597_3_lut_3_lut (.I0(n2381), .I1(n6088), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_5094));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33701_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n40531));
    defparam i33701_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_5108));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5148));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33597_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n40427));
    defparam i33597_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1595_3_lut_3_lut (.I0(n2381), .I1(n6086), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1198_3_lut_3_lut (.I0(n1778), .I1(n5980), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5146));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_5110));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1189_3_lut_3_lut (.I0(n1778), .I1(n5971), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5150));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_5112));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5149));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1583_3_lut_3_lut (.I0(n2381), .I1(n6074), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33540_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n40370));
    defparam i33540_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4731), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n666));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_5114));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1600_3_lut_3_lut (.I0(n2381), .I1(n6091), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1187_3_lut_3_lut (.I0(n1778), .I1(n5969), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1584_3_lut_3_lut (.I0(n2381), .I1(n6075), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1192_3_lut_3_lut (.I0(n1778), .I1(n5974), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5143));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5144));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    motorControl control (.duty({duty}), .GND_net(GND_net), .PWMLimit({PWMLimit}), 
            .\Kp[15] (Kp[15]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .\Kp[2] (Kp[2]), .\Kp[8] (Kp[8]), .\Kp[10] (Kp[10]), .clk32MHz(clk32MHz), 
            .\Kp[9] (Kp[9]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .VCC_net(VCC_net), .n25(n25), .IntegralLimit({IntegralLimit}), 
            .\Ki[3] (Ki[3]), .\Ki[2] (Ki[2]), .\Ki[0] (Ki[0]), .\Ki[1] (Ki[1]), 
            .n43164(n43164), .setpoint({setpoint}), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Ki[6] (Ki[6]), .motor_state({motor_state}), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
            .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15])) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(234[16] 247[4])
    SB_LUT4 div_46_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_5130));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1196_3_lut_3_lut (.I0(n1778), .I1(n5978), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33521_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n40351));
    defparam i33521_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5140));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1587_3_lut_3_lut (.I0(n2381), .I1(n6078), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5141));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5142));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1197_3_lut_3_lut (.I0(n1778), .I1(n5979), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_5132));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5131));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1195_3_lut_3_lut (.I0(n1778), .I1(n5977), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5133));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_5134));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33503_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n40333));
    defparam i33503_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_5136));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5135));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    \pwm(32000000,20000,32000000,23,1)  PWM (.pwm_setpoint({pwm_setpoint}), 
            .GND_net(GND_net), .\half_duty_new[0] (half_duty_new[0]), .CLK_c(CLK_c), 
            .PIN_19_c_0(PIN_19_c_0), .n18061(n18061), .\half_duty[0][1] (\half_duty[0] [1]), 
            .n18062(n18062), .\half_duty[0][2] (\half_duty[0] [2]), .n18063(n18063), 
            .\half_duty[0][3] (\half_duty[0] [3]), .n18064(n18064), .\half_duty[0][4] (\half_duty[0] [4]), 
            .n18066(n18066), .\half_duty[0][6] (\half_duty[0] [6]), .n18067(n18067), 
            .\half_duty[0][7] (\half_duty[0] [7]), .n1172(n1172), .VCC_net(VCC_net), 
            .\half_duty_new[1] (half_duty_new[1]), .\half_duty[0][0] (\half_duty[0] [0]), 
            .\half_duty_new[2] (half_duty_new[2]), .\half_duty_new[3] (half_duty_new[3]), 
            .\half_duty_new[4] (half_duty_new[4]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[7] (half_duty_new[7]), .n17424(n17424)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(153[43] 159[3])
    SB_LUT4 div_46_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5137));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1191_3_lut_3_lut (.I0(n1778), .I1(n5973), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5138));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5145));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33509_4_lut (.I0(n35_adj_5145), .I1(n23_adj_5138), .I2(n21_adj_5137), 
            .I3(n19_adj_5135), .O(n40339));
    defparam i33509_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34233_4_lut (.I0(n17_adj_5133), .I1(n15_adj_5131), .I2(n2464), 
            .I3(n98), .O(n41065));
    defparam i34233_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34759_4_lut (.I0(n23_adj_5138), .I1(n21_adj_5137), .I2(n19_adj_5135), 
            .I3(n41065), .O(n41591));
    defparam i34759_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34757_4_lut (.I0(n29_adj_5142), .I1(n27_adj_5141), .I2(n25_adj_5140), 
            .I3(n41591), .O(n41589));
    defparam i34757_4_lut.LUT_INIT = 16'hfeff;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, bit_ctr, VCC_net, 
            n40238, GND_net, n19, timer, n33435, n33465, n33467, 
            n33469, n33471, n33473, n33475, n33477, n33429, n33431, 
            n33443, n33445, n33451, n33453, n33455, n33457, n33497, 
            n33493, n33495, n33489, n33491, n33485, n33487, n33479, 
            n33481, n33483, n33463, n33461, n33433, \neo_pixel_transmitter.t0 , 
            n40237, n40231, \state_3__N_362[1] , \state[1] , n1166, 
            \state[0] , n4442, n40236, n40245, n40234, n24628, start, 
            n15744, \one_wire_N_513[10] , \one_wire_N_513[8] , \one_wire_N_513[5] , 
            \one_wire_N_513[11] , \one_wire_N_513[7] , \one_wire_N_513[9] , 
            \one_wire_N_513[6] , n35327, n33459, n33441, n33439, n17493, 
            n17492, n17491, n17490, n17489, n17488, n17487, n17486, 
            n17485, n17484, n17483, n17482, n17481, n17480, n17479, 
            n17478, n17477, n17476, n17475, n17474, n17473, n17472, 
            n17471, n17470, n17469, n17468, n17467, n17466, n17465, 
            n17464, n17463, n35462, n40230, n35424, n36115, n17431, 
            n40228, n17008, n35420, PIN_8_c, n36877, n40227, n11, 
            n40244, n33499, n17248, n40223, n40235, n40224, n40254, 
            n40253, n40252, n40251, n40226, n40225, n40250, n40249, 
            n40233, n40248, n40247, n40246, n40243, n40229, n40232, 
            n40242, n40241, n40240, n40239, \color[2] , \color[3] , 
            \color[4] , \color[1] , n24520) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output [31:0]bit_ctr;
    input VCC_net;
    output n40238;
    input GND_net;
    input n19;
    output [31:0]timer;
    input n33435;
    input n33465;
    input n33467;
    input n33469;
    input n33471;
    input n33473;
    input n33475;
    input n33477;
    input n33429;
    input n33431;
    input n33443;
    input n33445;
    input n33451;
    input n33453;
    input n33455;
    input n33457;
    input n33497;
    input n33493;
    input n33495;
    input n33489;
    input n33491;
    input n33485;
    input n33487;
    input n33479;
    input n33481;
    input n33483;
    input n33463;
    input n33461;
    input n33433;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output n40237;
    output n40231;
    output \state_3__N_362[1] ;
    output \state[1] ;
    output n1166;
    output \state[0] ;
    output n4442;
    output n40236;
    output n40245;
    output n40234;
    output n24628;
    output start;
    output n15744;
    output \one_wire_N_513[10] ;
    output \one_wire_N_513[8] ;
    output \one_wire_N_513[5] ;
    output \one_wire_N_513[11] ;
    output \one_wire_N_513[7] ;
    output \one_wire_N_513[9] ;
    output \one_wire_N_513[6] ;
    output n35327;
    input n33459;
    input n33441;
    input n33439;
    input n17493;
    input n17492;
    input n17491;
    input n17490;
    input n17489;
    input n17488;
    input n17487;
    input n17486;
    input n17485;
    input n17484;
    input n17483;
    input n17482;
    input n17481;
    input n17480;
    input n17479;
    input n17478;
    input n17477;
    input n17476;
    input n17475;
    input n17474;
    input n17473;
    input n17472;
    input n17471;
    input n17470;
    input n17469;
    input n17468;
    input n17467;
    input n17466;
    input n17465;
    input n17464;
    input n17463;
    input n35462;
    output n40230;
    output n35424;
    output n36115;
    input n17431;
    output n40228;
    output n17008;
    output n35420;
    output PIN_8_c;
    input n36877;
    output n40227;
    input n11;
    output n40244;
    input n33499;
    input n17248;
    output n40223;
    output n40235;
    output n40224;
    output n40254;
    output n40253;
    output n40252;
    output n40251;
    output n40226;
    output n40225;
    output n40250;
    output n40249;
    output n40233;
    output n40248;
    output n40247;
    output n40246;
    output n40243;
    output n40229;
    output n40232;
    output n40242;
    output n40241;
    output n40240;
    output n40239;
    input \color[2] ;
    input \color[3] ;
    input \color[4] ;
    input \color[1] ;
    output n24520;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n29297, n3090, n3116, n29298, n2408, n2309, n43140, n29098, 
        n29099, n3190, n3091, n29296, \neo_pixel_transmitter.done_N_570 , 
        n37261, n2409, n27764, n2291, n2192, n2225, n29097, n3191, 
        n3092, n29295, n2292, n2193, n29096;
    wire [31:0]one_wire_N_513;
    wire [31:0]n1;
    
    wire n28010, n3192, n3093, n29294, n2293, n2194, n29095, n3193, 
        n3094, n29293, n28011, n2294, n2195, n29094, n3194, n3095, 
        n29292, n2295, n2196, n29093, n3195, n3096, n29291, n2296, 
        n2197, n29092, n3196, n3097, n29290, n2297, n2198, n29091, 
        n3197, n3098, n29289, n2298, n2199, n29090, n3198, n3099, 
        n29288, n28009, n2299, n2200, n29089, n3199, n3100, n29287, 
        n2300, n2201, n29088, n3200, n3101, n29286, n2301, n2202, 
        n29087, n3201, n3102, n29285, n2302, n2203, n29086, n3202, 
        n3103, n29284, n2103, n2097, n18, n2109, n24514, n2093, 
        n2108, n2100, n30_adj_4539, n2098, n2094, n2099, n28, 
        n2105, n2096, n2095, n2102, n29, n2101, n2107, n2104, 
        n2106, n27, n2126, n43141, n2303, n2204, n29085, n3001, 
        n3002, n2994, n2991, n40, n2989, n2990, n2996, n3007, 
        n44, n3005, n3008, n2988, n2998, n42, n2986, n2995, 
        n2997, n2985, n43, n2984, n2992, n2993, n3003, n41, 
        n3006, n3009, n38, n3000, n2987, n46, n50, n2999, n3004, 
        n37, n3203, n3104, n29283, n3204, n3105, n29282, n3017, 
        n30079, n28008, n4, n3205, n3106, n29281, n3206, n3107, 
        n29280, n3207, n3108, n29279, n3208, n3109, n43139, n29278, 
        n3209, n2304, n2205, n29084, n3083, n29277, n2305, n2206, 
        n29083, n3084, n29276, n2306, n2207, n29082, n2307, n2208, 
        n29081, n1608, n1606, n1604, n1603, n20, n1602, n1609, 
        n13, n1598, n1600, n18_adj_4540, n1605, n1599, n22, n1601, 
        n1607, n1631, n3085, n29275, n2308, n2209, n29080, n3086, 
        n29274, n3087, n29273, n29079, n29078, n27765, n3088, 
        n29272, n3089, n29271, n29077, n29270, n29076, n29269, 
        n29268, n29267, n29266, n29075, n29074, n29265, n29264, 
        n29263, n29262, n29261, n29073, n29072, n29260, n29259, 
        n1730, n43151, n29071, n29070, n29069, n29068, n29067, 
        n27763, n29066, n30_adj_4541, n48, n46_adj_4542, n29258, 
        n29065, n27752, n29257, n29064, n29256, n29255, n43143, 
        n29063, n29254, n1994, n2027, n29062, n1995, n29061, n29253, 
        n43142, n29252, n1996, n29060, n47, n45, n1997, n29059, 
        n44_adj_4543, n43_adj_4544, n54, n49, n15745, n4414, n2885, 
        n2918, n29251, n2886, n29250, n1998, n29058, n2887, n29249, 
        n2888, n29248, n1999, n29057, n2889, n29247, n2000, n29056, 
        n2001, n29055, n2890, n29246;
    wire [31:0]n133;
    
    wire n28565, n2002, n29054, n2891, n29245, n28564, n28563, 
        n28562, n28561, n2892, n29244, n2003, n29053, n28560, 
        n28559, n2893, n29243, n2004, n29052, n2894, n29242, n2005, 
        n29051, n2895, n29241, n2006, n29050, n2896, n29240, n28558, 
        n2897, n29239, n2898, n29238, n2007, n29049, n28557, n2008, 
        n29048, n28556, n2009, n43144, n29047, n28555, n2899, 
        n29237, n2900, n29236, n28554, n1895, n1928, n29046, n28553, 
        n1896, n29045, n28552, n28551, n28550, n28549, n28548, 
        n28547, n28546, n28545, n28544, n28543, n28542, n27762, 
        n28541, n28540, n2901, n29235, n1897, n29044, n28539, 
        n28538, n1898, n29043, n28537, n1899, n29042, n2902, n29234, 
        n1900, n29041, n28536, n28535, n1901, n29040, n1902, n29039, 
        n2903, n29233, n1903, n29038, n1904, n29037, n2904, n29232, 
        n1905, n29036, n2905, n29231, n2906, n29230, n2907, n29229, 
        n1906, n29035, n2908, n29228, n1907, n29034, n27753, n2909, 
        n43145, n29227, n1908, n29033, n1909, n43146, n29032, 
        n2786, n2819, n29226, n2787, n29225, n2788, n29224, n1796, 
        n1829, n29031, n1797, n29030, n1798, n29029, n27751, n27761, 
        n2789, n29223, n2790, n29222, n2791, n29221, n2792, n29220, 
        n1799, n29028, n2793, n29219, n2794, n29218, n2795, n29217, 
        n1800, n29027, n2796, n29216, n2797, n29215, n2798, n29214, 
        n1801, n29026, n2799, n29213, n2800, n29212, n2801, n29211, 
        n1802, n29025, n1803, n29024, n2802, n29210, n2803, n29209, 
        n1804, n29023, n1805, n29022, n2804, n29208, n2805, n29207, 
        n1806, n29021, n2806, n29206, n1807, n29020, n2807, n29205, 
        n1808, n29019, n2808, n29204, n2809, n43148, n29203, n2687, 
        n2720, n29202, n2688, n29201, n2689, n29200, n1809, n43149, 
        n29018, n2690, n29199, n2691, n29198, n2692, n29197, n2693, 
        n29196, n1697, n29017, n2694, n29195, n1698, n29016, n2695, 
        n29194, n2696, n29193, n2697, n29192, n1699, n29015, n1700, 
        n29014, n2698, n29191, n1701, n29013, n1702, n29012, n2699, 
        n29190, n1703, n29011, n28_adj_4545, n32_adj_4546, n30_adj_4547, 
        n31_adj_4548, n29_adj_4549, n29824, n15631, n24324, n4_adj_4550, 
        n10, n15824, n14, n1704, n29010, n1506, n1503, n1500, 
        n1501, n18_adj_4551, n1504, n1502, n1499, n20_adj_4552, 
        n1505, n1509, n15, n1508, n1507, n1532, n27880, n21, 
        n23, n22_adj_4553, n24, n36, n25, n27_adj_4554, n26, n28_adj_4555, 
        n37_adj_4556, n29_adj_4557, n30_adj_4558, n34689, n35373, 
        n5, n34738, n116, n1705, n29009, n2700, n29189, n1706, 
        n29008, n2701, n29188, n27879, n1707, n29007, n27878, 
        n27877, n2702, n29187, n1708, n29006, n1709, n29005, n2703, 
        n29186, n27876, n2704, n29185, n29004, n2705, n29184, 
        n29003, n27875, n2706, n29183, n29002, n2707, n29182, 
        n29001, n27760, n2708, n29181, n29000, n27874, n2709, 
        n43150, n29180, n28999, n28998, n27873, n2588, n2621, 
        n29179, n28997, n27872, n2589, n29178, n28996, n27871, 
        n28995, n2590, n29177, n43153, n27870, n28994, n2591, 
        n29176, n35335, n36000, n35991, n2592, n29175, n2593, 
        n29174, n43154, n28993, n2594, n29173, n2595, n29172, 
        n27759, n2596, n29171, n2597, n29170, n2598, n29169, n2599, 
        n29168;
    wire [3:0]state_3__N_362;
    
    wire \neo_pixel_transmitter.done_N_576 , n16961, n35303, n14348, 
        n807, n838, n35416, n35313, n2600, n29167, n2601, n29166, 
        n2423, n43162, n2602, n29165, n2603, n29164, n2604, n29163, 
        n2605, n29162, n2606, n29161, n27758, n2607, n29160, n27750, 
        n2608, n29159;
    wire [31:0]n971;
    
    wire n905, n28195, n906, n28194, n27757, n2609, n43155, n29158, 
        n28193, n27749, n17101, n28192, n14346, n28191, n2489, 
        n2522, n29157, n2490, n29156, n2491, n29155, n27756, n2492, 
        n29154, n2493, n29153, n2494, n29152, n2495, n29151, n2496, 
        n29150, n2497, n29149, n1103, n4_adj_4578, n1037, n28162, 
        n1104, n1005, n28161, n1105, n1006, n28160, n2498, n29148, 
        n1106, n1007, n28159, n2499, n29147, n1107, n1008, n28158, 
        n2500, n29146, n27778, n1108, n1009, n43158, n28157, n27777, 
        n1109, n2501, n29145, n1202, n1136, n28156, n1203, n28155, 
        n1204, n28154, n2502, n29144, n27776, n2503, n29143, n1205, 
        n28153, n1206, n28152, n1207, n28151, n1208, n43159, n28150, 
        n1209, n2504, n29142, n27775, n1301, n1235, n28149, n1302, 
        n28148, n1303, n28147, n2505, n29141, n1304, n28146, n1305, 
        n28145, n1306, n28144, n2506, n29140, n2507, n29139, n1307, 
        n28143, n1308, n43160, n28142, n1309, n27748, n2508, n29138, 
        n27755, n2509, n43157, n29137, n1400, n1334, n28134, n1401, 
        n28133, n27774, n1402, n28132, n1403, n28131, n1404, n28130, 
        n1405, n28129, n1406, n28128, n27773, n1407, n28127, n1408, 
        n43161, n28126, n1409, n27754, n27772, n2390, n29136, 
        n2391, n29135, n2392, n29134, n2393, n29133, n27771, n27770, 
        n2394, n29132, n2395, n29131, n2396, n29130, n2397, n29129, 
        n2398, n29128, n1433, n28093, n28092, n28091, n2399, n29127, 
        n28090, n28089, n28088, n28087, n28086, n28085, n43163, 
        n28084, n2400, n29126, n27769, n2401, n29125, n2402, n29124, 
        n27768, n2403, n29123, n2404, n29122, n2405, n29121, n2406, 
        n29120, n2407, n29119, n27767, n29118, n29117, n2324, 
        n29116, n29115, n27766, n29114, n29113, n29112, n3182, 
        n29304, n3183, n29303, n29111, n29110, n3184, n29302, 
        n28038, n28037, n28036, n29109, n28035, n28034, n29108, 
        n29107, n29106, n3185, n29301, n28033, n28032, n3186, 
        n29300, n28031, n29105, n28030, n29104, n28029, n28028, 
        n28027, n28026, n28025, n28024, n3187, n29299, n29103, 
        n28023, n28022, n28021, n28020, n28019, n28018, n28017, 
        n28016, n29102, n29101, n28015, n29100, n28014, n3188, 
        n28013, n28012, n3189, n22_adj_4579, n15_adj_4580, n20_adj_4581, 
        n24_adj_4582, n28_adj_4583, n38_adj_4584, n24584, n36_adj_4585, 
        n42_adj_4586, n40_adj_4587, n41_adj_4588, n39, n24446, n16_adj_4589, 
        n17_adj_4590, n24_adj_4591, n22_adj_4592, n23_adj_4593, n27_adj_4594, 
        n21_adj_4595, n33_adj_4596, n32_adj_4597, n31_adj_4598, n35, 
        n37_adj_4599, n37_adj_4600, n40_adj_4601, n45_adj_4602, n38_adj_4603, 
        n39_adj_4604, n42_adj_4605, n32_adj_4606, n37_adj_4607, n34, 
        n42_adj_4608, n46_adj_4609, n33_adj_4610, n14_adj_4611, n15_adj_4612, 
        n44_adj_4613, n14_adj_4614, n9_adj_4615, n26_adj_4616, n19_adj_4617, 
        n16_adj_4618, n24_adj_4619, n28_adj_4620, n24154, n12_adj_4621, 
        n31265, n38102, n38124, n6_adj_4622, n34_adj_4623, n41_adj_4624, 
        n38_adj_4625, n43_adj_4626, n40_adj_4627, n46_adj_4628, n39_adj_4629, 
        n47_adj_4630, n18_adj_4631, n28_adj_4632, n26_adj_4633, n27_adj_4634, 
        n25_adj_4635, n24_adj_4636, n34_adj_4637, n22_adj_4638, n38_adj_4639, 
        n36_adj_4640, n37_adj_4641, n35_adj_4642, n22_adj_4643, n30_adj_4644, 
        n34_adj_4645, n32_adj_4646, n33_adj_4647, n31_adj_4648, n50_adj_4649, 
        n48_adj_4650, n60, n739, n30411, n708, n35452, n24408, 
        n35476, n103, n34609, n24462, n48_adj_4651, n46_adj_4652, 
        n47_adj_4653, n45_adj_4654, n44_adj_4655, n43_adj_4656, n54_adj_4657, 
        n49_adj_4658, n24464, n2_adj_4659, n4_adj_4660, n41190, n7_adj_4661, 
        n38086, n49_adj_4662, n1169, n13389, n36_adj_4663, n25_adj_4664, 
        n34_adj_4665, n40_adj_4666, n38_adj_4667, n39_adj_4668, n37_adj_4669, 
        n47_adj_4670;
    
    SB_CARRY mod_5_add_2143_22 (.CI(n29297), .I0(n3090), .I1(n3116), .CO(n29298));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n43140), 
            .I3(n29098), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n29098), .I0(n2309), .I1(n43140), .CO(n29099));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n29296), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n37261), .D(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n43140), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_21 (.CI(n29296), .I0(n3091), .I1(n3116), .CO(n29297));
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n43140), 
            .CO(n29098));
    SB_LUT4 add_21_19_lut (.I0(n19), .I1(bit_ctr[17]), .I2(GND_net), .I3(n27764), 
            .O(n40238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n29097), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n29295), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n29096), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n29295), .I0(n3092), .I1(n3116), .CO(n29296));
    SB_CARRY mod_5_add_1540_19 (.CI(n29096), .I0(n2193), .I1(n2225), .CO(n29097));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n28010), .O(one_wire_N_513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n29294), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n29095), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n29294), .I0(n3093), .I1(n3116), .CO(n29295));
    SB_CARRY mod_5_add_1540_18 (.CI(n29095), .I0(n2194), .I1(n2225), .CO(n29096));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n29293), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_5 (.CI(n28010), .I0(timer[3]), .I1(n1[3]), .CO(n28011));
    SB_CARRY mod_5_add_2143_18 (.CI(n29293), .I0(n3094), .I1(n3116), .CO(n29294));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n29094), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n29292), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n29094), .I0(n2195), .I1(n2225), .CO(n29095));
    SB_CARRY mod_5_add_2143_17 (.CI(n29292), .I0(n3095), .I1(n3116), .CO(n29293));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n29093), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n29291), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n29093), .I0(n2196), .I1(n2225), .CO(n29094));
    SB_CARRY mod_5_add_2143_16 (.CI(n29291), .I0(n3096), .I1(n3116), .CO(n29292));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n29092), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n29290), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n29092), .I0(n2197), .I1(n2225), .CO(n29093));
    SB_CARRY mod_5_add_2143_15 (.CI(n29290), .I0(n3097), .I1(n3116), .CO(n29291));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n29091), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n29289), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n29091), .I0(n2198), .I1(n2225), .CO(n29092));
    SB_CARRY mod_5_add_2143_14 (.CI(n29289), .I0(n3098), .I1(n3116), .CO(n29290));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n29090), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n29288), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n29090), .I0(n2199), .I1(n2225), .CO(n29091));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n28009), .O(one_wire_N_513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n29288), .I0(n3099), .I1(n3116), .CO(n29289));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n29089), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n29287), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n29089), .I0(n2200), .I1(n2225), .CO(n29090));
    SB_CARRY mod_5_add_2143_12 (.CI(n29287), .I0(n3100), .I1(n3116), .CO(n29288));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n29088), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n29286), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n29088), .I0(n2201), .I1(n2225), .CO(n29089));
    SB_CARRY sub_14_add_2_4 (.CI(n28009), .I0(timer[2]), .I1(n1[2]), .CO(n28010));
    SB_CARRY mod_5_add_2143_11 (.CI(n29286), .I0(n3101), .I1(n3116), .CO(n29287));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n29087), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n29087), .I0(n2202), .I1(n2225), .CO(n29088));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n29285), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n29086), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n33435));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n33465));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n33467));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n33469));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n33471));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n33473));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n33475));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n33477));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(VCC_net), 
            .D(n33429));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(VCC_net), 
            .D(n33431));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n33443));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n33445));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n33451));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n33453));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n33455));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n33457));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n33497));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n33493));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n33495));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n33489));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n33491));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n33485));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n33487));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n33479));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n33481));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n33483));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n33463));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n33461));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(VCC_net), 
            .D(n33433));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2143_10 (.CI(n29285), .I0(n3102), .I1(n3116), .CO(n29286));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n29284), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19788_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n24514));
    defparam i19788_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18), 
            .O(n30_adj_4539));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2098), .I1(n24514), .I2(n2094), .I3(n2099), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30_adj_4539), 
            .O(n2126));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36311_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43141));
    defparam i36311_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_9 (.CI(n29284), .I0(n3103), .I1(n3116), .CO(n29285));
    SB_CARRY mod_5_add_1540_9 (.CI(n29086), .I0(n2203), .I1(n2225), .CO(n29087));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n29085), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut (.I0(n3001), .I1(n3002), .I2(n2994), .I3(n2991), 
            .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n2989), .I1(n2990), .I2(n2996), .I3(n3007), 
            .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1585 (.I0(n3005), .I1(n3008), .I2(n2988), .I3(n2998), 
            .O(n42));
    defparam i16_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2986), .I1(n2995), .I2(n2997), .I3(n2985), 
            .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2984), .I1(n2992), .I2(n2993), .I3(n3003), 
            .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_3_lut (.I0(n3006), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n38));
    defparam i12_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i20_3_lut (.I0(n3000), .I1(n40), .I2(n2987), .I3(GND_net), 
            .O(n46));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_2_lut (.I0(n2999), .I1(n3004), .I2(GND_net), .I3(GND_net), 
            .O(n37));
    defparam i11_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n29283), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n29283), .I0(n3104), .I1(n3116), .CO(n29284));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n29282), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25_4_lut (.I0(n37), .I1(n50), .I2(n46), .I3(n38), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_7 (.CI(n29282), .I0(n3105), .I1(n3116), .CO(n29283));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4), .I1(timer[1]), .I2(n1[1]), .I3(n28008), 
            .O(n30079)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n29281), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n28008), .I0(timer[1]), .I1(n1[1]), .CO(n28009));
    SB_CARRY mod_5_add_2143_6 (.CI(n29281), .I0(n3106), .I1(n3116), .CO(n29282));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n29280), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n29280), .I0(n3107), .I1(n3116), .CO(n29281));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n29279), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n29085), .I0(n2204), .I1(n2225), .CO(n29086));
    SB_CARRY mod_5_add_2143_4 (.CI(n29279), .I0(n3108), .I1(n3116), .CO(n29280));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n43139), 
            .I3(n29278), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n29278), .I0(n3109), .I1(n43139), .CO(n29279));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n43139), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n29084), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_513[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1540_7 (.CI(n29084), .I0(n2205), .I1(n2225), .CO(n29085));
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n43139), 
            .CO(n29278));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n29277), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n29083), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n29083), .I0(n2206), .I1(n2225), .CO(n29084));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n29276), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n29082), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n29082), .I0(n2207), .I1(n2225), .CO(n29083));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n29081), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n29276), .I0(n2985), .I1(n3017), .CO(n29277));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), .I3(GND_net), 
            .O(n13));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n28008));
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4540));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1586 (.I0(n13), .I1(n20), .I2(n1605), .I3(n1599), 
            .O(n22));
    defparam i10_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1587 (.I0(n1601), .I1(n22), .I2(n18_adj_4540), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n29275), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n29081), .I0(n2208), .I1(n2225), .CO(n29082));
    SB_CARRY mod_5_add_2076_26 (.CI(n29275), .I0(n2986), .I1(n3017), .CO(n29276));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n43141), 
            .I3(n29080), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n29274), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_3 (.CI(n29080), .I0(n2209), .I1(n43141), .CO(n29081));
    SB_CARRY mod_5_add_2076_25 (.CI(n29274), .I0(n2987), .I1(n3017), .CO(n29275));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n43141), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n43141), 
            .CO(n29080));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n29273), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n29079), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n29078), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n29273), .I0(n2988), .I1(n3017), .CO(n29274));
    SB_CARRY add_21_19 (.CI(n27764), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27765));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n29272), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n29272), .I0(n2989), .I1(n3017), .CO(n29273));
    SB_CARRY mod_5_add_1473_18 (.CI(n29078), .I0(n2094), .I1(n2126), .CO(n29079));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n29271), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n29271), .I0(n2990), .I1(n3017), .CO(n29272));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n29077), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n29270), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n29077), .I0(n2095), .I1(n2126), .CO(n29078));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n29076), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n29270), .I0(n2991), .I1(n3017), .CO(n29271));
    SB_CARRY mod_5_add_1473_16 (.CI(n29076), .I0(n2096), .I1(n2126), .CO(n29077));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n29269), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n29269), .I0(n2992), .I1(n3017), .CO(n29270));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n29268), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n29268), .I0(n2993), .I1(n3017), .CO(n29269));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n29267), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n29267), .I0(n2994), .I1(n3017), .CO(n29268));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n29266), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n29266), .I0(n2995), .I1(n3017), .CO(n29267));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n29075), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n29075), .I0(n2097), .I1(n2126), .CO(n29076));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n29074), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n29265), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n29265), .I0(n2996), .I1(n3017), .CO(n29266));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n29264), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n29074), .I0(n2098), .I1(n2126), .CO(n29075));
    SB_CARRY mod_5_add_2076_15 (.CI(n29264), .I0(n2997), .I1(n3017), .CO(n29265));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n29263), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n29263), .I0(n2998), .I1(n3017), .CO(n29264));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n29262), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n29262), .I0(n2999), .I1(n3017), .CO(n29263));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n29261), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n29073), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n29073), .I0(n2099), .I1(n2126), .CO(n29074));
    SB_LUT4 i36309_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43139));
    defparam i36309_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n29072), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n29261), .I0(n3000), .I1(n3017), .CO(n29262));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n29260), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n29260), .I0(n3001), .I1(n3017), .CO(n29261));
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n29259), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36321_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43151));
    defparam i36321_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1473_12 (.CI(n29072), .I0(n2100), .I1(n2126), .CO(n29073));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n29071), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n29071), .I0(n2101), .I1(n2126), .CO(n29072));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n29070), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n29070), .I0(n2102), .I1(n2126), .CO(n29071));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n29069), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n29069), .I0(n2103), .I1(n2126), .CO(n29070));
    SB_CARRY mod_5_add_2076_10 (.CI(n29259), .I0(n3002), .I1(n3017), .CO(n29260));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n29068), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n29068), .I0(n2104), .I1(n2126), .CO(n29069));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n29067), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(n19), .I1(bit_ctr[16]), .I2(GND_net), .I3(n27763), 
            .O(n40237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1473_7 (.CI(n29067), .I0(n2105), .I1(n2126), .CO(n29068));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n29066), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4541));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1588 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46_adj_4542));
    defparam i18_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n29258), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n29258), .I0(n3003), .I1(n3017), .CO(n29259));
    SB_CARRY mod_5_add_1473_6 (.CI(n29066), .I0(n2106), .I1(n2126), .CO(n29067));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n29065), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n27752), 
            .O(n40231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n29257), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n29065), .I0(n2107), .I1(n2126), .CO(n29066));
    SB_CARRY mod_5_add_2076_8 (.CI(n29257), .I0(n3004), .I1(n3017), .CO(n29258));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n29064), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n29064), .I0(n2108), .I1(n2126), .CO(n29065));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n29256), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n29256), .I0(n3005), .I1(n3017), .CO(n29257));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n29255), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n43143), 
            .I3(n29063), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_6 (.CI(n29255), .I0(n3006), .I1(n3017), .CO(n29256));
    SB_CARRY mod_5_add_1473_3 (.CI(n29063), .I0(n2109), .I1(n43143), .CO(n29064));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n43143), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n29254), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n29254), .I0(n3007), .I1(n3017), .CO(n29255));
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n43143), 
            .CO(n29063));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n29062), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n29061), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n29253), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n29253), .I0(n3008), .I1(n3017), .CO(n29254));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n43142), 
            .I3(n29252), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_17 (.CI(n29061), .I0(n1995), .I1(n2027), .CO(n29062));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n29060), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_3 (.CI(n29252), .I0(n3009), .I1(n43142), .CO(n29253));
    SB_CARRY mod_5_add_1406_16 (.CI(n29060), .I0(n1996), .I1(n2027), .CO(n29061));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n43142), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i19_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1589 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n29059), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1590 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44_adj_4543));
    defparam i16_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1591 (.I0(bit_ctr[3]), .I1(n30_adj_4541), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43_adj_4544));
    defparam i15_4_lut_adj_1591.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46_adj_4542), .I3(n48), 
            .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43_adj_4544), .I3(n44_adj_4543), 
            .O(\state_3__N_362[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2057_3_lut (.I0(n15745), .I1(\state_3__N_362[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4414));
    defparam i2057_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n1166), .I2(n4414), .I3(\state[0] ), 
            .O(n4442));
    defparam i2_4_lut.LUT_INIT = 16'hf0ee;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n43142), 
            .CO(n29252));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n29251), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n29059), .I0(n1997), .I1(n2027), .CO(n29060));
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n29250), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n29250), .I0(n2886), .I1(n2918), .CO(n29251));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n29058), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n29249), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n29249), .I0(n2887), .I1(n2918), .CO(n29250));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n29248), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n29058), .I0(n1998), .I1(n2027), .CO(n29059));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n29057), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n29248), .I0(n2888), .I1(n2918), .CO(n29249));
    SB_CARRY mod_5_add_1406_13 (.CI(n29057), .I0(n1999), .I1(n2027), .CO(n29058));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n29247), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n29056), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n29056), .I0(n2000), .I1(n2027), .CO(n29057));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n29055), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n29247), .I0(n2889), .I1(n2918), .CO(n29248));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n29246), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n29055), .I0(n2001), .I1(n2027), .CO(n29056));
    SB_LUT4 timer_1186_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28565), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n29246), .I0(n2890), .I1(n2918), .CO(n29247));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n29054), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n29054), .I0(n2002), .I1(n2027), .CO(n29055));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n29245), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n29245), .I0(n2891), .I1(n2918), .CO(n29246));
    SB_LUT4 timer_1186_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28564), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_32 (.CI(n28564), .I0(GND_net), .I1(timer[30]), 
            .CO(n28565));
    SB_LUT4 timer_1186_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28563), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_31 (.CI(n28563), .I0(GND_net), .I1(timer[29]), 
            .CO(n28564));
    SB_LUT4 timer_1186_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28562), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_30 (.CI(n28562), .I0(GND_net), .I1(timer[28]), 
            .CO(n28563));
    SB_LUT4 timer_1186_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28561), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n29244), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1186_add_4_29 (.CI(n28561), .I0(GND_net), .I1(timer[27]), 
            .CO(n28562));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n29053), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1186_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28560), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_28 (.CI(n28560), .I0(GND_net), .I1(timer[26]), 
            .CO(n28561));
    SB_CARRY mod_5_add_2009_20 (.CI(n29244), .I0(n2892), .I1(n2918), .CO(n29245));
    SB_LUT4 timer_1186_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28559), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_27 (.CI(n28559), .I0(GND_net), .I1(timer[25]), 
            .CO(n28560));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n29243), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n29053), .I0(n2003), .I1(n2027), .CO(n29054));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n29052), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n29243), .I0(n2893), .I1(n2918), .CO(n29244));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n29242), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n29052), .I0(n2004), .I1(n2027), .CO(n29053));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n29051), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n29242), .I0(n2894), .I1(n2918), .CO(n29243));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n29241), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n29051), .I0(n2005), .I1(n2027), .CO(n29052));
    SB_CARRY mod_5_add_2009_17 (.CI(n29241), .I0(n2895), .I1(n2918), .CO(n29242));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n29050), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n29050), .I0(n2006), .I1(n2027), .CO(n29051));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n29240), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1186_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28558), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n29240), .I0(n2896), .I1(n2918), .CO(n29241));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n29239), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n29239), .I0(n2897), .I1(n2918), .CO(n29240));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n29238), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n29049), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n29049), .I0(n2007), .I1(n2027), .CO(n29050));
    SB_CARRY timer_1186_add_4_26 (.CI(n28558), .I0(GND_net), .I1(timer[24]), 
            .CO(n28559));
    SB_LUT4 timer_1186_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28557), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n29048), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n29048), .I0(n2008), .I1(n2027), .CO(n29049));
    SB_CARRY timer_1186_add_4_25 (.CI(n28557), .I0(GND_net), .I1(timer[23]), 
            .CO(n28558));
    SB_LUT4 timer_1186_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28556), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n43144), 
            .I3(n29047), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1186_add_4_24 (.CI(n28556), .I0(GND_net), .I1(timer[22]), 
            .CO(n28557));
    SB_CARRY mod_5_add_2009_14 (.CI(n29238), .I0(n2898), .I1(n2918), .CO(n29239));
    SB_LUT4 timer_1186_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28555), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_23 (.CI(n28555), .I0(GND_net), .I1(timer[21]), 
            .CO(n28556));
    SB_CARRY mod_5_add_1406_3 (.CI(n29047), .I0(n2009), .I1(n43144), .CO(n29048));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n29237), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n43144), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_13 (.CI(n29237), .I0(n2899), .I1(n2918), .CO(n29238));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n29236), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1186_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28554), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n29236), .I0(n2900), .I1(n2918), .CO(n29237));
    SB_CARRY timer_1186_add_4_22 (.CI(n28554), .I0(GND_net), .I1(timer[20]), 
            .CO(n28555));
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n43144), 
            .CO(n29047));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n29046), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1186_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28553), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n29045), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1186_add_4_21 (.CI(n28553), .I0(GND_net), .I1(timer[19]), 
            .CO(n28554));
    SB_LUT4 timer_1186_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28552), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_20 (.CI(n28552), .I0(GND_net), .I1(timer[18]), 
            .CO(n28553));
    SB_LUT4 timer_1186_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28551), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_19 (.CI(n28551), .I0(GND_net), .I1(timer[17]), 
            .CO(n28552));
    SB_LUT4 timer_1186_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28550), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_18 (.CI(n28550), .I0(GND_net), .I1(timer[16]), 
            .CO(n28551));
    SB_LUT4 timer_1186_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28549), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_17 (.CI(n28549), .I0(GND_net), .I1(timer[15]), 
            .CO(n28550));
    SB_LUT4 timer_1186_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28548), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_16 (.CI(n28548), .I0(GND_net), .I1(timer[14]), 
            .CO(n28549));
    SB_CARRY add_21_18 (.CI(n27763), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27764));
    SB_LUT4 timer_1186_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28547), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_15 (.CI(n28547), .I0(GND_net), .I1(timer[13]), 
            .CO(n28548));
    SB_LUT4 timer_1186_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28546), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_14 (.CI(n28546), .I0(GND_net), .I1(timer[12]), 
            .CO(n28547));
    SB_LUT4 timer_1186_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28545), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_13 (.CI(n28545), .I0(GND_net), .I1(timer[11]), 
            .CO(n28546));
    SB_LUT4 timer_1186_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28544), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_12 (.CI(n28544), .I0(GND_net), .I1(timer[10]), 
            .CO(n28545));
    SB_LUT4 timer_1186_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28543), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_11 (.CI(n28543), .I0(GND_net), .I1(timer[9]), 
            .CO(n28544));
    SB_LUT4 timer_1186_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28542), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_10 (.CI(n28542), .I0(GND_net), .I1(timer[8]), 
            .CO(n28543));
    SB_LUT4 add_21_17_lut (.I0(n19), .I1(bit_ctr[15]), .I2(GND_net), .I3(n27762), 
            .O(n40236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1186_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28541), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_9 (.CI(n28541), .I0(GND_net), .I1(timer[7]), 
            .CO(n28542));
    SB_LUT4 timer_1186_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28540), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n29235), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n29045), .I0(n1896), .I1(n1928), .CO(n29046));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n29044), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1186_add_4_8 (.CI(n28540), .I0(GND_net), .I1(timer[6]), 
            .CO(n28541));
    SB_LUT4 timer_1186_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28539), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_7 (.CI(n28539), .I0(GND_net), .I1(timer[5]), 
            .CO(n28540));
    SB_LUT4 timer_1186_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28538), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_6 (.CI(n28538), .I0(GND_net), .I1(timer[4]), 
            .CO(n28539));
    SB_CARRY mod_5_add_1339_15 (.CI(n29044), .I0(n1897), .I1(n1928), .CO(n29045));
    SB_CARRY mod_5_add_2009_11 (.CI(n29235), .I0(n2901), .I1(n2918), .CO(n29236));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n29043), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n29043), .I0(n1898), .I1(n1928), .CO(n29044));
    SB_LUT4 timer_1186_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28537), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n29042), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n29042), .I0(n1899), .I1(n1928), .CO(n29043));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n29234), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n29041), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1186_add_4_5 (.CI(n28537), .I0(GND_net), .I1(timer[3]), 
            .CO(n28538));
    SB_LUT4 timer_1186_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28536), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_4 (.CI(n28536), .I0(GND_net), .I1(timer[2]), 
            .CO(n28537));
    SB_LUT4 timer_1186_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28535), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1186_add_4_3 (.CI(n28535), .I0(GND_net), .I1(timer[1]), 
            .CO(n28536));
    SB_LUT4 timer_1186_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1186_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n29041), .I0(n1900), .I1(n1928), .CO(n29042));
    SB_CARRY timer_1186_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28535));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n29040), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n29234), .I0(n2902), .I1(n2918), .CO(n29235));
    SB_CARRY mod_5_add_1339_11 (.CI(n29040), .I0(n1901), .I1(n1928), .CO(n29041));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n29039), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n29233), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n29039), .I0(n1902), .I1(n1928), .CO(n29040));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n29038), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n29038), .I0(n1903), .I1(n1928), .CO(n29039));
    SB_CARRY mod_5_add_2009_9 (.CI(n29233), .I0(n2903), .I1(n2918), .CO(n29234));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n29037), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n29037), .I0(n1904), .I1(n1928), .CO(n29038));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n29232), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n29036), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n29232), .I0(n2904), .I1(n2918), .CO(n29233));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n29231), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n29231), .I0(n2905), .I1(n2918), .CO(n29232));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n29230), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n29036), .I0(n1905), .I1(n1928), .CO(n29037));
    SB_CARRY mod_5_add_2009_6 (.CI(n29230), .I0(n2906), .I1(n2918), .CO(n29231));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n29229), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n29229), .I0(n2907), .I1(n2918), .CO(n29230));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n29035), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n29035), .I0(n1906), .I1(n1928), .CO(n29036));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n29228), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n29034), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n29228), .I0(n2908), .I1(n2918), .CO(n29229));
    SB_CARRY mod_5_add_1339_5 (.CI(n29034), .I0(n1907), .I1(n1928), .CO(n29035));
    SB_CARRY add_21_7 (.CI(n27752), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27753));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n43145), 
            .I3(n29227), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n29033), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_3 (.CI(n29227), .I0(n2909), .I1(n43145), .CO(n29228));
    SB_CARRY add_21_17 (.CI(n27762), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27763));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n43145), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n43145), 
            .CO(n29227));
    SB_CARRY mod_5_add_1339_4 (.CI(n29033), .I0(n1908), .I1(n1928), .CO(n29034));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n43146), 
            .I3(n29032), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n29226), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n29225), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n29225), .I0(n2787), .I1(n2819), .CO(n29226));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n29224), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_3 (.CI(n29032), .I0(n1909), .I1(n43146), .CO(n29033));
    SB_CARRY mod_5_add_1942_24 (.CI(n29224), .I0(n2788), .I1(n2819), .CO(n29225));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n43146), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n43146), 
            .CO(n29032));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n29031), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n29030), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n29030), .I0(n1797), .I1(n1829), .CO(n29031));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n29029), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n27751), 
            .O(n40245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n27761), 
            .O(n40234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n29223), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n29223), .I0(n2789), .I1(n2819), .CO(n29224));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n29222), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n29222), .I0(n2790), .I1(n2819), .CO(n29223));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n29221), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n29029), .I0(n1798), .I1(n1829), .CO(n29030));
    SB_CARRY mod_5_add_1942_21 (.CI(n29221), .I0(n2791), .I1(n2819), .CO(n29222));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n29220), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n29220), .I0(n2792), .I1(n2819), .CO(n29221));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n29028), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n29219), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n29219), .I0(n2793), .I1(n2819), .CO(n29220));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n29218), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n29028), .I0(n1799), .I1(n1829), .CO(n29029));
    SB_CARRY mod_5_add_1942_18 (.CI(n29218), .I0(n2794), .I1(n2819), .CO(n29219));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n29217), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n29217), .I0(n2795), .I1(n2819), .CO(n29218));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n29027), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n29216), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n29027), .I0(n1800), .I1(n1829), .CO(n29028));
    SB_CARRY mod_5_add_1942_16 (.CI(n29216), .I0(n2796), .I1(n2819), .CO(n29217));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n29215), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n29215), .I0(n2797), .I1(n2819), .CO(n29216));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n29214), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n29214), .I0(n2798), .I1(n2819), .CO(n29215));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n29026), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n29213), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n29213), .I0(n2799), .I1(n2819), .CO(n29214));
    SB_CARRY mod_5_add_1272_11 (.CI(n29026), .I0(n1801), .I1(n1829), .CO(n29027));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n29212), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n29212), .I0(n2800), .I1(n2819), .CO(n29213));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n29211), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n29025), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n29025), .I0(n1802), .I1(n1829), .CO(n29026));
    SB_CARRY mod_5_add_1942_11 (.CI(n29211), .I0(n2801), .I1(n2819), .CO(n29212));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n29024), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n29210), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n29024), .I0(n1803), .I1(n1829), .CO(n29025));
    SB_CARRY mod_5_add_1942_10 (.CI(n29210), .I0(n2802), .I1(n2819), .CO(n29211));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n29209), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n29023), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n29209), .I0(n2803), .I1(n2819), .CO(n29210));
    SB_CARRY mod_5_add_1272_8 (.CI(n29023), .I0(n1804), .I1(n1829), .CO(n29024));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n29022), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n29208), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n29022), .I0(n1805), .I1(n1829), .CO(n29023));
    SB_CARRY mod_5_add_1942_8 (.CI(n29208), .I0(n2804), .I1(n2819), .CO(n29209));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n29207), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n29021), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n29207), .I0(n2805), .I1(n2819), .CO(n29208));
    SB_CARRY mod_5_add_1272_6 (.CI(n29021), .I0(n1806), .I1(n1829), .CO(n29022));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n29206), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n29020), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n29206), .I0(n2806), .I1(n2819), .CO(n29207));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n29205), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n29020), .I0(n1807), .I1(n1829), .CO(n29021));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n29019), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n29019), .I0(n1808), .I1(n1829), .CO(n29020));
    SB_CARRY mod_5_add_1942_5 (.CI(n29205), .I0(n2807), .I1(n2819), .CO(n29206));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n29204), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n29204), .I0(n2808), .I1(n2819), .CO(n29205));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n43148), 
            .I3(n29203), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n29203), .I0(n2809), .I1(n43148), .CO(n29204));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n43148), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n43148), 
            .CO(n29203));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n29202), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n29201), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n29201), .I0(n2688), .I1(n2720), .CO(n29202));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n29200), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n43149), 
            .I3(n29018), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_23 (.CI(n29200), .I0(n2689), .I1(n2720), .CO(n29201));
    SB_CARRY mod_5_add_1272_3 (.CI(n29018), .I0(n1809), .I1(n43149), .CO(n29019));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n29199), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n43149), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_22 (.CI(n29199), .I0(n2690), .I1(n2720), .CO(n29200));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n29198), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n29198), .I0(n2691), .I1(n2720), .CO(n29199));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n29197), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n29197), .I0(n2692), .I1(n2720), .CO(n29198));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n29196), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1186__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n43149), 
            .CO(n29018));
    SB_CARRY mod_5_add_1875_19 (.CI(n29196), .I0(n2693), .I1(n2720), .CO(n29197));
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n29017), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n29195), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n29016), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_16 (.CI(n27761), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27762));
    SB_CARRY mod_5_add_1875_18 (.CI(n29195), .I0(n2694), .I1(n2720), .CO(n29196));
    SB_CARRY mod_5_add_1205_14 (.CI(n29016), .I0(n1698), .I1(n1730), .CO(n29017));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n29194), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n29194), .I0(n2695), .I1(n2720), .CO(n29195));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n29193), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n29193), .I0(n2696), .I1(n2720), .CO(n29194));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n29192), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n29015), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n29015), .I0(n1699), .I1(n1730), .CO(n29016));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n29014), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n29014), .I0(n1700), .I1(n1730), .CO(n29015));
    SB_CARRY mod_5_add_1875_15 (.CI(n29192), .I0(n2697), .I1(n2720), .CO(n29193));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n29191), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n29013), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n29191), .I0(n2698), .I1(n2720), .CO(n29192));
    SB_CARRY mod_5_add_1205_11 (.CI(n29013), .I0(n1701), .I1(n1730), .CO(n29014));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n29012), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n29190), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n29012), .I0(n1702), .I1(n1730), .CO(n29013));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n29011), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n29011), .I0(n1703), .I1(n1730), .CO(n29012));
    SB_CARRY mod_5_add_1875_13 (.CI(n29190), .I0(n2699), .I1(n2720), .CO(n29191));
    SB_LUT4 i10_4_lut_adj_1592 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4545));
    defparam i10_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1593 (.I0(n2203), .I1(n28_adj_4545), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4546));
    defparam i14_4_lut_adj_1593.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1594 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4547));
    defparam i12_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1595 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4548));
    defparam i13_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1596 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4549));
    defparam i11_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1597 (.I0(n29_adj_4549), .I1(n31_adj_4548), .I2(n30_adj_4547), 
            .I3(n32_adj_4546), .O(n2225));
    defparam i17_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[4]), .I2(one_wire_N_513[2]), 
            .I3(GND_net), .O(n29824));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i19901_2_lut (.I0(n29824), .I1(n15631), .I2(GND_net), .I3(GND_net), 
            .O(n24628));
    defparam i19901_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1598 (.I0(n24324), .I1(one_wire_N_513[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4550));
    defparam i1_2_lut_adj_1598.LUT_INIT = 16'heeee;
    SB_LUT4 equal_335_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n15744));
    defparam equal_335_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut_adj_1599 (.I0(\one_wire_N_513[10] ), .I1(\one_wire_N_513[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/neopixel.v(62[15:42])
    defparam i2_2_lut_adj_1599.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(\one_wire_N_513[5] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[7] ), .I3(n15824), .O(n14));   // verilog/neopixel.v(62[15:42])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(\one_wire_N_513[9] ), .I1(n14), .I2(n10), .I3(\one_wire_N_513[6] ), 
            .O(n15631));   // verilog/neopixel.v(62[15:42])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28566_2_lut (.I0(\state[1] ), .I1(n15745), .I2(GND_net), 
            .I3(GND_net), .O(n35327));
    defparam i28566_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n29010), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n33459));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i7_4_lut_adj_1600 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4551));
    defparam i7_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1504), .I1(n18_adj_4551), .I2(n1502), .I3(n1499), 
            .O(n20_adj_4552));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), .I3(GND_net), 
            .O(n15));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1601 (.I0(n15), .I1(n20_adj_4552), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n33441));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n33439));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17493));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17492));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17491));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17490));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17489));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17488));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17487));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17486));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17485));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17484));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17483));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17482));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17481));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17480));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17479));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17478));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17477));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17476));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17475));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17474));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17473));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17472));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17471));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17470));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17469));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17468));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17467));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17466));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17465));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17464));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17463));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n27880), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1602 (.I0(n21), .I1(n23), .I2(n22_adj_4553), 
            .I3(n24), .O(n36));   // verilog/neopixel.v(62[15:42])
    defparam i16_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1603 (.I0(n25), .I1(n27_adj_4554), .I2(n26), 
            .I3(n28_adj_4555), .O(n37_adj_4556));   // verilog/neopixel.v(62[15:42])
    defparam i17_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1604 (.I0(n37_adj_4556), .I1(n29_adj_4557), .I2(n36), 
            .I3(n30_adj_4558), .O(n15824));   // verilog/neopixel.v(62[15:42])
    defparam i19_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1605 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34689));
    defparam i1_2_lut_adj_1605.LUT_INIT = 16'h2222;
    SB_LUT4 i28609_2_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[2]), 
            .I2(GND_net), .I3(GND_net), .O(n35373));
    defparam i28609_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19598_2_lut (.I0(n30079), .I1(one_wire_N_513[3]), .I2(GND_net), 
            .I3(GND_net), .O(n24324));
    defparam i19598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1606 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_1606.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_513[4]), .I1(n34738), .I2(n24324), 
            .I3(n35373), .O(n116));
    defparam i1_4_lut.LUT_INIT = 16'h45cd;
    SB_LUT4 i36287_3_lut (.I0(n35462), .I1(n116), .I2(n15824), .I3(GND_net), 
            .O(n37261));
    defparam i36287_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY mod_5_add_1205_8 (.CI(n29010), .I0(n1704), .I1(n1730), .CO(n29011));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n29009), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n29189), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n29009), .I0(n1705), .I1(n1730), .CO(n29010));
    SB_CARRY mod_5_add_1875_12 (.CI(n29189), .I0(n2700), .I1(n2720), .CO(n29190));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n29008), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n29188), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n29008), .I0(n1706), .I1(n1730), .CO(n29009));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n27879), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n29188), .I0(n2701), .I1(n2720), .CO(n29189));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n29007), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n27879), .I0(n1500), .I1(n1532), .CO(n27880));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n27878), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n27878), .I0(n1501), .I1(n1532), .CO(n27879));
    SB_CARRY mod_5_add_1205_5 (.CI(n29007), .I0(n1707), .I1(n1730), .CO(n29008));
    SB_CARRY add_21_6 (.CI(n27751), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27752));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n27877), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n29187), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n29006), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n29187), .I0(n2702), .I1(n2720), .CO(n29188));
    SB_CARRY mod_5_add_1205_4 (.CI(n29006), .I0(n1708), .I1(n1730), .CO(n29007));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n43151), 
            .I3(n29005), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n29186), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_3 (.CI(n29005), .I0(n1709), .I1(n43151), .CO(n29006));
    SB_CARRY mod_5_add_1071_10 (.CI(n27877), .I0(n1502), .I1(n1532), .CO(n27878));
    SB_CARRY mod_5_add_1875_9 (.CI(n29186), .I0(n2703), .I1(n2720), .CO(n29187));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n43151), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n27876), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n29185), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n43151), 
            .CO(n29005));
    SB_CARRY mod_5_add_1071_9 (.CI(n27876), .I0(n1503), .I1(n1532), .CO(n27877));
    SB_CARRY mod_5_add_1875_8 (.CI(n29185), .I0(n2704), .I1(n2720), .CO(n29186));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n29004), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n29184), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n29003), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n29184), .I0(n2705), .I1(n2720), .CO(n29185));
    SB_CARRY mod_5_add_1138_13 (.CI(n29003), .I0(n1599), .I1(n1631), .CO(n29004));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n27875), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n29183), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n29002), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n29183), .I0(n2706), .I1(n2720), .CO(n29184));
    SB_CARRY mod_5_add_1138_12 (.CI(n29002), .I0(n1600), .I1(n1631), .CO(n29003));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n29182), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n29001), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n27760), 
            .O(n40230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_5 (.CI(n29182), .I0(n2707), .I1(n2720), .CO(n29183));
    SB_CARRY mod_5_add_1138_11 (.CI(n29001), .I0(n1601), .I1(n1631), .CO(n29002));
    SB_CARRY mod_5_add_1071_8 (.CI(n27875), .I0(n1504), .I1(n1532), .CO(n27876));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n29181), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n29000), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n27874), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n29181), .I0(n2708), .I1(n2720), .CO(n29182));
    SB_CARRY mod_5_add_1138_10 (.CI(n29000), .I0(n1602), .I1(n1631), .CO(n29001));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n43150), 
            .I3(n29180), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n28999), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_3 (.CI(n29180), .I0(n2709), .I1(n43150), .CO(n29181));
    SB_CARRY mod_5_add_1138_9 (.CI(n28999), .I0(n1603), .I1(n1631), .CO(n29000));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n43150), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n28998), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n27874), .I0(n1505), .I1(n1532), .CO(n27875));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n27873), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n43150), 
            .CO(n29180));
    SB_CARRY mod_5_add_1138_8 (.CI(n28998), .I0(n1604), .I1(n1631), .CO(n28999));
    SB_CARRY mod_5_add_1071_6 (.CI(n27873), .I0(n1506), .I1(n1532), .CO(n27874));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n29179), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n28997), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n27872), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n29178), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n28997), .I0(n1605), .I1(n1631), .CO(n28998));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n28996), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n27872), .I0(n1507), .I1(n1532), .CO(n27873));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n27871), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_15 (.CI(n27760), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27761));
    SB_CARRY mod_5_add_1808_23 (.CI(n29178), .I0(n2589), .I1(n2621), .CO(n29179));
    SB_CARRY mod_5_add_1138_6 (.CI(n28996), .I0(n1606), .I1(n1631), .CO(n28997));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n28995), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n27871), .I0(n1508), .I1(n1532), .CO(n27872));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n29177), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n28995), .I0(n1607), .I1(n1631), .CO(n28996));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n43153), 
            .I3(n27870), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_22 (.CI(n29177), .I0(n2590), .I1(n2621), .CO(n29178));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n28994), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28658_4_lut (.I0(n15631), .I1(n29824), .I2(n4_adj_4550), 
            .I3(\state[0] ), .O(n35424));
    defparam i28658_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n29176), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_4_lut (.I0(n5), .I1(\state[1] ), .I2(n15631), .I3(n35335), 
            .O(n36000));
    defparam i3_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut_adj_1607 (.I0(\state[1] ), .I1(n36000), .I2(start), 
            .I3(n35991), .O(n36115));
    defparam i2_4_lut_adj_1607.LUT_INIT = 16'h8c00;
    SB_CARRY mod_5_add_1808_21 (.CI(n29176), .I0(n2591), .I1(n2621), .CO(n29177));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17431));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_3 (.CI(n27870), .I0(n1509), .I1(n43153), .CO(n27871));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n29175), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n29175), .I0(n2592), .I1(n2621), .CO(n29176));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n29174), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n28994), .I0(n1608), .I1(n1631), .CO(n28995));
    SB_CARRY mod_5_add_1808_19 (.CI(n29174), .I0(n2593), .I1(n2621), .CO(n29175));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n43154), 
            .I3(n28993), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n28993), .I0(n1609), .I1(n43154), .CO(n28994));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n43153), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n29173), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n29173), .I0(n2594), .I1(n2621), .CO(n29174));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n43154), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n43154), 
            .CO(n28993));
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n43153), 
            .CO(n27870));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n29172), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n27759), 
            .O(n40228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_17 (.CI(n29172), .I0(n2595), .I1(n2621), .CO(n29173));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n29171), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n29171), .I0(n2596), .I1(n2621), .CO(n29172));
    SB_CARRY add_21_14 (.CI(n27759), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27760));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n29170), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n29170), .I0(n2597), .I1(n2621), .CO(n29171));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n29169), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n29169), .I0(n2598), .I1(n2621), .CO(n29170));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n29168), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17008), .D(state_3__N_362[0]), 
            .S(n35420));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n16961), .D(\neo_pixel_transmitter.done_N_576 ), 
            .R(n36877));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1808_13 (.CI(n29168), .I0(n2599), .I1(n2621), .CO(n29169));
    SB_LUT4 i3_4_lut_4_lut (.I0(n35303), .I1(n14348), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14348), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n35303), .O(n35416));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28552_2_lut_4_lut (.I0(bit_ctr[28]), .I1(bit_ctr[29]), .I2(bit_ctr[30]), 
            .I3(bit_ctr[31]), .O(n35313));
    defparam i28552_2_lut_4_lut.LUT_INIT = 16'h8208;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n29167), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n29167), .I0(n2600), .I1(n2621), .CO(n29168));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n29166), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36332_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43162));
    defparam i36332_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_11 (.CI(n29166), .I0(n2601), .I1(n2621), .CO(n29167));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n29165), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n29165), .I0(n2602), .I1(n2621), .CO(n29166));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n29164), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n29164), .I0(n2603), .I1(n2621), .CO(n29165));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n29163), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n29163), .I0(n2604), .I1(n2621), .CO(n29164));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n29162), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n29162), .I0(n2605), .I1(n2621), .CO(n29163));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n29161), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n29161), .I0(n2606), .I1(n2621), .CO(n29162));
    SB_LUT4 add_21_13_lut (.I0(n11), .I1(bit_ctr[11]), .I2(GND_net), .I3(n27758), 
            .O(n40227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n29160), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n27750), 
            .O(n40244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_13 (.CI(n27758), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27759));
    SB_DFF timer_1186__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1186__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n33499));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17248));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_5 (.CI(n27750), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27751));
    SB_CARRY mod_5_add_1808_5 (.CI(n29160), .I0(n2607), .I1(n2621), .CO(n29161));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n29159), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n28195), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28194), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_12_lut (.I0(n11), .I1(bit_ctr[10]), .I2(GND_net), .I3(n27757), 
            .O(n40223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_669_6 (.CI(n28194), .I0(n906), .I1(VCC_net), .CO(n28195));
    SB_CARRY mod_5_add_1808_4 (.CI(n29159), .I0(n2608), .I1(n2621), .CO(n29160));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n43155), 
            .I3(n29158), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n35416), .I2(VCC_net), 
            .I3(n28193), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_3 (.CI(n29158), .I0(n2609), .I1(n43155), .CO(n29159));
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n27749), 
            .O(n40235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n43155), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_669_5 (.CI(n28193), .I0(n35416), .I1(VCC_net), 
            .CO(n28194));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17101), .I2(VCC_net), 
            .I3(n28192), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n28192), .I0(n17101), .I1(VCC_net), 
            .CO(n28193));
    SB_CARRY add_21_12 (.CI(n27757), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27758));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n43155), 
            .CO(n29158));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14346), .I2(GND_net), 
            .I3(n28191), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n29157), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_3 (.CI(n28191), .I0(n14346), .I1(GND_net), 
            .CO(n28192));
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n29156), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n29156), .I0(n2490), .I1(n2522), .CO(n29157));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n27749), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27750));
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28191));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n29155), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(n11), .I1(bit_ctr[9]), .I2(GND_net), .I3(n27756), 
            .O(n40224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_21 (.CI(n29155), .I0(n2491), .I1(n2522), .CO(n29156));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n29154), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n29154), .I0(n2492), .I1(n2522), .CO(n29155));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n29153), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n29153), .I0(n2493), .I1(n2522), .CO(n29154));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n29152), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n29152), .I0(n2494), .I1(n2522), .CO(n29153));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n29151), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n29151), .I0(n2495), .I1(n2522), .CO(n29152));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n29150), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n29150), .I0(n2496), .I1(n2522), .CO(n29151));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n29149), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n29149), .I0(n2497), .I1(n2522), .CO(n29150));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4578), .I1(n4_adj_4578), .I2(n1037), 
            .I3(n28162), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28161), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28161), .I0(n1005), .I1(n1037), .CO(n28162));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28160), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n28160), .I0(n1006), .I1(n1037), .CO(n28161));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n29148), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28159), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28159), .I0(n1007), .I1(n1037), .CO(n28160));
    SB_CARRY mod_5_add_1741_14 (.CI(n29148), .I0(n2498), .I1(n2522), .CO(n29149));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n29147), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n29147), .I0(n2499), .I1(n2522), .CO(n29148));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28158), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n29146), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n27778), 
            .O(n40254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_736_4 (.CI(n28158), .I0(n1008), .I1(n1037), .CO(n28159));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n43158), 
            .I3(n28157), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n27777), 
            .O(n40253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_736_3 (.CI(n28157), .I0(n1009), .I1(n43158), .CO(n28158));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n43158), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_32 (.CI(n27777), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27778));
    SB_CARRY mod_5_add_1741_12 (.CI(n29146), .I0(n2500), .I1(n2522), .CO(n29147));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n29145), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n43158), 
            .CO(n28157));
    SB_CARRY mod_5_add_1741_11 (.CI(n29145), .I0(n2501), .I1(n2522), .CO(n29146));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28156), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28155), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28155), .I0(n1104), .I1(n1136), .CO(n28156));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28154), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n27756), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27757));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n29144), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n29144), .I0(n2502), .I1(n2522), .CO(n29145));
    SB_LUT4 add_21_31_lut (.I0(n19), .I1(bit_ctr[29]), .I2(GND_net), .I3(n27776), 
            .O(n40252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_803_7 (.CI(n28154), .I0(n1105), .I1(n1136), .CO(n28155));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n29143), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28153), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28153), .I0(n1106), .I1(n1136), .CO(n28154));
    SB_CARRY mod_5_add_1741_9 (.CI(n29143), .I0(n2503), .I1(n2522), .CO(n29144));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28152), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28152), .I0(n1107), .I1(n1136), .CO(n28153));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28151), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28151), .I0(n1108), .I1(n1136), .CO(n28152));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n43159), 
            .I3(n28150), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_31 (.CI(n27776), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27777));
    SB_CARRY mod_5_add_803_3 (.CI(n28150), .I0(n1109), .I1(n43159), .CO(n28151));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n43159), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n43159), 
            .CO(n28150));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n29142), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(n19), .I1(bit_ctr[28]), .I2(GND_net), .I3(n27775), 
            .O(n40251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28149), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28148), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28148), .I0(n1203), .I1(n1235), .CO(n28149));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28147), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n29142), .I0(n2504), .I1(n2522), .CO(n29143));
    SB_CARRY mod_5_add_870_8 (.CI(n28147), .I0(n1204), .I1(n1235), .CO(n28148));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n29141), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28146), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28146), .I0(n1205), .I1(n1235), .CO(n28147));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28145), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28145), .I0(n1206), .I1(n1235), .CO(n28146));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28144), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n29141), .I0(n2505), .I1(n2522), .CO(n29142));
    SB_CARRY mod_5_add_870_5 (.CI(n28144), .I0(n1207), .I1(n1235), .CO(n28145));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n29140), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n29140), .I0(n2506), .I1(n2522), .CO(n29141));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n29139), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28143), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n28143), .I0(n1208), .I1(n1235), .CO(n28144));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n43160), 
            .I3(n28142), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n28142), .I0(n1209), .I1(n43160), .CO(n28143));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n43160), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_5 (.CI(n29139), .I0(n2507), .I1(n2522), .CO(n29140));
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n43160), 
            .CO(n28142));
    SB_CARRY add_21_30 (.CI(n27775), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27776));
    SB_LUT4 add_21_3_lut (.I0(n11), .I1(bit_ctr[1]), .I2(GND_net), .I3(n27748), 
            .O(n40226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n29138), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(n11), .I1(bit_ctr[8]), .I2(GND_net), .I3(n27755), 
            .O(n40225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_4 (.CI(n29138), .I0(n2508), .I1(n2522), .CO(n29139));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n43157), 
            .I3(n29137), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28134), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28133), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28133), .I0(n1302), .I1(n1334), .CO(n28134));
    SB_LUT4 add_21_29_lut (.I0(n19), .I1(bit_ctr[27]), .I2(GND_net), .I3(n27774), 
            .O(n40250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28132), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28132), .I0(n1303), .I1(n1334), .CO(n28133));
    SB_CARRY add_21_29 (.CI(n27774), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27775));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28131), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n28131), .I0(n1304), .I1(n1334), .CO(n28132));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28130), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_3 (.CI(n29137), .I0(n2509), .I1(n43157), .CO(n29138));
    SB_CARRY mod_5_add_937_7 (.CI(n28130), .I0(n1305), .I1(n1334), .CO(n28131));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28129), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28129), .I0(n1306), .I1(n1334), .CO(n28130));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28128), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28128), .I0(n1307), .I1(n1334), .CO(n28129));
    SB_LUT4 add_21_28_lut (.I0(n19), .I1(bit_ctr[26]), .I2(GND_net), .I3(n27773), 
            .O(n40249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28127), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n43157), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_4 (.CI(n28127), .I0(n1308), .I1(n1334), .CO(n28128));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n43161), 
            .I3(n28126), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n28126), .I0(n1309), .I1(n43161), .CO(n28127));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n43161), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n43157), 
            .CO(n29137));
    SB_CARRY add_21_10 (.CI(n27755), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27756));
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n27754), 
            .O(n40233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_28 (.CI(n27773), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27774));
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n43161), 
            .CO(n28126));
    SB_LUT4 add_21_27_lut (.I0(n19), .I1(bit_ctr[25]), .I2(GND_net), .I3(n27772), 
            .O(n40248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n29136), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n29135), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n29135), .I0(n2391), .I1(n2423), .CO(n29136));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n29134), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n27748), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27749));
    SB_CARRY add_21_9 (.CI(n27754), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27755));
    SB_CARRY mod_5_add_1674_20 (.CI(n29134), .I0(n2392), .I1(n2423), .CO(n29135));
    SB_CARRY add_21_27 (.CI(n27772), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27773));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n29133), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_26_lut (.I0(n19), .I1(bit_ctr[24]), .I2(GND_net), .I3(n27771), 
            .O(n40247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_26 (.CI(n27771), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27772));
    SB_LUT4 add_21_25_lut (.I0(n19), .I1(bit_ctr[23]), .I2(GND_net), .I3(n27770), 
            .O(n40246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_19 (.CI(n29133), .I0(n2393), .I1(n2423), .CO(n29134));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n29132), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n29132), .I0(n2394), .I1(n2423), .CO(n29133));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n29131), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n29131), .I0(n2395), .I1(n2423), .CO(n29132));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n29130), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n29130), .I0(n2396), .I1(n2423), .CO(n29131));
    SB_CARRY add_21_25 (.CI(n27770), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27771));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n29129), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n29129), .I0(n2397), .I1(n2423), .CO(n29130));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n29128), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n29128), .I0(n2398), .I1(n2423), .CO(n29129));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28093), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28092), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28092), .I0(n1401), .I1(n1433), .CO(n28093));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28091), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n29127), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n28091), .I0(n1402), .I1(n1433), .CO(n28092));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28090), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n28090), .I0(n1403), .I1(n1433), .CO(n28091));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28089), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n28089), .I0(n1404), .I1(n1433), .CO(n28090));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28088), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n28088), .I0(n1405), .I1(n1433), .CO(n28089));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28087), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28087), .I0(n1406), .I1(n1433), .CO(n28088));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28086), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n29127), .I0(n2399), .I1(n2423), .CO(n29128));
    SB_CARRY mod_5_add_1004_5 (.CI(n28086), .I0(n1407), .I1(n1433), .CO(n28087));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28085), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28085), .I0(n1408), .I1(n1433), .CO(n28086));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n43163), 
            .I3(n28084), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n29126), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n29126), .I0(n2400), .I1(n2423), .CO(n29127));
    SB_CARRY mod_5_add_1004_3 (.CI(n28084), .I0(n1409), .I1(n43163), .CO(n28085));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n43163), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n43163), 
            .CO(n28084));
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n27769), 
            .O(n40243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n29125), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n29125), .I0(n2401), .I1(n2423), .CO(n29126));
    SB_CARRY add_21_24 (.CI(n27769), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27770));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n29124), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n40229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n27753), 
            .O(n40232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_23_lut (.I0(n19), .I1(bit_ctr[21]), .I2(GND_net), .I3(n27768), 
            .O(n40242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_10 (.CI(n29124), .I0(n2402), .I1(n2423), .CO(n29125));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n29123), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n29123), .I0(n2403), .I1(n2423), .CO(n29124));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n29122), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n29122), .I0(n2404), .I1(n2423), .CO(n29123));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n29121), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n29121), .I0(n2405), .I1(n2423), .CO(n29122));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n29120), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n29120), .I0(n2406), .I1(n2423), .CO(n29121));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n29119), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n29119), .I0(n2407), .I1(n2423), .CO(n29120));
    SB_CARRY add_21_23 (.CI(n27768), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27769));
    SB_LUT4 add_21_22_lut (.I0(n19), .I1(bit_ctr[20]), .I2(GND_net), .I3(n27767), 
            .O(n40241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n29118), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n29118), .I0(n2408), .I1(n2423), .CO(n29119));
    SB_CARRY add_21_22 (.CI(n27767), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27768));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n43162), 
            .I3(n29117), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n29117), .I0(n2409), .I1(n43162), .CO(n29118));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n43162), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n43162), 
            .CO(n29117));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n29116), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n29115), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(n19), .I1(bit_ctr[19]), .I2(GND_net), .I3(n27766), 
            .O(n40240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_21 (.CI(n27766), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27767));
    SB_CARRY mod_5_add_1607_20 (.CI(n29115), .I0(n2292), .I1(n2324), .CO(n29116));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n29114), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n29114), .I0(n2293), .I1(n2324), .CO(n29115));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n29113), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n29113), .I0(n2294), .I1(n2324), .CO(n29114));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n29112), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n29112), .I0(n2295), .I1(n2324), .CO(n29113));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n29304), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n29303), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n29111), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n29303), .I0(n3084), .I1(n3116), .CO(n29304));
    SB_CARRY mod_5_add_1607_16 (.CI(n29111), .I0(n2296), .I1(n2324), .CO(n29112));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n29110), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n29302), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n29110), .I0(n2297), .I1(n2324), .CO(n29111));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_513[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n28038), .O(n22_adj_4553)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_513[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n28037), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n28037), .I0(timer[30]), .I1(n1[30]), 
            .CO(n28038));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_513[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n28036), .O(n28_adj_4555)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n28036), .I0(timer[29]), .I1(n1[29]), 
            .CO(n28037));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n29109), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_513[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n28035), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n28035), .I0(timer[28]), .I1(n1[28]), 
            .CO(n28036));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_513[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n28034), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2143_27 (.CI(n29302), .I0(n3085), .I1(n3116), .CO(n29303));
    SB_CARRY mod_5_add_1607_14 (.CI(n29109), .I0(n2298), .I1(n2324), .CO(n29110));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n29108), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n29108), .I0(n2299), .I1(n2324), .CO(n29109));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n29107), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n29107), .I0(n2300), .I1(n2324), .CO(n29108));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n29106), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_29 (.CI(n28034), .I0(timer[27]), .I1(n1[27]), 
            .CO(n28035));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n29301), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n28033), .O(one_wire_N_513[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_26 (.CI(n29301), .I0(n3086), .I1(n3116), .CO(n29302));
    SB_CARRY sub_14_add_2_28 (.CI(n28033), .I0(timer[26]), .I1(n1[26]), 
            .CO(n28034));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n28032), .O(one_wire_N_513[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n29300), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n29106), .I0(n2301), .I1(n2324), .CO(n29107));
    SB_CARRY sub_14_add_2_27 (.CI(n28032), .I0(timer[25]), .I1(n1[25]), 
            .CO(n28033));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n28031), .O(one_wire_N_513[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n28031), .I0(timer[24]), .I1(n1[24]), 
            .CO(n28032));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n29105), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n29105), .I0(n2302), .I1(n2324), .CO(n29106));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_513[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n28030), .O(n30_adj_4558)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2143_25 (.CI(n29300), .I0(n3087), .I1(n3116), .CO(n29301));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n29104), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n29104), .I0(n2303), .I1(n2324), .CO(n29105));
    SB_CARRY sub_14_add_2_25 (.CI(n28030), .I0(timer[23]), .I1(n1[23]), 
            .CO(n28031));
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_513[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n28029), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n28029), .I0(timer[22]), .I1(n1[22]), 
            .CO(n28030));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_513[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n28028), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n28028), .I0(timer[21]), .I1(n1[21]), 
            .CO(n28029));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_513[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n28027), .O(n29_adj_4557)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n28027), .I0(timer[20]), .I1(n1[20]), 
            .CO(n28028));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n28026), .O(one_wire_N_513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_21 (.CI(n28026), .I0(timer[19]), .I1(n1[19]), 
            .CO(n28027));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n28025), .O(one_wire_N_513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n28025), .I0(timer[18]), .I1(n1[18]), 
            .CO(n28026));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_513[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n28024), .O(n27_adj_4554)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n29299), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n28024), .I0(timer[17]), .I1(n1[17]), 
            .CO(n28025));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n29103), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n28023), .O(one_wire_N_513[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n28023), .I0(timer[16]), .I1(n1[16]), 
            .CO(n28024));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n28022), .O(one_wire_N_513[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n28022), .I0(timer[15]), .I1(n1[15]), 
            .CO(n28023));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n28021), .O(one_wire_N_513[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n28021), .I0(timer[14]), .I1(n1[14]), 
            .CO(n28022));
    SB_CARRY mod_5_add_1607_8 (.CI(n29103), .I0(n2304), .I1(n2324), .CO(n29104));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n28020), .O(one_wire_N_513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n28020), .I0(timer[13]), .I1(n1[13]), 
            .CO(n28021));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n28019), .O(one_wire_N_513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n28019), .I0(timer[12]), .I1(n1[12]), 
            .CO(n28020));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n28018), .O(\one_wire_N_513[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n28018), .I0(timer[11]), .I1(n1[11]), 
            .CO(n28019));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n28017), .O(\one_wire_N_513[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n28017), .I0(timer[10]), .I1(n1[10]), 
            .CO(n28018));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n28016), .O(\one_wire_N_513[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n28016), .I0(timer[9]), .I1(n1[9]), 
            .CO(n28017));
    SB_CARRY mod_5_add_2143_24 (.CI(n29299), .I0(n3088), .I1(n3116), .CO(n29300));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n29102), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n29102), .I0(n2305), .I1(n2324), .CO(n29103));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n29101), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n28015), .O(\one_wire_N_513[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n28015), .I0(timer[8]), .I1(n1[8]), 
            .CO(n28016));
    SB_CARRY mod_5_add_1607_6 (.CI(n29101), .I0(n2306), .I1(n2324), .CO(n29102));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n29100), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n28014), .O(\one_wire_N_513[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n29298), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n29100), .I0(n2307), .I1(n2324), .CO(n29101));
    SB_CARRY sub_14_add_2_9 (.CI(n28014), .I0(timer[7]), .I1(n1[7]), .CO(n28015));
    SB_CARRY mod_5_add_2143_23 (.CI(n29298), .I0(n3089), .I1(n3116), .CO(n29299));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n28013), .O(\one_wire_N_513[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n28013), .I0(timer[6]), .I1(n1[6]), .CO(n28014));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n28012), .O(\one_wire_N_513[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n28012), .I0(timer[5]), .I1(n1[5]), .CO(n28013));
    SB_CARRY add_21_8 (.CI(n27753), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27754));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n28011), .O(one_wire_N_513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n29099), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_6 (.CI(n28011), .I0(timer[4]), .I1(n1[4]), .CO(n28012));
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n27765), 
            .O(n40239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n29297), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n27765), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27766));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27748));
    SB_CARRY mod_5_add_1607_4 (.CI(n29099), .I0(n2308), .I1(n2324), .CO(n29100));
    SB_LUT4 i9_4_lut_adj_1608 (.I0(n1701), .I1(n1708), .I2(n1707), .I3(n1700), 
            .O(n22_adj_4579));
    defparam i9_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1609 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n15_adj_4580));
    defparam i2_3_lut_adj_1609.LUT_INIT = 16'hecec;
    SB_LUT4 i7_3_lut (.I0(n1703), .I1(n1698), .I2(n1705), .I3(GND_net), 
            .O(n20_adj_4581));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1610 (.I0(n15_adj_4580), .I1(n22_adj_4579), .I2(n1704), 
            .I3(n1706), .O(n24_adj_4582));
    defparam i11_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1611 (.I0(n1697), .I1(n24_adj_4582), .I2(n20_adj_4581), 
            .I3(n1702), .O(n1730));
    defparam i12_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i36333_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43163));
    defparam i36333_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36319_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43149));
    defparam i36319_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4583));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1612 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4584));
    defparam i15_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i19858_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24584));
    defparam i19858_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1613 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24584), 
            .O(n36_adj_4585));
    defparam i13_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1614 (.I0(n2700), .I1(n38_adj_4584), .I2(n28_adj_4583), 
            .I3(n2705), .O(n42_adj_4586));
    defparam i19_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1615 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4587));
    defparam i17_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1616 (.I0(n2687), .I1(n36_adj_4585), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4588));
    defparam i18_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1617 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39));
    defparam i16_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i19720_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24446));
    defparam i19720_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1618 (.I0(n1405), .I1(n24446), .I2(n1401), .I3(n1406), 
            .O(n16_adj_4589));
    defparam i6_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1619 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4590));
    defparam i7_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1620 (.I0(n17_adj_4590), .I1(n1408), .I2(n16_adj_4589), 
            .I3(n1403), .O(n1433));
    defparam i9_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41_adj_4588), .I2(n40_adj_4587), 
            .I3(n42_adj_4586), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36318_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43148));
    defparam i36318_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1621 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4591));
    defparam i10_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1622 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4592));
    defparam i8_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1623 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4593));
    defparam i9_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1624 (.I0(bit_ctr[11]), .I1(n2399), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4594));
    defparam i7_3_lut_adj_1624.LUT_INIT = 16'hecec;
    SB_LUT4 i7_3_lut_adj_1625 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4595));
    defparam i7_3_lut_adj_1625.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1626 (.I0(n2392), .I1(n2390), .I2(n2394), .I3(n2407), 
            .O(n33_adj_4596));
    defparam i13_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1627 (.I0(n2396), .I1(n2401), .I2(n2403), .I3(n2400), 
            .O(n32_adj_4597));
    defparam i12_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1628 (.I0(n2406), .I1(n2405), .I2(n2391), .I3(n2402), 
            .O(n31_adj_4598));
    defparam i11_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1629 (.I0(n2393), .I1(n2397), .I2(n2408), .I3(n2395), 
            .O(n35));
    defparam i15_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1630 (.I0(n33_adj_4596), .I1(n27_adj_4594), .I2(n2404), 
            .I3(n2398), .O(n37_adj_4599));
    defparam i17_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1631 (.I0(n21_adj_4595), .I1(n23_adj_4593), .I2(n22_adj_4592), 
            .I3(n24_adj_4591), .O(n1829));
    defparam i13_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1632 (.I0(n37_adj_4599), .I1(n35), .I2(n31_adj_4598), 
            .I3(n32_adj_4597), .O(n2423));
    defparam i19_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_3_lut (.I0(bit_ctr[4]), .I1(n3101), .I2(n3109), .I3(GND_net), 
            .O(n37_adj_4600));
    defparam i10_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1633 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4601));
    defparam i16_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1634 (.I0(n3091), .I1(n3094), .I2(n3106), .I3(n3096), 
            .O(n45_adj_4602));
    defparam i18_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1635 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4603));
    defparam i14_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1636 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4604));
    defparam i15_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1637 (.I0(n3089), .I1(n3105), .I2(n3107), .I3(n3100), 
            .O(n42_adj_4605));
    defparam i15_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i36331_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43161));
    defparam i36331_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut_adj_1638 (.I0(n3097), .I1(n3092), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4606));
    defparam i5_2_lut_adj_1638.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1639 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4607));
    defparam i13_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1640 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4608));
    defparam i18_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1641 (.I0(n37_adj_4607), .I1(n39_adj_4604), .I2(n38_adj_4603), 
            .I3(n40_adj_4601), .O(n46_adj_4609));
    defparam i22_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4610));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4610), .I1(n46_adj_4609), .I2(n42_adj_4608), 
            .I3(n34), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36316_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43146));
    defparam i36316_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(n1301), .I1(n1302), .I2(bit_ctr[22]), .I3(n1309), 
            .O(n14_adj_4611));
    defparam i5_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i36315_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43145));
    defparam i36315_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1642 (.I0(n1304), .I1(n1305), .I2(n1306), .I3(n1307), 
            .O(n15_adj_4612));
    defparam i6_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1643 (.I0(n15_adj_4612), .I1(n1308), .I2(n14_adj_4611), 
            .I3(n1303), .O(n1334));
    defparam i8_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i36327_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43157));
    defparam i36327_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1644 (.I0(n3098), .I1(n3084), .I2(n3099), .I3(n3083), 
            .O(n44_adj_4613));
    defparam i17_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i36330_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43160));
    defparam i36330_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1645 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4614));
    defparam i6_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1646 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4615));
    defparam i1_3_lut_adj_1646.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1647 (.I0(n9_adj_4615), .I1(n14_adj_4614), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1648 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4616));
    defparam i11_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i36329_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43159));
    defparam i36329_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1649 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4617));
    defparam i4_3_lut_adj_1649.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1650 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4618));
    defparam i1_2_lut_adj_1650.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1651 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4619));
    defparam i9_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1652 (.I0(n19_adj_4617), .I1(n26_adj_4616), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4620));
    defparam i13_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1653 (.I0(n1896), .I1(n28_adj_4620), .I2(n24_adj_4619), 
            .I3(n16_adj_4618), .O(n1928));
    defparam i14_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i19432_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24154));
    defparam i19432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1654 (.I0(n1105), .I1(n1103), .I2(n24154), .I3(n1108), 
            .O(n12_adj_4621));
    defparam i5_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1655 (.I0(n1107), .I1(n12_adj_4621), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i36314_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43144));
    defparam i36314_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36328_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43158));
    defparam i36328_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36298_2_lut (.I0(n31265), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i36298_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i36300_2_lut (.I0(n31265), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i36300_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n31265), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31336_3_lut (.I0(n905), .I1(n906), .I2(n35416), .I3(GND_net), 
            .O(n38102));
    defparam i31336_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n38102), .I2(n17101), .I3(n14346), 
            .O(n31265));
    defparam i4_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n31265), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14346), .I1(n971[27]), .I2(n31265), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31357_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n38124));
    defparam i31357_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1656 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4622));
    defparam i2_3_lut_adj_1656.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1657 (.I0(n31265), .I1(n6_adj_4622), .I2(n1005), 
            .I3(n38124), .O(n1037));
    defparam i3_4_lut_adj_1657.LUT_INIT = 16'hfdfc;
    SB_LUT4 i36296_2_lut (.I0(n31265), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4578));   // verilog/neopixel.v(22[26:36])
    defparam i36296_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i9_3_lut_adj_1658 (.I0(bit_ctr[6]), .I1(n2904), .I2(n2909), 
            .I3(GND_net), .O(n34_adj_4623));
    defparam i9_3_lut_adj_1658.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1659 (.I0(n2897), .I1(n2905), .I2(n2895), .I3(n2901), 
            .O(n41_adj_4624));
    defparam i16_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2885), .I3(GND_net), 
            .O(n38_adj_4625));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1660 (.I0(n2898), .I1(n2902), .I2(n2907), .I3(n2903), 
            .O(n43_adj_4626));
    defparam i18_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1661 (.I0(n2888), .I1(n2890), .I2(n2894), .I3(n2908), 
            .O(n40_adj_4627));
    defparam i15_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1662 (.I0(n41_adj_4624), .I1(n2896), .I2(n34_adj_4623), 
            .I3(n2899), .O(n46_adj_4628));
    defparam i21_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1663 (.I0(n2893), .I1(n2886), .I2(n2892), .I3(n2889), 
            .O(n39_adj_4629));
    defparam i14_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1664 (.I0(n43_adj_4626), .I1(n2891), .I2(n38_adj_4625), 
            .I3(n2900), .O(n47_adj_4630));
    defparam i22_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1665 (.I0(n47_adj_4630), .I1(n39_adj_4629), .I2(n46_adj_4628), 
            .I3(n40_adj_4627), .O(n2918));
    defparam i24_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 i36312_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43142));
    defparam i36312_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1666 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4631));
    defparam i2_2_lut_adj_1666.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1667 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4632));
    defparam i12_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1668 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4633));
    defparam i10_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1669 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4634));
    defparam i11_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1670 (.I0(bit_ctr[15]), .I1(n18_adj_4631), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4635));
    defparam i9_4_lut_adj_1670.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1671 (.I0(n25_adj_4635), .I1(n27_adj_4634), .I2(n26_adj_4633), 
            .I3(n28_adj_4632), .O(n2027));
    defparam i15_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i36313_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43143));
    defparam i36313_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4636));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1672 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4637));
    defparam i13_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1673 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4638));
    defparam i1_3_lut_adj_1673.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1674 (.I0(n2490), .I1(n34_adj_4637), .I2(n24_adj_4636), 
            .I3(n2494), .O(n38_adj_4639));
    defparam i17_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1675 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4640));
    defparam i15_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1676 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4638), 
            .O(n37_adj_4641));
    defparam i16_4_lut_adj_1676.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1677 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4642));
    defparam i14_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1678 (.I0(n35_adj_4642), .I1(n37_adj_4641), .I2(n36_adj_4640), 
            .I3(n38_adj_4639), .O(n2522));
    defparam i20_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1679 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4643));
    defparam i3_2_lut_adj_1679.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1680 (.I0(bit_ctr[12]), .I1(n22_adj_4643), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4644));
    defparam i11_4_lut_adj_1680.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1681 (.I0(n2294), .I1(n30_adj_4644), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4645));
    defparam i15_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1682 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4646));
    defparam i13_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1683 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4647));
    defparam i14_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1684 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4648));
    defparam i12_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1685 (.I0(n45_adj_4602), .I1(n37_adj_4600), .I2(n3087), 
            .I3(n3088), .O(n50_adj_4649));
    defparam i23_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1686 (.I0(n31_adj_4648), .I1(n33_adj_4647), .I2(n32_adj_4646), 
            .I3(n34_adj_4645), .O(n2324));
    defparam i18_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1687 (.I0(n3102), .I1(n42_adj_4605), .I2(n3108), 
            .I3(n3093), .O(n48_adj_4650));
    defparam i21_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1688 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14346));
    defparam i1_2_lut_adj_1688.LUT_INIT = 16'h9999;
    SB_LUT4 i36310_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43140));
    defparam i36310_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36325_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43155));
    defparam i36325_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_2_lut_adj_1689 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n14348));
    defparam i1_2_lut_adj_1689.LUT_INIT = 16'h6666;
    SB_LUT4 i34046_3_lut (.I0(n30411), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n35303));
    defparam i34046_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n35313), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i28686_2_lut (.I0(one_wire_N_513[4]), .I1(n35373), .I2(GND_net), 
            .I3(GND_net), .O(n35452));
    defparam i28686_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i130_4_lut (.I0(n24408), .I1(n35476), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n103));
    defparam i130_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n35462), .I1(n35452), .I2(n4_adj_4550), 
            .I3(n34689), .O(n34609));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'h1505;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n15824), .I1(\state[0] ), .I2(n34609), 
            .I3(n103), .O(n16961));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'h5150;
    SB_LUT4 i96_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_576 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i96_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19736_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n24462));
    defparam i19736_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1692 (.I0(n3184), .I1(n3182), .I2(n3201), .I3(n3200), 
            .O(n48_adj_4651));
    defparam i20_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1693 (.I0(n3204), .I1(n3203), .I2(n3187), .I3(n3207), 
            .O(n46_adj_4652));
    defparam i18_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1694 (.I0(n3188), .I1(n3194), .I2(n3208), .I3(n3196), 
            .O(n47_adj_4653));
    defparam i19_4_lut_adj_1694.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1695 (.I0(n3186), .I1(n3195), .I2(n3205), .I3(n3191), 
            .O(n45_adj_4654));
    defparam i17_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1696 (.I0(n3183), .I1(n3199), .I2(n3197), .I3(n24462), 
            .O(n44_adj_4655));
    defparam i16_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1697 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n3206), 
            .O(n43_adj_4656));
    defparam i15_4_lut_adj_1697.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1698 (.I0(n45_adj_4654), .I1(n47_adj_4653), .I2(n46_adj_4652), 
            .I3(n48_adj_4651), .O(n54_adj_4657));
    defparam i26_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1699 (.I0(n3190), .I1(n3192), .I2(n3185), .I3(n3202), 
            .O(n49_adj_4658));
    defparam i21_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1700 (.I0(n49_adj_4658), .I1(n54_adj_4657), .I2(n43_adj_4656), 
            .I3(n44_adj_4655), .O(n24464));
    defparam i27_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 color_bit_I_0_i2_3_lut (.I0(\color[2] ), .I1(\color[3] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n2_adj_4659));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1701 (.I0(bit_ctr[0]), .I1(\color[4] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4660));
    defparam i1_2_lut_adj_1701.LUT_INIT = 16'h4444;
    SB_LUT4 i34358_4_lut (.I0(\color[1] ), .I1(n2_adj_4659), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n41190));   // verilog/neopixel.v(22[26:36])
    defparam i34358_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 color_bit_I_0_i7_4_lut (.I0(n41190), .I1(bit_ctr[1]), .I2(bit_ctr[2]), 
            .I3(n4_adj_4660), .O(n7_adj_4661));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i7_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i31320_4_lut (.I0(\state_3__N_362[1] ), .I1(n3209), .I2(bit_ctr[3]), 
            .I3(n24464), .O(n38086));
    defparam i31320_4_lut.LUT_INIT = 16'hbeee;
    SB_LUT4 i3_4_lut_adj_1702 (.I0(n38086), .I1(n7_adj_4661), .I2(bit_ctr[3]), 
            .I3(n24464), .O(state_3__N_362[0]));
    defparam i3_4_lut_adj_1702.LUT_INIT = 16'h4004;
    SB_LUT4 i22_4_lut_adj_1703 (.I0(n3085), .I1(n44_adj_4613), .I2(n32_adj_4606), 
            .I3(n3095), .O(n49_adj_4662));
    defparam i22_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i36324_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43154));
    defparam i36324_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19682_3_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(GND_net), .O(n24408));
    defparam i19682_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i237_2_lut (.I0(n24520), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1169));   // verilog/neopixel.v(103[9] 111[12])
    defparam i237_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(\state[0] ), .I1(n13389), .I2(n1169), 
            .I3(\state[1] ), .O(n17008));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'haf33;
    SB_LUT4 i15_4_lut_adj_1705 (.I0(n13389), .I1(n1169), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n35420));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1705.LUT_INIT = 16'h0535;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(GND_net), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 i1_2_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(GND_net), .O(n30411));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h9292;
    SB_LUT4 i1_2_lut_3_lut (.I0(n35424), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n13389));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i19794_2_lut_4_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(n15824), .O(n24520));
    defparam i19794_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i28710_2_lut_3_lut (.I0(n35462), .I1(one_wire_N_513[4]), .I2(n35373), 
            .I3(GND_net), .O(n35476));
    defparam i28710_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i34051_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17101));
    defparam i34051_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_LUT4 i2804_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n35303), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i2804_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 i2_3_lut_4_lut (.I0(n35424), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(\state[1] ), .O(n35991));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i23_3_lut_4_lut (.I0(n24324), .I1(one_wire_N_513[4]), .I2(n29824), 
            .I3(\state[0] ), .O(n35335));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 mux_668_Mux_0_i3_3_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_668_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34738));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36323_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43153));
    defparam i36323_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1706 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4663));
    defparam i14_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_4664));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1707 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4665));
    defparam i12_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1708 (.I0(n25_adj_4664), .I1(n36_adj_4663), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4666));
    defparam i18_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1709 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4667));
    defparam i16_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4665), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4668));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1710 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4669));
    defparam i15_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1711 (.I0(n37_adj_4669), .I1(n39_adj_4668), .I2(n38_adj_4667), 
            .I3(n40_adj_4666), .O(n2621));
    defparam i21_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i36320_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43150));
    defparam i36320_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(n29824), .I1(n15631), .I2(\neo_pixel_transmitter.done ), 
            .I3(start), .O(n1166));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff1f;
    SB_LUT4 i1_3_lut_4_lut (.I0(n15631), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n4_adj_4550), .O(n15745));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i20_4_lut_adj_1712 (.I0(n3103), .I1(n3086), .I2(n3104), .I3(n3090), 
            .O(n47_adj_4670));
    defparam i20_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n739));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h49db;
    SB_LUT4 i26_4_lut_adj_1713 (.I0(n47_adj_4670), .I1(n49_adj_4662), .I2(n48_adj_4650), 
            .I3(n50_adj_4649), .O(n3116));
    defparam i26_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, \data_in_frame[5] , GND_net, n34179, byte_transmit_counter, 
            n34135, n18046, setpoint, n18047, \data_in_frame[12] , 
            n34037, n34001, n34177, \byte_transmit_counter[1] , n18057, 
            n18058, n18059, n18060, n18048, n18049, n18050, n18051, 
            n18052, n18053, n18054, n18055, n18056, n43329, n18042, 
            n18043, n18044, n18045, n18040, n18041, n18038, n18039, 
            n17960, PWMLimit, n17961, n17936, \data_in_frame[24] , 
            n17937, n17938, n17939, n17940, n17941, n17942, \data_in_frame[21] , 
            n17962, n17963, n17964, n17965, \data_in_frame[20] , n17956, 
            n17957, n17958, n17959, n17954, n17955, n17952, n17953, 
            n17950, n17951, n17948, n17949, n17946, n17947, n17943, 
            n17944, n17945, n17935, \data_in_frame[22] , \data_in_frame[4] , 
            \data_in_frame[11] , \data_in_frame[3] , \data_in_frame[2] , 
            \FRAME_MATCHER.state[1] , \data_out_frame[5] , \data_out_frame[6] , 
            \data_out_frame[7] , \byte_transmit_counter[0] , rx_data, 
            \data_in_frame[1] , \data_in_frame[2][0] , \data_in_frame[2][2] , 
            n17743, control_mode, n17742, n17741, n17740, n17739, 
            n17738, n17737, n17736, \data_out_frame[20] , n17735, 
            \data_in_frame[10] , n17734, rx_data_ready, n17733, n17732, 
            tx_active, n63, n17731, n17730, n17729, n17728, \data_out_frame[19] , 
            n17727, n17726, n17725, n17724, n17723, n17722, n17721, 
            n17720, \data_out_frame[18] , n17719, n17718, n17717, 
            n17716, n17714, \data_out_frame[18][1] , n17713, \data_out_frame[18][0] , 
            n17712, \data_out_frame[17] , n17711, n17710, \data_in_frame[13] , 
            n17709, n17708, n17707, n17706, n17705, n17704, \data_out_frame[16] , 
            n17703, n17702, n17701, n17700, n17699, n17698, n17697, 
            n17696, \data_out_frame[15] , n17695, n17694, n17693, 
            n17692, n17691, n17690, n17689, n17688, \data_out_frame[14] , 
            n17687, n17686, n17685, n17684, n17683, n17682, n17681, 
            n17680, \data_out_frame[13] , n17679, n17678, n17677, 
            n17676, n17675, n17674, n17673, n17672, \data_out_frame[12] , 
            n17671, n17670, n17669, n17668, n17667, n17666, n17665, 
            n17664, \data_out_frame[11] , n17663, n17662, n17661, 
            n17660, n17659, n17658, n17657, n17656, \data_out_frame[10] , 
            n17655, n17654, n17653, n17652, n17651, n17650, n17649, 
            n17648, \data_out_frame[9] , n17647, n17646, n17645, n17644, 
            n17643, n17642, n17641, n17640, \data_out_frame[8] , n17639, 
            n17638, n17637, n17636, n17635, n17634, n17633, n17632, 
            n17631, n17630, n17629, n17628, n17627, n17626, n17625, 
            n17624, n17623, n17622, n17621, n17620, n17619, n17618, 
            n17617, n17616, n17615, n17614, n17613, n17612, n17611, 
            n17610, n17609, n17608, \data_in[3] , n17607, n17606, 
            n17605, n17604, n17603, n17602, n17601, n17600, \data_in[2] , 
            n17599, n17598, n17597, n17596, n17595, n17594, n17593, 
            n17592, \data_in[1] , n17591, n17590, n17589, n17588, 
            n17587, n17586, n17585, n17584, \data_in[0] , n17583, 
            n17582, n17581, n17580, n17579, n17578, n17577, \Ki[15] , 
            n17576, \Ki[14] , n17575, \Ki[13] , n17574, \Ki[12] , 
            n17573, \Ki[11] , n17572, \Ki[10] , n30070, n17571, 
            \Ki[9] , n17570, \Ki[8] , n17569, \Ki[7] , n17568, \Ki[6] , 
            n17567, \Ki[5] , n17566, \Ki[4] , n17565, \Ki[3] , n17564, 
            \Ki[2] , n17563, \Ki[1] , n17562, \Kp[15] , n17561, 
            \Kp[14] , n17560, \Kp[13] , n17559, \Kp[12] , n17558, 
            \Kp[11] , n17557, \Kp[10] , \Kp[9] , n17555, \Kp[8] , 
            n17554, \Kp[7] , n17553, \Kp[6] , n17552, \Kp[5] , n17551, 
            \Kp[4] , n17550, \Kp[3] , n17549, \Kp[2] , n17548, \Kp[1] , 
            n17547, gearBoxRatio, n4351, n17546, n17545, n17544, 
            n17543, n17542, n4350, \data_in_frame[9] , n17541, n17540, 
            n17539, n17538, n17537, n17536, n17535, n4353, n17534, 
            n17533, n4352, n17532, n17531, n17530, n17529, n17528, 
            n17527, n4357, n17526, n17525, n17523, IntegralLimit, 
            n17522, n4356, n4355, n4354, n17521, n17520, n17519, 
            n788, n17518, n17517, n17516, n17515, n17514, n17513, 
            n17512, n17511, n17510, n17509, n17508, n122, n9001, 
            n34675, \FRAME_MATCHER.i_31__N_2621 , n17507, n17506, n3894, 
            n17505, n5, n17504, n17503, n17502, n17501, n34173, 
            n4368, n4367, n4366, n4365, n4364, n4363, n4362, n4361, 
            n4360, n17417, n4372, n4371, \data_in_frame[8] , n4370, 
            LED_c, n4369, n34067, n17398, n17396, n17395, n17394, 
            \Ki[0] , n17393, \Kp[0] , n17392, \FRAME_MATCHER.i_31__N_2625 , 
            n17249, n40273, n40274, n40275, n40278, n40277, n40276, 
            n36887, n24391, n4359, \displacement[18] , n13263, \FRAME_MATCHER.state_31__N_2661[2] , 
            n7, \FRAME_MATCHER.state_31__N_2661[0] , n4349, n2957, n36881, 
            n4358, n17314, r_Bit_Index, n17311, r_SM_Main, n17446, 
            n17412, n17411, n17410, tx_o, VCC_net, \r_SM_Main_2__N_3579[1] , 
            n17058, n43694, n4670, n17189, n4, n3, n8936, n10627, 
            tx_enable, n17338, r_Bit_Index_adj_11, n17341, n24450, 
            \r_SM_Main[1]_adj_6 , r_Rx_Data, PIN_13_N_105, \r_SM_Main[2]_adj_7 , 
            n40218, n40217, n17452, n17462, n4_adj_8, n17429, n17428, 
            n17427, n17426, n17425, n17403, n17052, n17180, n4648, 
            n17343, n17342, n43211, n15734, n15626, n23653, n4_adj_9, 
            n4_adj_10) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    output [7:0]\data_in_frame[5] ;
    input GND_net;
    input n34179;
    output [7:0]byte_transmit_counter;
    input n34135;
    input n18046;
    output [23:0]setpoint;
    input n18047;
    output [7:0]\data_in_frame[12] ;
    input n34037;
    input n34001;
    input n34177;
    output \byte_transmit_counter[1] ;
    input n18057;
    input n18058;
    input n18059;
    input n18060;
    input n18048;
    input n18049;
    input n18050;
    input n18051;
    input n18052;
    input n18053;
    input n18054;
    input n18055;
    input n18056;
    input n43329;
    input n18042;
    input n18043;
    input n18044;
    input n18045;
    input n18040;
    input n18041;
    input n18038;
    input n18039;
    input n17960;
    output [23:0]PWMLimit;
    input n17961;
    input n17936;
    output [7:0]\data_in_frame[24] ;
    input n17937;
    input n17938;
    input n17939;
    input n17940;
    input n17941;
    input n17942;
    output [7:0]\data_in_frame[21] ;
    input n17962;
    input n17963;
    input n17964;
    input n17965;
    output [7:0]\data_in_frame[20] ;
    input n17956;
    input n17957;
    input n17958;
    input n17959;
    input n17954;
    input n17955;
    input n17952;
    input n17953;
    input n17950;
    input n17951;
    input n17948;
    input n17949;
    input n17946;
    input n17947;
    input n17943;
    input n17944;
    input n17945;
    input n17935;
    output [7:0]\data_in_frame[22] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[2] ;
    output \FRAME_MATCHER.state[1] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output \byte_transmit_counter[0] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[1] ;
    output \data_in_frame[2][0] ;
    output \data_in_frame[2][2] ;
    input n17743;
    output [7:0]control_mode;
    input n17742;
    input n17741;
    input n17740;
    input n17739;
    input n17738;
    input n17737;
    input n17736;
    output [7:0]\data_out_frame[20] ;
    input n17735;
    output [7:0]\data_in_frame[10] ;
    input n17734;
    output rx_data_ready;
    input n17733;
    input n17732;
    output tx_active;
    output n63;
    input n17731;
    input n17730;
    input n17729;
    input n17728;
    output [7:0]\data_out_frame[19] ;
    input n17727;
    input n17726;
    input n17725;
    input n17724;
    input n17723;
    input n17722;
    input n17721;
    input n17720;
    output [7:0]\data_out_frame[18] ;
    input n17719;
    input n17718;
    input n17717;
    input n17716;
    input n17714;
    output \data_out_frame[18][1] ;
    input n17713;
    output \data_out_frame[18][0] ;
    input n17712;
    output [7:0]\data_out_frame[17] ;
    input n17711;
    input n17710;
    output [7:0]\data_in_frame[13] ;
    input n17709;
    input n17708;
    input n17707;
    input n17706;
    input n17705;
    input n17704;
    output [7:0]\data_out_frame[16] ;
    input n17703;
    input n17702;
    input n17701;
    input n17700;
    input n17699;
    input n17698;
    input n17697;
    input n17696;
    output [7:0]\data_out_frame[15] ;
    input n17695;
    input n17694;
    input n17693;
    input n17692;
    input n17691;
    input n17690;
    input n17689;
    input n17688;
    output [7:0]\data_out_frame[14] ;
    input n17687;
    input n17686;
    input n17685;
    input n17684;
    input n17683;
    input n17682;
    input n17681;
    input n17680;
    output [7:0]\data_out_frame[13] ;
    input n17679;
    input n17678;
    input n17677;
    input n17676;
    input n17675;
    input n17674;
    input n17673;
    input n17672;
    output [7:0]\data_out_frame[12] ;
    input n17671;
    input n17670;
    input n17669;
    input n17668;
    input n17667;
    input n17666;
    input n17665;
    input n17664;
    output [7:0]\data_out_frame[11] ;
    input n17663;
    input n17662;
    input n17661;
    input n17660;
    input n17659;
    input n17658;
    input n17657;
    input n17656;
    output [7:0]\data_out_frame[10] ;
    input n17655;
    input n17654;
    input n17653;
    input n17652;
    input n17651;
    input n17650;
    input n17649;
    input n17648;
    output [7:0]\data_out_frame[9] ;
    input n17647;
    input n17646;
    input n17645;
    input n17644;
    input n17643;
    input n17642;
    input n17641;
    input n17640;
    output [7:0]\data_out_frame[8] ;
    input n17639;
    input n17638;
    input n17637;
    input n17636;
    input n17635;
    input n17634;
    input n17633;
    input n17632;
    input n17631;
    input n17630;
    input n17629;
    input n17628;
    input n17627;
    input n17626;
    input n17625;
    input n17624;
    input n17623;
    input n17622;
    input n17621;
    input n17620;
    input n17619;
    input n17618;
    input n17617;
    input n17616;
    input n17615;
    input n17614;
    input n17613;
    input n17612;
    input n17611;
    input n17610;
    input n17609;
    input n17608;
    output [7:0]\data_in[3] ;
    input n17607;
    input n17606;
    input n17605;
    input n17604;
    input n17603;
    input n17602;
    input n17601;
    input n17600;
    output [7:0]\data_in[2] ;
    input n17599;
    input n17598;
    input n17597;
    input n17596;
    input n17595;
    input n17594;
    input n17593;
    input n17592;
    output [7:0]\data_in[1] ;
    input n17591;
    input n17590;
    input n17589;
    input n17588;
    input n17587;
    input n17586;
    input n17585;
    input n17584;
    output [7:0]\data_in[0] ;
    input n17583;
    input n17582;
    input n17581;
    input n17580;
    input n17579;
    input n17578;
    input n17577;
    output \Ki[15] ;
    input n17576;
    output \Ki[14] ;
    input n17575;
    output \Ki[13] ;
    input n17574;
    output \Ki[12] ;
    input n17573;
    output \Ki[11] ;
    input n17572;
    output \Ki[10] ;
    output n30070;
    input n17571;
    output \Ki[9] ;
    input n17570;
    output \Ki[8] ;
    input n17569;
    output \Ki[7] ;
    input n17568;
    output \Ki[6] ;
    input n17567;
    output \Ki[5] ;
    input n17566;
    output \Ki[4] ;
    input n17565;
    output \Ki[3] ;
    input n17564;
    output \Ki[2] ;
    input n17563;
    output \Ki[1] ;
    input n17562;
    output \Kp[15] ;
    input n17561;
    output \Kp[14] ;
    input n17560;
    output \Kp[13] ;
    input n17559;
    output \Kp[12] ;
    input n17558;
    output \Kp[11] ;
    input n17557;
    output \Kp[10] ;
    output \Kp[9] ;
    input n17555;
    output \Kp[8] ;
    input n17554;
    output \Kp[7] ;
    input n17553;
    output \Kp[6] ;
    input n17552;
    output \Kp[5] ;
    input n17551;
    output \Kp[4] ;
    input n17550;
    output \Kp[3] ;
    input n17549;
    output \Kp[2] ;
    input n17548;
    output \Kp[1] ;
    input n17547;
    output [23:0]gearBoxRatio;
    output n4351;
    input n17546;
    input n17545;
    input n17544;
    input n17543;
    input n17542;
    output n4350;
    output [7:0]\data_in_frame[9] ;
    input n17541;
    input n17540;
    input n17539;
    input n17538;
    input n17537;
    input n17536;
    input n17535;
    output n4353;
    input n17534;
    input n17533;
    output n4352;
    input n17532;
    input n17531;
    input n17530;
    input n17529;
    input n17528;
    input n17527;
    output n4357;
    input n17526;
    input n17525;
    input n17523;
    output [23:0]IntegralLimit;
    input n17522;
    output n4356;
    output n4355;
    output n4354;
    input n17521;
    input n17520;
    input n17519;
    output n788;
    input n17518;
    input n17517;
    input n17516;
    input n17515;
    input n17514;
    input n17513;
    input n17512;
    input n17511;
    input n17510;
    input n17509;
    input n17508;
    output n122;
    output n9001;
    output n34675;
    output \FRAME_MATCHER.i_31__N_2621 ;
    input n17507;
    input n17506;
    output n3894;
    input n17505;
    output n5;
    input n17504;
    input n17503;
    input n17502;
    input n17501;
    input n34173;
    output n4368;
    output n4367;
    output n4366;
    output n4365;
    output n4364;
    output n4363;
    output n4362;
    output n4361;
    output n4360;
    input n17417;
    output n4372;
    output n4371;
    output [7:0]\data_in_frame[8] ;
    output n4370;
    output LED_c;
    output n4369;
    input n34067;
    input n17398;
    input n17396;
    input n17395;
    input n17394;
    output \Ki[0] ;
    input n17393;
    output \Kp[0] ;
    input n17392;
    output \FRAME_MATCHER.i_31__N_2625 ;
    input n17249;
    output n40273;
    output n40274;
    output n40275;
    output n40278;
    output n40277;
    output n40276;
    output n36887;
    output n24391;
    output n4359;
    input \displacement[18] ;
    output n13263;
    output \FRAME_MATCHER.state_31__N_2661[2] ;
    output n7;
    output \FRAME_MATCHER.state_31__N_2661[0] ;
    output n4349;
    output n2957;
    output n36881;
    output n4358;
    input n17314;
    output [2:0]r_Bit_Index;
    input n17311;
    output [2:0]r_SM_Main;
    input n17446;
    input n17412;
    input n17411;
    input n17410;
    output tx_o;
    input VCC_net;
    output \r_SM_Main_2__N_3579[1] ;
    output n17058;
    input n43694;
    output n4670;
    output n17189;
    output n4;
    output n3;
    output n8936;
    output n10627;
    output tx_enable;
    input n17338;
    output [2:0]r_Bit_Index_adj_11;
    input n17341;
    input n24450;
    output \r_SM_Main[1]_adj_6 ;
    output r_Rx_Data;
    input PIN_13_N_105;
    output \r_SM_Main[2]_adj_7 ;
    output n40218;
    output n40217;
    input n17452;
    input n17462;
    output n4_adj_8;
    input n17429;
    input n17428;
    input n17427;
    input n17426;
    input n17425;
    input n17403;
    output n17052;
    output n17180;
    output n4648;
    input n17343;
    input n17342;
    output n43211;
    output n15734;
    output n15626;
    output n23653;
    output n4_adj_9;
    output n4_adj_10;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n17900;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    
    wire n17899, n17898, n17897, n17896, n17895, n17894;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    
    wire n17893, n17892, n17891, n17890, n17889, n17888, n17790, 
        n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n3_c, n17887, n17886;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    
    wire n17885, n17884, n17789, n17883, n27809, n27810, n2_adj_4257, 
        n27808, n2060, n17804;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    
    wire n17803, n17802, n17801, n17800, n17799, n17798;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    
    wire n17797, n17796, n17844, n18093;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(100[12:33])
    
    wire n18094, n17843, n17842, n17841;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n17928;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(94[12:25])
    
    wire n17929, n17930, n17931, n17932, n17933, n17917, n17918, 
        n17795, n17788, n17787, n17901, n17902, n17903, n17786, 
        n17785, n17784, n17783, n17934, n17919, n17920, n17921, 
        n17922, n17923, n17924, n17925, n17926, n17927, n17782, 
        n17840, n17839, n17838, n17837, n17836, n17781, n17780, 
        n17915, n17916, n17913, n17914, n17911, n17912, n17909, 
        n17910, n17907, n17908, n17904, n17905, n17906, n17779, 
        n17778, n17777, n17776, n17775, n17774, n17773, n17772, 
        n17771, n17770, n17856;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n17835, n17834, n17769, n17794, n17768, n17793, n17767, 
        n17766, n17792, n17765, n17833, n17764, n17763, n17762, 
        n2_adj_4258, n27807, n24676, n34704, n24683, tx_transmit_N_3479, 
        n23565, n40143, n24684;
    wire [0:0]n3295;
    
    wire n17882, n40568, n5_c, n8, n34707, n40044, n38201, n43199, 
        n38203, n2_adj_4259, n27806;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(94[12:25])
    
    wire n38, n25;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n38112, n38114, n39, n43, n9, n38122;
    wire [31:0]\FRAME_MATCHER.state_31__N_2725 ;
    
    wire n17761, n17760, n17759, n17881, n17758, n17757, n17756, 
        n17755, n17754, n17753, n17752, n17751, n17750, n17749, 
        n17748, n17747, n17746, n17832, n17745, n17744, n17831, 
        n17830, n13355, n31, n31_adj_4260, n29, n35082, n34943, 
        n16448;
    wire [2:0]r_SM_Main_2__N_3582;
    
    wire n34694, \FRAME_MATCHER.rx_data_ready_prev , n17880, n15876, 
        n23620, n17879, n17878;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n17877, n17829, n17845, n17828, n17855, n17876, n17715;
    wire [7:0]\data_out_frame[18]_c ;   // verilog/coms.v(95[12:26])
    
    wire n2_adj_4261, n27805, n35063, n16033, n2_adj_4262, n27804, 
        n8_adj_4263, n34723, n17857, n17858, n2_adj_4264, n27803, 
        n17859, n17860, n2_adj_4265, n27802, n17861, n17862, n17854, 
        n17853, n2_adj_4266, n27801, n17852, n26, n17851, n17850, 
        n2_adj_4267, n27821, n2_adj_4268, n27820, n34961, n2_adj_4269, 
        n27819, n16427, n4_c, n16716, n34864, n16706, n34749, 
        n16666, n16663, n34900, n34978, n31329, n16292, n31129, 
        n31392, n6, n16053, n34806, n34786, n34800, n35227, n17849, 
        n2_adj_4270, n27800, n2_adj_4271, n27818, n2_adj_4272, n27817, 
        n2_adj_4273, n27799, n2_adj_4274, n27798, n34765, n17848, 
        n2_adj_4275, n27816, n34883, n29_adj_4276, n36028, n16, 
        n16430, n34880, n17, n2_adj_4277, n27815, n2_adj_4278, n27797, 
        n2_adj_4279, n27796, n2_adj_4280, n27814, n5_adj_4281, n2_adj_4282, 
        n27795, n17556, n4348, n8_adj_4283, n17815, n17816, n17817, 
        n17818, n17819, n17820, n4_adj_4284, n15839, n15645, n20, 
        n19, n17821, n38108, n63_adj_4285, n10, n14, n16_adj_4286, 
        n17_adj_4287, n15728, n10_adj_4288, n15741, n14_adj_4289, 
        n15, n16_adj_4290, n17_adj_4291, n63_adj_4292, n17822, n34948, 
        n10_adj_4293, n1713, n31414, n35100, n18, n20_adj_4294, 
        n15_adj_4295, n63_adj_4296, n16815, n31306, n15731, n15648, 
        n44, n42, n43_adj_4297, n41, n16742, n40, n39_adj_4298, 
        n50, n45, n7_c, n37049, n16299, n24610, n30545, n35233, 
        n12, n31381, n19504, n2774, n30491, n31281, n1211, n34790, 
        n34927, n15489, n6_adj_4300, n16760, n34940, n16029, n34991, 
        n34771, n16660, n31435, n10_adj_4301, n36954, n35025, n15422, 
        n35142, n6_adj_4302, n31390, n35057, n35058, n34994, n34995, 
        n31394, n35221, n10_adj_4303, n15426, n35781, n34906, n10_adj_4304;
    wire [31:0]n92;
    
    wire n34681, n29937, n34051, n10337, n50_adj_4305, n27214, n34065, 
        n34105, n2_adj_4306, n27813, n2_adj_4307, n27812, n27811, 
        n2_adj_4308, n27794, n34107, n2_adj_4309, n3_adj_4310, n17827, 
        n12_adj_4311, n28, n32, n34063, n34069, n34129, n17806, 
        n2_adj_4312, n2_adj_4313, n27793, n34109, n2_adj_4314, n27792, 
        n2_adj_4315, n34111, n17826, n17825, n27791, n17824, n17823, 
        n3_adj_4316, n24311, n3_adj_4317, n3_adj_4318, n3_adj_4319, 
        n3_adj_4320, n3_adj_4321, n3_adj_4322, n3_adj_4323, n3_adj_4324, 
        n3_adj_4325, n3_adj_4326, n3_adj_4327, n3_adj_4328, n3_adj_4329, 
        n3_adj_4330, n3_adj_4331, n3_adj_4332, n2_adj_4333, n3_adj_4334, 
        n3_adj_4335, n3_adj_4336, n3_adj_4337, n3_adj_4338, n3_adj_4339, 
        n3_adj_4340, n3_adj_4341, n3_adj_4342, n3_adj_4343, n3_adj_4344, 
        n3_adj_4345, n3_adj_4346, n37121, n17010;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n36413, n36072, n36454, n36358, n36643, n36919, n37102, 
        n34972;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n35055, n34964, n35194, n34829, n37115, n43574, n24309, 
        n34113, n34115, n34053, n34193, n23582, n34059, n34195, 
        n34055, n34197, n34127, n34199, n34125, n34201, n34123, 
        n34203, n34121, n23584, n24305, n34205, n34119, n23586, 
        n24307, n34207, n34117, n34209, n7_adj_4347, n8_adj_4348, 
        n34211, n23588, n23590, n34213, n34215, n7_adj_4349, n8_adj_4350, 
        n34187, n7_adj_4351, n8_adj_4352, n34221, n23592, n34217, 
        n7_adj_4353, n8_adj_4354, n34219, n7_adj_4355, n8_adj_4356, 
        n23594, n7_adj_4357, n8_adj_4358, n49, n37, n43298, n16641, 
        n6_adj_4359, n16382, n35179, n34955, n14_adj_4360, n10_adj_4361, 
        n31060, Kp_23__N_1186, n41_adj_4362, n36824, n36660, n6_adj_4363, 
        n8_adj_4364, n35006, n35022, n31439, n17875, n17874, n161, 
        n24351;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    
    wire n17863, n17864, n34837, n17865, n17866, n43301, n43292, 
        n43295, n43286, n43289, n43280, n43283, n43274, n43277, 
        n43268, n43271, n43262, n43265, n43256, n17873, n17872, 
        n17871, n17867, n17868, n17869, n17870, n10_adj_4365, n34697, 
        n17807, n17814, n17847, n17397, n17808, n17809, n17810, 
        n17811, n43259, n17812, n17813, n31141, n15435, n30525, 
        n35785, n30999, n31320, n31310, n31273, n14249, n6_adj_4366, 
        n27, n31368, n6_adj_4367, n27212, n35182, n34746, n35170, 
        n10_adj_4368, n31327, n31298, n34897, n17805, n38252, n38253, 
        n38256, n38255, n38246, n38247, n38250, n38249, n38240, 
        n38241, n38244, n38243, n16_adj_4369, n17_adj_4370, n40113, 
        n19_adj_4371, n16_adj_4372, n17_adj_4373, n40133, n19_adj_4374, 
        n38282, n38283, n38286, n38285, n34603, n19503, n43250, 
        n8_adj_4375, n43253, n8_adj_4376, n17846, n17791, n40145, 
        n27854, n40179, n27853, \FRAME_MATCHER.i_31__N_2624 , n27852, 
        n27851, n27850, n27849, n35212, n27848, n34987, n34715, 
        n43244, n10_adj_4377, n10_adj_4378, n43247, n15414, n35200, 
        n16631, n30861, n16537, n15957, n12_adj_4379, n81, n16869, 
        n34831, n35131, n31006, n15983, n13, Kp_23__N_1535, n31386, 
        n34849, n15942, n34775, n36773, n35051, n34855, n14_adj_4380, 
        n10_adj_4381, n35091, n16570, n43238, n43241, n43232, n35029, 
        n35190, n10_adj_4382, n30549, n43235, n43226, n30562, n35196, 
        n16188, n35251, n43229, n43220, n43223, n35032, n43202, 
        n43205, n43196, n43184, n37031, n34852, n14247, n43187, 
        n35038, Kp_23__N_1783, n10_adj_4383, n34848, n34871, n16610, 
        n10_adj_4384, n35003, n16096, n30974, n14_adj_4385, n43178, 
        n35230, n7_adj_4386, n35094, n31094, Kp_23__N_1189, n14_adj_4387, 
        n10_adj_4388, n37090, n16160, n35069, n34874, n35137, n31030, 
        n16414, n30843, n35048, n35375, n34683, n35016, n34984, 
        n15_adj_4389, n4_adj_4390, n14_adj_4391, n30543, n36905, n31283, 
        n35245, n10_adj_4392, n16252, n16064, n35060, n43181, n34974, 
        n12_adj_4393, n15970, n35173, Kp_23__N_760, n35185, n16892, 
        n16_adj_4394, n30481, n17_adj_4395, n30426, Kp_23__N_1276, 
        n36240, n48, n46, n47, n45_adj_4396, n35248, n44_adj_4397, 
        n43_adj_4398, n54, n49_adj_4399, n35269, n15950, n35209, 
        n35108, n34796, n35260, n36645, n35160, n14_adj_4400, n35115, 
        n15_adj_4401, n10_adj_4402, n34, n14_adj_4404, n10_adj_4405, 
        n35105, n35266, n35122, n28_adj_4406, n19_adj_4407, n38238, 
        n40641, n5_adj_4408, n38239, n38189, n38191, n26_adj_4409, 
        n19_adj_4410, n40636, n5_adj_4411, n38235, n27_adj_4412, n38236, 
        n38219, n14136, n25_adj_4413, n36911, n38221, n34877, n48_adj_4414, 
        n38220, n46_adj_4415, n35167, n35045, n47_adj_4416, n19_adj_4417, 
        n40627, n5_adj_4418, n38232, n38233, n38216, n34867, n45_adj_4419, 
        n35242, n44_adj_4420, n16178, n43_adj_4421, n38218, n54_adj_4422, 
        n38217, n49_adj_4423, n19_adj_4424, n6_adj_4425, n5_adj_4426, 
        n38229, n38230, n38213, n38215, n38214, n19_adj_4427, n6_adj_4428, 
        n5_adj_4429, n38226, n38227, n38210, n38212, n38211, n19_adj_4430, 
        n38223, n6_adj_4431, n5_adj_4432, n38224, n38207, n14_adj_4433, 
        n38209, n40613, n5_adj_4434, Kp_23__N_1183, n38204, n38206, 
        n43172, n43175, n35134, n6_adj_4435, n34969, n6_adj_4436, 
        n37203, n35855, n10_adj_4437, n16354, n10_adj_4438, n30625, 
        n34981, n6_adj_4439, n8_adj_4440, Kp_23__N_731, n6_adj_4441, 
        n34952, n16273, n16503, n16_adj_4442, n31275, n34845, n4_adj_4443, 
        n12_adj_4444, n6_adj_4445, n1, n28_adj_4446, n26_adj_4447, 
        n34997, n34793, n35164, n34934, n16889, n16482, n6_adj_4448, 
        n16312, n34930, n34834, n34911, n6_adj_4449, n16072, n35203, 
        n12_adj_4450, n16229, n16499, n6_adj_4451, n16124, n16020, 
        n35236, n35239, n16376, n16404, n10_adj_4452, n34937, n35151, 
        n1336, n5_adj_4453, n14_adj_4454, n1_adj_4455, n6_adj_4456, 
        n35078, n34809, n35097, n31342, n35035, n35193, n31340, 
        n35224, n34966, n16060, n34824, n6_adj_4457, n36635, n6_adj_4458, 
        n34755, n35072, n34886, n6_adj_4459, n35075, n35176, n30432, 
        n14_adj_4460, n7_adj_4461, n37156, n16593, n18_adj_4462, n6_adj_4463, 
        n27_adj_4464, n25_adj_4465, n16_adj_4466, n34782, n1765, n8_adj_4467, 
        n36296, n20_adj_4468, n6_adj_4469, n35019, n30889, n35088, 
        n16130, n16753, n16857, n12_adj_4470, n16736, n31427, n15974, 
        n28_adj_4471, n34924, n35148, n10_adj_4472, n16370, n16401, 
        n35257, n16886, n26_adj_4473, n27_adj_4474, n16839, n16699, 
        n16417, n16212, n34921, n35145, n10_adj_4475, n25_adj_4476, 
        n6_adj_4477, n12_adj_4478, n31322, n34903, n10_adj_4479, n30994, 
        n34812, n16_adj_4480, n35188, n35254, n17_adj_4481, n30859, 
        n8_adj_4482, n16791, n34759, n34762, n35157, n10_adj_4483, 
        n35118, n36985, n30424, n11, n1558, n16875, n14_adj_4484, 
        n18_adj_4485, n15_adj_4486, n35042, n16324, n19_adj_4487, 
        n16_adj_4488, n35206, n17_adj_4489, n35154, n12_adj_4490, 
        n10_adj_4491, n19260, n42402, n31421, n12_adj_4492, n36936, 
        n10_adj_4493, n34821, n16530, n14_adj_4494, n12_adj_4495, 
        n16713, n15_adj_4496, n16634, n16851, n15_adj_4497, n35009, 
        n6_adj_4498, n16526, n12_adj_4499, n8_adj_4500, n37062, n43807, 
        n10_adj_4501, n37063, n14_adj_4502, n4_adj_4503, n13_adj_4504, 
        n34768, n6_adj_4505, n42_adj_4506, n60, n31302, n34815, 
        n58, n4_adj_4507, n68, n64, n16276, n62, n36809, n34842, 
        n63_adj_4508, n34803, n61, n15886, n66, n72, n38096, n36304, 
        n22, n16016, n65, n73, n38120, n36959, n9_adj_4509, n35263, 
        n35215, n14_adj_4510, n36997, n18_adj_4511, n13_adj_4512, 
        n20_adj_4513, n32_adj_4514, n31_adj_4515, n35, n38098, n30, 
        n25_adj_4516, n34_adj_4517, n38_adj_4518, n6_adj_4519, n33, 
        n8_adj_4520, n6_adj_4521, n16103, n12_adj_4522, n16_adj_4523, 
        n18_adj_4524, n17_adj_4525, n37123, n7_adj_4526, n35111, n35218, 
        n16794, n6_adj_4527, n43166, n43169;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n17900));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n17899));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n17898));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n17897));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n17896));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n17895));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n17894));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n17893));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n17892));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n17891));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n17890));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n17889));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n17888));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17790));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3_c));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n17887));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n17886));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n17885));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n17884));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17789));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n17883));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_21 (.CI(n27809), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27810));
    SB_LUT4 add_44_20_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27808), .O(n2_adj_4257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_20 (.CI(n27808), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27809));
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17804));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17803));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17802));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17801));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17800));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17799));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n17798));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17797));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17796));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n34179));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n34135));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n18046));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n18047));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n17844));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n34037));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n34001));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
           .D(n18093));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
           .D(n18094));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), .C(clk32MHz), 
           .D(n34177));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n17843));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n17842));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n17841));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n18057));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n18058));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n18059));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n18060));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n18048));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n18049));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n18050));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n18051));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n18052));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n18053));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n18054));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n18055));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n18056));   // verilog/coms.v(126[12] 292[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n43329));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n18042));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n18043));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n18044));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n18045));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n18040));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n18041));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n18038));   // verilog/coms.v(126[12] 292[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n18039));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n17960));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n17961));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i194 (.Q(\data_in_frame[24] [1]), .C(clk32MHz), 
           .D(n17936));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i195 (.Q(\data_in_frame[24] [2]), .C(clk32MHz), 
           .D(n17937));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i196 (.Q(\data_in_frame[24] [3]), .C(clk32MHz), 
           .D(n17938));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i197 (.Q(\data_in_frame[24] [4]), .C(clk32MHz), 
           .D(n17939));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i198 (.Q(\data_in_frame[24] [5]), .C(clk32MHz), 
           .D(n17940));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i199 (.Q(\data_in_frame[24] [6]), .C(clk32MHz), 
           .D(n17941));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i200 (.Q(\data_in_frame[24] [7]), .C(clk32MHz), 
           .D(n17942));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i186 (.Q(\data_in_frame[23] [1]), .C(clk32MHz), 
           .D(n17928));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i187 (.Q(\data_in_frame[23] [2]), .C(clk32MHz), 
           .D(n17929));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i188 (.Q(\data_in_frame[23] [3]), .C(clk32MHz), 
           .D(n17930));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i189 (.Q(\data_in_frame[23] [4]), .C(clk32MHz), 
           .D(n17931));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i190 (.Q(\data_in_frame[23] [5]), .C(clk32MHz), 
           .D(n17932));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i191 (.Q(\data_in_frame[23] [6]), .C(clk32MHz), 
           .D(n17933));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n17917));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n17918));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17795));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n17962));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n17963));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n17964));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n17965));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17788));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17787));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n17901));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n17902));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n17903));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n17956));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n17957));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n17958));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n17959));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17786));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17785));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17784));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n17954));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n17955));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n17952));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n17953));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n17950));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n17951));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n17948));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n17949));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n17946));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n17947));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17783));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n17943));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n17944));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n17945));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i192 (.Q(\data_in_frame[23] [7]), .C(clk32MHz), 
           .D(n17934));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i193 (.Q(\data_in_frame[24] [0]), .C(clk32MHz), 
           .D(n17935));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i177 (.Q(\data_in_frame[22] [0]), .C(clk32MHz), 
           .D(n17919));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i178 (.Q(\data_in_frame[22] [1]), .C(clk32MHz), 
           .D(n17920));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i179 (.Q(\data_in_frame[22] [2]), .C(clk32MHz), 
           .D(n17921));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i180 (.Q(\data_in_frame[22] [3]), .C(clk32MHz), 
           .D(n17922));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i181 (.Q(\data_in_frame[22] [4]), .C(clk32MHz), 
           .D(n17923));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i182 (.Q(\data_in_frame[22] [5]), .C(clk32MHz), 
           .D(n17924));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i183 (.Q(\data_in_frame[22] [6]), .C(clk32MHz), 
           .D(n17925));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i184 (.Q(\data_in_frame[22] [7]), .C(clk32MHz), 
           .D(n17926));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i185 (.Q(\data_in_frame[23] [0]), .C(clk32MHz), 
           .D(n17927));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17782));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n17840));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n17839));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n17838));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n17837));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n17836));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17781));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17780));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n17915));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n17916));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n17913));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n17914));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n17911));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n17912));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n17909));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n17910));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n17907));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n17908));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n17904));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n17905));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n17906));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17779));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17778));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17777));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17776));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17775));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17774));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17773));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17772));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17771));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17770));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n17856));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n17835));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n17834));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17769));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17794));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17768));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17793));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17767));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17766));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17792));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17765));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n17833));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17764));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17763));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17762));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_19_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27807), .O(n2_adj_4258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i19954_4_lut (.I0(n24676), .I1(\FRAME_MATCHER.state [0]), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n34704), .O(n24683));   // verilog/coms.v(110[11:16])
    defparam i19954_4_lut.LUT_INIT = 16'hfaea;
    SB_LUT4 i34357_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(tx_transmit_N_3479), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(n23565), .O(n40143));   // verilog/coms.v(110[11:16])
    defparam i34357_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i14794_4_lut (.I0(n24684), .I1(n40143), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n3295[0]));   // verilog/coms.v(110[11:16])
    defparam i14794_4_lut.LUT_INIT = 16'hc5c0;
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n17882));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_3_lut (.I0(\data_out_frame[5] [0]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40568));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13038_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n17767));
    defparam i13038_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31371_4_lut (.I0(n5_c), .I1(\byte_transmit_counter[0] ), .I2(n40044), 
            .I3(n40568), .O(n38201));
    defparam i31371_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31373_4_lut (.I0(n38201), .I1(n43199), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38203));
    defparam i31373_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_44_19 (.CI(n27807), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27808));
    SB_LUT4 i13039_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n17768));
    defparam i13039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13040_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n17769));
    defparam i13040_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_18_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27806), .O(n2_adj_4259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2]_c [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [6]), .O(n38));
    defparam i14_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31346_4_lut (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[2] [7]), .O(n38112));
    defparam i31346_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31348_4_lut (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[0] [3]), .O(n38114));
    defparam i31348_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2][2] ), .I3(\data_in_frame[0] [5]), .O(n39));
    defparam i15_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i19_4_lut (.I0(n25), .I1(n38), .I2(\data_in_frame[0] [4]), 
            .I3(\data_in_frame[1] [3]), .O(n43));
    defparam i19_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i13041_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n17770));
    defparam i13041_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31355_4_lut (.I0(n38112), .I1(\data_in_frame[0] [0]), .I2(n9), 
            .I3(\data_in_frame[2] [6]), .O(n38122));
    defparam i31355_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n38122), .I1(n43), .I2(n39), .I3(n38114), 
            .O(\FRAME_MATCHER.state_31__N_2725 [3]));
    defparam i23_4_lut.LUT_INIT = 16'h0040;
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2][2] ), .C(clk32MHz), 
           .D(n17761));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13042_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n17771));
    defparam i13042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2]_c [1]), .C(clk32MHz), 
           .D(n17760));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2][0] ), .C(clk32MHz), 
           .D(n17759));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n17881));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17758));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17757));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17756));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17755));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17754));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17753));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17752));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17751));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17750));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17749));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17748));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17747));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17746));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n17832));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17745));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17744));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n17743));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n17742));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n17741));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n17740));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n17739));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n17738));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n17831));   // verilog/coms.v(126[12] 292[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n17737));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17736));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13043_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n17772));
    defparam i13043_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17735));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n17830));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13044_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n17773));
    defparam i13044_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13045_3_lut_4_lut (.I0(n8), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n17774));
    defparam i13045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17734));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_4_lut (.I0(n13355), .I1(n31), .I2(n31_adj_4260), .I3(\FRAME_MATCHER.state[1] ), 
            .O(n29));   // verilog/coms.v(110[11:16])
    defparam i1_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35082));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[1] [3]), .I1(n34943), .I2(\data_in_frame[3] [5]), 
            .I3(\data_in_frame[5] [7]), .O(n16448));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSR tx_transmit_3490 (.Q(r_SM_Main_2__N_3582[0]), .C(clk32MHz), 
            .D(n3295[0]), .R(n24683));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34694));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'hbbbb;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3491  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17733));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17732));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n17880));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i3_4_lut_adj_1006 (.I0(\FRAME_MATCHER.state[1] ), .I1(n34694), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n24676), .O(n15876));
    defparam i3_4_lut_adj_1006.LUT_INIT = 16'hffdf;
    SB_LUT4 i18858_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3582[0]), .I2(GND_net), 
            .I3(GND_net), .O(n23565));
    defparam i18858_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18906_2_lut (.I0(n15876), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n23620));
    defparam i18906_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17731));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17730));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17729));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17728));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n17879));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n17878));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n17877));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17727));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17726));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17725));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17724));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17723));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17722));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17721));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17720));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17719));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17718));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n17829));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17717));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n17845));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n17828));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n17855));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17716));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n17876));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18]_c [2]), .C(clk32MHz), 
           .D(n17715));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_18 (.CI(n27806), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27807));
    SB_LUT4 add_44_17_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27805), .O(n2_adj_4261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1007 (.I0(\data_in_frame[4] [1]), .I1(n35063), 
            .I2(\data_in_frame[2][0] ), .I3(\data_in_frame[1] [5]), .O(n16033));   // verilog/coms.v(228[9:81])
    defparam i3_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18][1] ), .C(clk32MHz), 
           .D(n17714));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18][0] ), .C(clk32MHz), 
           .D(n17713));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17712));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_17 (.CI(n27805), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27806));
    SB_LUT4 add_44_16_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27804), .O(n2_adj_4262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13128_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n17857));
    defparam i13128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13129_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n17858));
    defparam i13129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_16 (.CI(n27804), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27805));
    SB_LUT4 add_44_15_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27803), .O(n2_adj_4264)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_15 (.CI(n27803), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27804));
    SB_LUT4 i13130_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n17859));
    defparam i13130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13131_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n17860));
    defparam i13131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17711));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_14_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27802), .O(n2_adj_4265)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17710));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13132_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n17861));
    defparam i13132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_14 (.CI(n27802), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27803));
    SB_LUT4 i13133_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n17862));
    defparam i13133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13126_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n17855));
    defparam i13126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n17854));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13127_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n17856));
    defparam i13127_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n17853));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_13_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27801), .O(n2_adj_4266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_13 (.CI(n27801), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27802));
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n17852));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17709));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i9_3_lut (.I0(\FRAME_MATCHER.state [15]), .I1(\FRAME_MATCHER.state [26]), 
            .I2(\FRAME_MATCHER.state [13]), .I3(GND_net), .O(n26));   // verilog/coms.v(126[12] 292[6])
    defparam i9_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n17851));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n17850));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17708));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17707));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_33_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27821), .O(n2_adj_4267)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_32_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27820), .O(n2_adj_4268)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1008 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [6]), .O(n34961));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_CARRY add_44_32 (.CI(n27820), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27821));
    SB_LUT4 add_44_31_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27819), .O(n2_adj_4269)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[4] [5]), .I1(n16427), .I2(n4_c), 
            .I3(GND_net), .O(n16716));   // verilog/coms.v(228[9:81])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(\data_in_frame[1] [7]), .I1(n34864), 
            .I2(\data_in_frame[2]_c [1]), .I3(GND_net), .O(n16706));   // verilog/coms.v(228[9:81])
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\data_in_frame[4] [4]), .I1(n34749), 
            .I2(GND_net), .I3(GND_net), .O(n16666));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\data_in_frame[1] [4]), .I1(n34961), 
            .I2(GND_net), .I3(GND_net), .O(n16663));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(n34900), .I1(n34978), .I2(GND_net), 
            .I3(GND_net), .O(n31329));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1013 (.I0(n16292), .I1(n31129), .I2(\data_in_frame[5] [1]), 
            .I3(GND_net), .O(n31392));
    defparam i2_3_lut_adj_1013.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(n6), .O(n16053));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1014 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n34806));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1014.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[1] [4]), .I1(n34806), 
            .I2(GND_net), .I3(GND_net), .O(n34786));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1016 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n16427));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_adj_1016.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1017 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(163[9:87])
    defparam i2_3_lut_adj_1017.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n34943));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n34800));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35227));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17706));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17705));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n17849));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17704));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_12_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27800), .O(n2_adj_4270)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_31 (.CI(n27819), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27820));
    SB_LUT4 add_44_30_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27818), .O(n2_adj_4271)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_30 (.CI(n27818), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27819));
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17703));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17702));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17701));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_29_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27817), .O(n2_adj_4272)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_12 (.CI(n27800), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27801));
    SB_CARRY add_44_29 (.CI(n27817), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27818));
    SB_LUT4 add_44_11_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27799), .O(n2_adj_4273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17700));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_11 (.CI(n27799), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27800));
    SB_LUT4 add_44_10_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27798), .O(n2_adj_4274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1021 (.I0(\data_in_frame[2]_c [1]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[2][0] ), .I3(GND_net), .O(n34765));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17699));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17698));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17697));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17696));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17695));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17694));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17693));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17692));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17691));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17690));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17689));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17688));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n17848));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17687));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17686));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17685));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17684));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17683));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17682));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17681));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17680));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17679));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_28_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27816), .O(n2_adj_4275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17678));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17677));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17676));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17675));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17674));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17673));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17672));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17671));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17670));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17669));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17668));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17667));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17666));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17665));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17664));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17663));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17662));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17661));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17660));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17659));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17658));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34883));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17657));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17656));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17655));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17654));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17653));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17652));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17651));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17650));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17649));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17648));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17647));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17646));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17645));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_28 (.CI(n27816), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27817));
    SB_LUT4 i12_4_lut (.I0(\FRAME_MATCHER.state [12]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(\FRAME_MATCHER.state [9]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n29_adj_4276));   // verilog/coms.v(126[12] 292[6])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17644));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35063));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1024 (.I0(n35063), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(\data_in_frame[0] [2]), .O(n36028));   // verilog/coms.v(94[12:25])
    defparam i3_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n34883), .I1(n34765), .I2(n35227), .I3(n36028), 
            .O(n16));   // verilog/coms.v(71[16:34])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n34800), .I1(n34943), .I2(n16430), .I3(n34880), 
            .O(n17));   // verilog/coms.v(71[16:34])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n34786), .I2(n16), .I3(\data_in_frame[2] [7]), 
            .O(n31129));   // verilog/coms.v(71[16:34])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17643));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17642));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17641));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17640));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17639));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17638));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17637));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17636));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17635));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17634));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17633));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17632));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17631));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17630));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17629));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_27_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27815), .O(n2_adj_4277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17628));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17627));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17626));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17625));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_27 (.CI(n27815), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27816));
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17624));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17623));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17622));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17621));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17620));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17619));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17618));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17617));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17616));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17615));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17614));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17613));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17612));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17611));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17610));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17609));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17608));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17607));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17606));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17605));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17604));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17603));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17602));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17601));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17600));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17599));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17598));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_10 (.CI(n27798), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27799));
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17597));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_9_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27797), .O(n2_adj_4278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17596));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17595));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17594));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17593));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17592));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17591));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17590));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17589));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17588));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17587));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17586));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17585));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_9 (.CI(n27797), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27798));
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n17584));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n17583));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n17582));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n17581));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n17580));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_8_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27796), .O(n2_adj_4279)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17579));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n17578));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n17577));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n17576));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n17575));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n17574));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n17573));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_26_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27814), .O(n2_adj_4280)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_26 (.CI(n27814), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27815));
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n17572));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i2_4_lut (.I0(n13355), .I1(n5_adj_4281), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state[1] ), .O(n30070));
    defparam i2_4_lut.LUT_INIT = 16'hffef;
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n17571));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n17570));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17569));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17568));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17567));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_8 (.CI(n27796), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27797));
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17566));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17565));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17564));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17563));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n17562));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n17561));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n17560));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n17559));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n17558));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n17557));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_7_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27795), .O(n2_adj_4282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n17556));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n17555));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17554));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17553));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17552));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17551));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17550));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17549));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17548));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n17547));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4348), .I3(GND_net), .O(n4351));
    defparam mux_1055_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n17546));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n17545));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n17544));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n17543));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n17542));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4348), .I3(GND_net), .O(n4350));
    defparam mux_1055_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13086_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n17815));
    defparam i13086_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n17541));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n17540));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n17539));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13087_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n17816));
    defparam i13087_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n17538));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n17537));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n17536));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n17535));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4348), .I3(GND_net), .O(n4353));
    defparam mux_1055_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n17534));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n17533));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4348), .I3(GND_net), .O(n4352));
    defparam mux_1055_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n17532));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n17531));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n17530));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n17529));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13088_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n17817));
    defparam i13088_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13089_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n17818));
    defparam i13089_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n17528));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n17527));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2][0] ), 
            .I2(n4348), .I3(GND_net), .O(n4357));
    defparam mux_1055_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n17526));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n17525));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17523));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17522));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4348), .I3(GND_net), .O(n4356));
    defparam mux_1055_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1055_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4348), .I3(GND_net), .O(n4355));
    defparam mux_1055_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1055_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4348), .I3(GND_net), .O(n4354));
    defparam mux_1055_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13090_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n17819));
    defparam i13090_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17521));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13091_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n17820));
    defparam i13091_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17520));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17519));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i19012_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_4284), .I3(\FRAME_MATCHER.i [1]), .O(n788));   // verilog/coms.v(154[9:60])
    defparam i19012_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i8_4_lut (.I0(n15839), .I1(\data_in[1] [3]), .I2(n15645), 
            .I3(\data_in[2] [0]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1025 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_1025.LUT_INIT = 16'hfeff;
    SB_LUT4 i13092_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n17821));
    defparam i13092_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17518));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17517));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17516));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17515));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i31342_4_lut (.I0(\data_in[0] [5]), .I1(\data_in[2] [5]), .I2(\data_in[1] [2]), 
            .I3(\data_in[3] [2]), .O(n38108));
    defparam i31342_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n38108), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n63_adj_4285));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1026 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14));
    defparam i6_4_lut_adj_1026.LUT_INIT = 16'hfeff;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17514));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17513));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17512));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i7_4_lut_adj_1027 (.I0(\data_in[3] [6]), .I1(n14), .I2(n10), 
            .I3(\data_in[2] [1]), .O(n15839));
    defparam i7_4_lut_adj_1027.LUT_INIT = 16'hfffd;
    SB_LUT4 i6_4_lut_adj_1028 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4286));
    defparam i6_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1029 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4287));
    defparam i7_4_lut_adj_1029.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1030 (.I0(n17_adj_4287), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4286), .I3(\data_in[3] [7]), .O(n15728));
    defparam i9_4_lut_adj_1030.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1031 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4288));
    defparam i4_4_lut_adj_1031.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut (.I0(\data_in[3] [4]), .I1(n10_adj_4288), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n15741));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17511));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i5_3_lut_adj_1032 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4289));
    defparam i5_3_lut_adj_1032.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1033 (.I0(\data_in[0] [6]), .I1(n15741), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15));
    defparam i6_4_lut_adj_1033.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1034 (.I0(n15), .I1(\data_in[2] [2]), .I2(n14_adj_4289), 
            .I3(\data_in[3] [0]), .O(n15645));
    defparam i8_4_lut_adj_1034.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1035 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n15645), .O(n16_adj_4290));
    defparam i6_4_lut_adj_1035.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1036 (.I0(n15728), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4291));
    defparam i7_4_lut_adj_1036.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1037 (.I0(n17_adj_4291), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4290), .I3(\data_in[3] [3]), .O(n63_adj_4292));
    defparam i9_4_lut_adj_1037.LUT_INIT = 16'hfbff;
    SB_LUT4 i13093_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n17822));
    defparam i13093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17510));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17509));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17508));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n34948), .I1(n10_adj_4293), .I2(n1713), 
            .I3(n31414), .O(n35100));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1038 (.I0(\data_in[2] [4]), .I1(n15839), .I2(\data_in[1] [5]), 
            .I3(n15741), .O(n18));
    defparam i7_4_lut_adj_1038.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1039 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n15728), .O(n20_adj_4294));
    defparam i9_4_lut_adj_1039.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4295));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4295), .I1(n20_adj_4294), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_4296));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4296), 
            .I2(n63_adj_4292), .I3(GND_net), .O(n122));   // verilog/coms.v(110[11:16])
    defparam i1_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i4349_2_lut (.I0(n63_adj_4285), .I1(n788), .I2(GND_net), .I3(GND_net), 
            .O(n9001));   // verilog/coms.v(154[6] 156[9])
    defparam i4349_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(\FRAME_MATCHER.state[1] ), .I1(n34675), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2621 ));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_adj_1041 (.I0(n34948), .I1(n10_adj_4293), .I2(n1713), 
            .I3(n16815), .O(n31306));
    defparam i1_2_lut_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1042 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n15731), .I3(GND_net), .O(n15648));
    defparam i2_3_lut_adj_1042.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[9] [2]), .O(n34948));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17507));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4297));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1043 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_1043.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n16742));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_1044 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4298));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43_adj_4297), .I2(n42), .I3(n44), 
            .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1045 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39_adj_4298), .I3(n40), 
            .O(n15731));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17506));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i2_4_lut_adj_1046 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n7_c), .I3(\FRAME_MATCHER.i [3]), .O(n37049));
    defparam i2_4_lut_adj_1046.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_3_lut_adj_1047 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n16299));
    defparam i1_2_lut_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i19019_3_lut (.I0(n37049), .I1(\FRAME_MATCHER.i [31]), .I2(n15731), 
            .I3(GND_net), .O(n3894));   // verilog/coms.v(248[9:58])
    defparam i19019_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i19005_2_lut (.I0(\byte_transmit_counter[1] ), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n40044));
    defparam i19005_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36253_4_lut (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter[5]), .I3(n24610), .O(tx_transmit_N_3479));
    defparam i36253_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1048 (.I0(\data_out_frame[16] [4]), .I1(n30545), 
            .I2(n35233), .I3(GND_net), .O(n12));
    defparam i1_2_lut_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34704));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17505));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[16] [4]), .I1(n30545), .I2(\data_out_frame[14] [5]), 
            .I3(n31414), .O(n31381));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1050 (.I0(n23620), .I1(n34704), .I2(n2060), .I3(n19504), 
            .O(n2774));
    defparam i2_4_lut_adj_1050.LUT_INIT = 16'h0a02;
    SB_LUT4 i2_3_lut_4_lut_adj_1051 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[15] [5]), .I3(n30491), .O(n31281));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1052 (.I0(n2774), .I1(n1211), .I2(n15876), .I3(GND_net), 
            .O(n5));
    defparam i1_3_lut_adj_1052.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_3_lut_adj_1053 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[13] [2]), .I3(GND_net), .O(n34790));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1053.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17504));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17503));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17502));   // verilog/coms.v(126[12] 292[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17501));   // verilog/coms.v(126[12] 292[6])
    SB_DFF byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), .C(clk32MHz), 
           .D(n34173));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1054 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(n34927), .I3(GND_net), .O(n15489));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1055 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n6_adj_4300));
    defparam i1_2_lut_3_lut_adj_1055.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1056 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [1]), .I3(n16760), .O(n34927));
    defparam i2_3_lut_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1057 (.I0(\data_out_frame[13] [2]), .I1(n34940), 
            .I2(n16029), .I3(\data_out_frame[17] [5]), .O(n34991));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 equal_107_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_c));   // verilog/coms.v(151[7:23])
    defparam equal_107_i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1058 (.I0(\data_out_frame[13] [2]), .I1(n34940), 
            .I2(n34771), .I3(GND_net), .O(n16660));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1058.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1059 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(n31414), .I3(GND_net), .O(n31435));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1059.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(\data_out_frame[16] [3]), .I3(n10_adj_4301), .O(n36954));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1060 (.I0(\data_out_frame[15] [7]), .I1(n35025), 
            .I2(n15422), .I3(\data_out_frame[18] [3]), .O(n35142));
    defparam i1_2_lut_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1061 (.I0(\data_out_frame[15] [7]), .I1(n35025), 
            .I2(n15422), .I3(\data_out_frame[17] [7]), .O(n6_adj_4302));
    defparam i1_2_lut_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1062 (.I0(n31390), .I1(\data_out_frame[20] [1]), 
            .I2(n35057), .I3(GND_net), .O(n35058));
    defparam i1_2_lut_3_lut_adj_1062.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1063 (.I0(n31390), .I1(\data_out_frame[20] [1]), 
            .I2(n34994), .I3(GND_net), .O(n34995));
    defparam i1_2_lut_3_lut_adj_1063.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[4] [7]), .I1(n31394), .I2(\data_in_frame[7] [2]), 
            .I3(GND_net), .O(n35221));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut_adj_1064 (.I0(\data_in_frame[4] [7]), .I1(n31394), 
            .I2(\data_in_frame[6] [6]), .I3(GND_net), .O(n10_adj_4303));
    defparam i2_2_lut_3_lut_adj_1064.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1065 (.I0(\data_in_frame[4] [7]), .I1(n31394), 
            .I2(n31392), .I3(n15426), .O(n35781));
    defparam i2_3_lut_4_lut_adj_1065.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1066 (.I0(\data_in_frame[4] [7]), .I1(n31394), 
            .I2(n34906), .I3(GND_net), .O(n10_adj_4304));
    defparam i2_2_lut_3_lut_adj_1066.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1067 (.I0(n92[1]), .I1(n63_adj_4285), .I2(n34681), 
            .I3(GND_net), .O(n29937));   // verilog/coms.v(141[4] 143[7])
    defparam i1_2_lut_3_lut_adj_1067.LUT_INIT = 16'hb0b0;
    SB_LUT4 i1_2_lut_3_lut_adj_1068 (.I0(n92[1]), .I1(n63_adj_4285), .I2(n5), 
            .I3(GND_net), .O(n34051));   // verilog/coms.v(141[4] 143[7])
    defparam i1_2_lut_3_lut_adj_1068.LUT_INIT = 16'hb0b0;
    SB_LUT4 i19042_2_lut_3_lut (.I0(n63_adj_4296), .I1(n63_adj_4292), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(138[7:80])
    defparam i19042_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1069 (.I0(n63_adj_4296), .I1(n63_adj_4292), 
            .I2(n63_adj_4285), .I3(GND_net), .O(n10337));   // verilog/coms.v(138[7:80])
    defparam i1_2_lut_3_lut_adj_1069.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1070 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n34065));
    defparam i1_2_lut_3_lut_adj_1070.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1071 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n34105));
    defparam i1_2_lut_3_lut_adj_1071.LUT_INIT = 16'he0e0;
    SB_LUT4 add_44_25_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27813), .O(n2_adj_4306)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_25 (.CI(n27813), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27814));
    SB_LUT4 add_44_24_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27812), .O(n2_adj_4307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_22 (.CI(n27810), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27811));
    SB_CARRY add_44_7 (.CI(n27795), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27796));
    SB_LUT4 add_44_6_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27794), .O(n2_adj_4308)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_1055_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4348), .I3(GND_net), .O(n4368));
    defparam mux_1055_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1072 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n34107));
    defparam i1_2_lut_3_lut_adj_1072.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1055_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4348), .I3(GND_net), .O(n4367));
    defparam mux_1055_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4309), .S(n3_adj_4310));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n17827));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i5_4_lut (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n12_adj_4311));   // verilog/coms.v(126[12] 292[6])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [8]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n28));   // verilog/coms.v(126[12] 292[6])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1073 (.I0(n29_adj_4276), .I1(\FRAME_MATCHER.state [14]), 
            .I2(n26), .I3(\FRAME_MATCHER.state [29]), .O(n32));   // verilog/coms.v(126[12] 292[6])
    defparam i15_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1074 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n34063));
    defparam i1_2_lut_3_lut_adj_1074.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1075 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n34069));
    defparam i1_2_lut_3_lut_adj_1075.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1055_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4348), .I3(GND_net), .O(n4366));
    defparam mux_1055_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1076 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n34129));
    defparam i1_2_lut_3_lut_adj_1076.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17806));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4348), .I3(GND_net), .O(n4365));
    defparam mux_1055_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_44_6 (.CI(n27794), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27795));
    SB_LUT4 add_44_23_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27811), .O(n2_adj_4312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_23 (.CI(n27811), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27812));
    SB_LUT4 add_44_5_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27793), .O(n2_adj_4313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1077 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n34109));
    defparam i1_2_lut_3_lut_adj_1077.LUT_INIT = 16'he0e0;
    SB_CARRY add_44_5 (.CI(n27793), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27794));
    SB_LUT4 add_44_4_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27792), .O(n2_adj_4314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_22_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27810), .O(n2_adj_4315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_4 (.CI(n27792), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27793));
    SB_LUT4 i1_2_lut_3_lut_adj_1078 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n34111));
    defparam i1_2_lut_3_lut_adj_1078.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n17826));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n17825));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 add_44_3_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27791), .O(n2_adj_4309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n17824));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n17823));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n17822));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4314), .S(n3_adj_4316));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i19585_2_lut_3_lut (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n24311));
    defparam i19585_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4313), .S(n3_adj_4317));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4308), .S(n3_adj_4318));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4282), .S(n3_adj_4319));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4279), .S(n3_adj_4320));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4278), .S(n3_adj_4321));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4274), .S(n3_adj_4322));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4273), .S(n3_adj_4323));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4270), .S(n3_adj_4324));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4266), .S(n3_adj_4325));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4265), .S(n3_adj_4326));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4264), .S(n3_adj_4327));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4262), .S(n3_adj_4328));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4261), .S(n3_adj_4329));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4259), .S(n3_adj_4330));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4258), .S(n3_adj_4331));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4257), .S(n3_adj_4332));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4333), .S(n3_adj_4334));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4315), .S(n3_adj_4335));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4312), .S(n3_adj_4336));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4307), .S(n3_adj_4337));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4306), .S(n3_adj_4338));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4280), .S(n3_adj_4339));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4277), .S(n3_adj_4340));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4275), .S(n3_adj_4341));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4272), .S(n3_adj_4342));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4271), .S(n3_adj_4343));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4269), .S(n3_adj_4344));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4268), .S(n3_adj_4345));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4267), .S(n3_adj_4346));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n17010), .D(n37121));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4348), .I3(GND_net), .O(n4364));
    defparam mux_1055_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n17010), .D(n36413));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n17010), .D(n36072));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n17010), .D(n36454));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n17010), .D(n36358));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n17010), .D(n36643));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n17010), .D(n36919));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n17010), .D(n37102));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n17010), .D(n34972));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n17010), .D(n35055));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n17010), .D(n34995));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n17010), .D(n35058));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n17010), .D(n34964));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n17010), .D(n35194));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n17010), .D(n34829));   // verilog/coms.v(126[12] 292[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n17010), .D(n37115));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state[1] ), .C(clk32MHz), 
            .D(n34051), .S(n43574));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1079 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n24309));
    defparam i1_2_lut_3_lut_adj_1079.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1080 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n34113));
    defparam i1_2_lut_3_lut_adj_1080.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1081 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n34115));
    defparam i1_2_lut_3_lut_adj_1081.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n34053), .S(n34193));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n23582), .S(n34059));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n34195), .S(n34055));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n34197), .S(n34127));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n34199), .S(n34125));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n34201), .S(n34123));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n34203), .S(n34121));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n23584), .S(n24305));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n34205), .S(n34119));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n23586), .S(n24307));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n34207), .S(n34117));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n34209), .S(n34115));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_4347), .S(n8_adj_4348));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n34211), .S(n34113));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n23588), .S(n24309));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n23590), .S(n24311));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n34213), .S(n34111));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n34215), .S(n34109));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n7_adj_4349), .S(n8_adj_4350));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n34187), .S(n34129));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_4351), .S(n8_adj_4352));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n34221), .S(n34069));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n23592), .S(n34063));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n34217), .S(n34107));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_4353), .S(n8_adj_4354));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n34219), .S(n34105));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n7_adj_4355), .S(n8_adj_4356));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n23594), .S(n34065));   // verilog/coms.v(126[12] 292[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4357), .S(n8_adj_4358));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n17821));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 mux_1055_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4348), .I3(GND_net), .O(n4363));
    defparam mux_1055_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1055_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4348), .I3(GND_net), .O(n4362));
    defparam mux_1055_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1082 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n34117));
    defparam i1_2_lut_3_lut_adj_1082.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1083 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n34119));
    defparam i1_2_lut_3_lut_adj_1083.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1084 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n34121));
    defparam i1_2_lut_3_lut_adj_1084.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1085 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n34123));
    defparam i1_2_lut_3_lut_adj_1085.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1086 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n34125));
    defparam i1_2_lut_3_lut_adj_1086.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1055_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4348), .I3(GND_net), .O(n4361));
    defparam mux_1055_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1055_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4348), .I3(GND_net), .O(n4360));
    defparam mux_1055_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1087 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n34127));
    defparam i1_2_lut_3_lut_adj_1087.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1088 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n34055));
    defparam i1_2_lut_3_lut_adj_1088.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1089 (.I0(n50_adj_4305), .I1(n27214), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n34059));
    defparam i1_2_lut_3_lut_adj_1089.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1090 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [31]), .O(n8_adj_4358));
    defparam i1_2_lut_4_lut_adj_1090.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1091 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [29]), .O(n8_adj_4356));
    defparam i1_2_lut_4_lut_adj_1091.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1092 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [27]), .O(n8_adj_4354));
    defparam i1_2_lut_4_lut_adj_1092.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43298));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17417));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1093 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [23]), .O(n8_adj_4352));
    defparam i1_2_lut_4_lut_adj_1093.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1094 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [21]), .O(n8_adj_4350));
    defparam i1_2_lut_4_lut_adj_1094.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n17820));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1095 (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [15]), .O(n8_adj_4348));
    defparam i1_2_lut_4_lut_adj_1095.LUT_INIT = 16'hfe00;
    SB_LUT4 i19583_2_lut_4_lut (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [12]), .O(n24307));
    defparam i19583_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i19582_2_lut_4_lut (.I0(n49), .I1(n37), .I2(n50_adj_4305), 
            .I3(\FRAME_MATCHER.state [10]), .O(n24305));
    defparam i19582_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1096 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[7] [0]), .I3(GND_net), .O(n16641));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1055_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4348), .I3(GND_net), .O(n4372));
    defparam mux_1055_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1097 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(n34961), .I3(GND_net), .O(n6_adj_4359));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1097.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1055_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4348), .I3(GND_net), .O(n4371));
    defparam mux_1055_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1098 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [4]), .I3(n16382), .O(n35179));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_3_lut (.I0(\data_in_frame[12] [6]), .I1(n34955), .I2(n16382), 
            .I3(GND_net), .O(n14_adj_4360));   // verilog/coms.v(83[17:28])
    defparam i6_4_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1099 (.I0(n16706), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[8] [6]), .I3(n10_adj_4361), .O(n31060));   // verilog/coms.v(72[16:43])
    defparam i5_3_lut_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1100 (.I0(n16706), .I1(\data_in_frame[6] [4]), 
            .I2(n16033), .I3(\data_in_frame[6] [3]), .O(Kp_23__N_1186));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1055_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4348), .I3(GND_net), .O(n4370));
    defparam mux_1055_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_44_24 (.CI(n27812), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27813));
    SB_DFFESR LED_3493 (.Q(LED_c), .C(clk32MHz), .E(n36824), .D(n41_adj_4362), 
            .R(n36660));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i2_3_lut_adj_1101 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n6_adj_4363));   // verilog/coms.v(163[9:87])
    defparam i2_3_lut_adj_1101.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1055_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4348), .I3(GND_net), .O(n4369));
    defparam mux_1055_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13030_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[2][0] ), .O(n17759));
    defparam i13030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13031_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[2]_c [1]), .O(n17760));
    defparam i13031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_3_lut (.I0(n35006), .I1(n35179), .I2(\data_in_frame[13] [7]), 
            .I3(GND_net), .O(n35022));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_2_lut (.I0(n35179), .I1(\data_in_frame[12] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n31439));
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n17819));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n17818));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n17875));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i1_2_lut_adj_1102 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34880));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n17874));   // verilog/coms.v(126[12] 292[6])
    SB_CARRY add_44_3 (.CI(n27791), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27792));
    SB_LUT4 add_44_2_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27791));
    SB_LUT4 i13134_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n17863));
    defparam i13134_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13135_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n17864));
    defparam i13135_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1103 (.I0(\data_in_frame[0] [5]), .I1(n34837), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [7]), .O(n16292));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i13136_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n17865));
    defparam i13136_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13032_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[2][2] ), .O(n17761));
    defparam i13032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13137_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n17866));
    defparam i13137_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n43298_bdd_4_lut (.I0(n43298), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43301));
    defparam n43298_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36445 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43292));
    defparam byte_transmit_counter_0__bdd_4_lut_36445.LUT_INIT = 16'he4aa;
    SB_LUT4 n43292_bdd_4_lut (.I0(n43292), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43295));
    defparam n43292_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36440 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43286));
    defparam byte_transmit_counter_0__bdd_4_lut_36440.LUT_INIT = 16'he4aa;
    SB_LUT4 n43286_bdd_4_lut (.I0(n43286), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43289));
    defparam n43286_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36435 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43280));
    defparam byte_transmit_counter_0__bdd_4_lut_36435.LUT_INIT = 16'he4aa;
    SB_LUT4 n43280_bdd_4_lut (.I0(n43280), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43283));
    defparam n43280_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36430 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43274));
    defparam byte_transmit_counter_0__bdd_4_lut_36430.LUT_INIT = 16'he4aa;
    SB_LUT4 n43274_bdd_4_lut (.I0(n43274), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43277));
    defparam n43274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36425 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43268));
    defparam byte_transmit_counter_0__bdd_4_lut_36425.LUT_INIT = 16'he4aa;
    SB_LUT4 n43268_bdd_4_lut (.I0(n43268), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43271));
    defparam n43268_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36420 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43262));
    defparam byte_transmit_counter_0__bdd_4_lut_36420.LUT_INIT = 16'he4aa;
    SB_LUT4 n43262_bdd_4_lut (.I0(n43262), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43265));
    defparam n43262_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36415 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43256));
    defparam byte_transmit_counter_0__bdd_4_lut_36415.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n17873));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n17872));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n17871));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i18086_3_lut (.I0(\Kp[9] ), .I1(\data_in_frame[2]_c [1]), .I2(n30070), 
            .I3(GND_net), .O(n17556));
    defparam i18086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13033_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n17762));
    defparam i13033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13138_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n17867));
    defparam i13138_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13139_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n17868));
    defparam i13139_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13140_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n17869));
    defparam i13140_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13141_3_lut_4_lut (.I0(n24351), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n17870));
    defparam i13141_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13078_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n17807));
    defparam i13078_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n34067));   // verilog/coms.v(126[12] 292[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17398));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n17870));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13034_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n17763));
    defparam i13034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n17869));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n17868));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n17867));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n17866));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n17817));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n17816));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n17815));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n17814));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n17847));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17397));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13079_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n17808));
    defparam i13079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13080_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n17809));
    defparam i13080_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13081_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n17810));
    defparam i13081_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13082_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n17811));
    defparam i13082_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17396));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 n43256_bdd_4_lut (.I0(n43256), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43259));
    defparam n43256_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13083_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n17812));
    defparam i13083_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n17395));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n17394));   // verilog/coms.v(126[12] 292[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17393));   // verilog/coms.v(126[12] 292[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n17392));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13084_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n17813));
    defparam i13084_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13085_3_lut_4_lut (.I0(n10_adj_4365), .I1(n34697), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n17814));
    defparam i13085_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1104 (.I0(\FRAME_MATCHER.state [18]), .I1(n12_adj_4311), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [20]), 
            .O(n31141));   // verilog/coms.v(126[12] 292[6])
    defparam i6_4_lut_adj_1104.LUT_INIT = 16'hfffe;
    SB_LUT4 i13035_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n17764));
    defparam i13035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34837));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1106 (.I0(\data_in_frame[14] [1]), .I1(n15435), 
            .I2(\data_in_frame[16] [3]), .I3(n30525), .O(n35785));
    defparam i2_3_lut_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1107 (.I0(\data_in_frame[14] [1]), .I1(n15435), 
            .I2(\data_in_frame[16] [2]), .I3(n30999), .O(n31320));
    defparam i2_3_lut_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1108 (.I0(\data_in_frame[15] [7]), .I1(n31310), 
            .I2(\data_in_frame[16] [1]), .I3(n30999), .O(n31273));
    defparam i2_3_lut_4_lut_adj_1108.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1109 (.I0(\data_in_frame[15] [7]), .I1(n31310), 
            .I2(\data_in_frame[18] [0]), .I3(n14249), .O(n6_adj_4366));
    defparam i2_3_lut_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1110 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [10]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n27));   // verilog/coms.v(126[12] 292[6])
    defparam i10_4_lut_adj_1110.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1111 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[13] [4]), 
            .I2(n31368), .I3(GND_net), .O(n6_adj_4367));
    defparam i1_2_lut_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1112 (.I0(n27), .I1(n31141), .I2(n32), .I3(n28), 
            .O(n27212));   // verilog/coms.v(126[12] 292[6])
    defparam i1_4_lut_adj_1112.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1113 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[16] [6]), .I3(GND_net), .O(n35182));
    defparam i1_2_lut_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1114 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [0]), 
            .I2(\data_in_frame[21] [3]), .I3(GND_net), .O(n34746));
    defparam i1_2_lut_3_lut_adj_1114.LUT_INIT = 16'h9696;
    SB_LUT4 i13036_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n17765));
    defparam i13036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1115 (.I0(n35170), .I1(n10_adj_4368), .I2(n31327), 
            .I3(\data_in_frame[17] [7]), .O(n31298));
    defparam i1_2_lut_4_lut_adj_1115.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1116 (.I0(n35170), .I1(n10_adj_4368), .I2(n31327), 
            .I3(\data_in_frame[20] [1]), .O(n34897));
    defparam i1_2_lut_4_lut_adj_1116.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17805));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i31422_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38252));
    defparam i31422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31423_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38253));
    defparam i31423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31426_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38256));
    defparam i31426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31425_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38255));
    defparam i31425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31416_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38246));
    defparam i31416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31417_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38247));
    defparam i31417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31420_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38250));
    defparam i31420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31419_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38249));
    defparam i31419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31410_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38240));
    defparam i31410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31411_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38241));
    defparam i31411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31414_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38244));
    defparam i31414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31413_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38243));
    defparam i31413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14561_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n16_adj_4369));   // verilog/coms.v(100[12:33])
    defparam i14561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18][1] ), 
            .I1(\data_out_frame[19] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4370));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33739_2_lut (.I0(\data_out_frame[22] [1]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n40113));
    defparam i33739_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4371));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n16_adj_4372));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18][0] ), 
            .I1(\data_out_frame[19] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4373));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33745_2_lut (.I0(\data_out_frame[22] [0]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n40133));
    defparam i33745_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4374));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31452_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38282));
    defparam i31452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31453_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38283));
    defparam i31453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31456_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38286));
    defparam i31456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31455_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n38285));
    defparam i31455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13037_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n17766));
    defparam i13037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13022_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n17751));
    defparam i13022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1117 (.I0(\FRAME_MATCHER.state [7]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [4]), 
            .O(n34603));
    defparam i3_4_lut_adj_1117.LUT_INIT = 16'hfffe;
    SB_LUT4 i19948_2_lut (.I0(n34603), .I1(n27212), .I2(GND_net), .I3(GND_net), 
            .O(n24676));
    defparam i19948_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1118 (.I0(n19503), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n34675));
    defparam i2_3_lut_adj_1118.LUT_INIT = 16'h0404;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36410 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n43250));
    defparam byte_transmit_counter_0__bdd_4_lut_36410.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n19503), .O(\FRAME_MATCHER.i_31__N_2625 ));   // verilog/coms.v(126[12] 292[6])
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'h0040;
    SB_LUT4 i13023_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n17752));
    defparam i13023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(150[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_adj_1120 (.I0(\FRAME_MATCHER.i_31__N_2625 ), .I1(n34675), 
            .I2(GND_net), .I3(GND_net), .O(n2060));
    defparam i2_2_lut_adj_1120.LUT_INIT = 16'heeee;
    SB_LUT4 i13024_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n17753));
    defparam i13024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13025_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n17754));
    defparam i13025_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n17813));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n17812));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13026_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n17755));
    defparam i13026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n17811));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n17810));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n17809));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13118_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n17847));
    defparam i13118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13119_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n17848));
    defparam i13119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13120_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n17849));
    defparam i13120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13121_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n17850));
    defparam i13121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13122_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n17851));
    defparam i13122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13123_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n17852));
    defparam i13123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13124_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n17853));
    defparam i13124_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13125_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n17854));
    defparam i13125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_21_lut (.I0(n2060), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27809), .O(n2_adj_4333)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n43250_bdd_4_lut (.I0(n43250), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n43253));
    defparam n43250_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13027_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n17756));
    defparam i13027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n17249));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13028_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n17757));
    defparam i13028_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13117_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n17846));
    defparam i13117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13116_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n17845));
    defparam i13116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17791));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13110_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n17839));
    defparam i13110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13111_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n17840));
    defparam i13111_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13112_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n17841));
    defparam i13112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n17846));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13113_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n17842));
    defparam i13113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n17865));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13029_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n17758));
    defparam i13029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3591_9_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n27854), .O(n40145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3591_8_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n27853), .O(n40179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_8 (.CI(n27853), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n27854));
    SB_LUT4 add_3591_7_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n27852), .O(n40273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_7 (.CI(n27852), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n27853));
    SB_LUT4 i13114_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n17843));
    defparam i13114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3591_6_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n27851), .O(n40274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_6 (.CI(n27851), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n27852));
    SB_LUT4 add_3591_5_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n27850), .O(n40275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_5 (.CI(n27850), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n27851));
    SB_LUT4 i13115_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n17844));
    defparam i13115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3591_4_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n27849), .O(n40278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_4 (.CI(n27849), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n27850));
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35212));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 add_3591_3_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n27848), .O(n40277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_3 (.CI(n27848), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n27849));
    SB_LUT4 add_3591_2_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3479), .I3(GND_net), .O(n40276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3591_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3591_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3479), .CO(n27848));
    SB_LUT4 i1_3_lut_adj_1122 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(n34900), .I3(GND_net), .O(n34987));
    defparam i1_3_lut_adj_1122.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n17864));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n17863));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n17862));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17808));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17807));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n17861));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13173_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n17902));
    defparam i13173_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n17860));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36405 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43244));
    defparam byte_transmit_counter_0__bdd_4_lut_36405.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n17859));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13172_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n17901));
    defparam i13172_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n17858));   // verilog/coms.v(126[12] 292[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n17857));   // verilog/coms.v(126[12] 292[6])
    SB_LUT4 i13166_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n17895));
    defparam i13166_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13167_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n17896));
    defparam i13167_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13168_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n17897));
    defparam i13168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13169_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n17898));
    defparam i13169_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13170_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n17899));
    defparam i13170_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13171_3_lut_4_lut (.I0(n8), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n17900));
    defparam i13171_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1123 (.I0(n2060), .I1(n161), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n7_c), .O(n34697));
    defparam i2_3_lut_4_lut_adj_1123.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(n2060), .I1(n161), .I2(n10_adj_4365), 
            .I3(GND_net), .O(n34723));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(n2060), .I1(n161), .I2(n10_adj_4377), 
            .I3(GND_net), .O(n34707));
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1126 (.I0(n2060), .I1(n161), .I2(n10_adj_4378), 
            .I3(GND_net), .O(n34715));
    defparam i1_2_lut_3_lut_adj_1126.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_4_lut_adj_1127 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n34697), .I3(\FRAME_MATCHER.i [3]), .O(n36887));   // verilog/coms.v(151[7:23])
    defparam i2_3_lut_4_lut_adj_1127.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_112_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4378));   // verilog/coms.v(151[7:23])
    defparam equal_112_i10_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_113_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(151[7:23])
    defparam equal_113_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 equal_122_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4364));   // verilog/coms.v(151[7:23])
    defparam equal_122_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i13158_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n17887));
    defparam i13158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13159_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n17888));
    defparam i13159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13160_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n17889));
    defparam i13160_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13161_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n17890));
    defparam i13161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13162_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n17891));
    defparam i13162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n43244_bdd_4_lut (.I0(n43244), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43247));
    defparam n43244_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13163_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n17892));
    defparam i13163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13164_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n17893));
    defparam i13164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13165_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n17894));
    defparam i13165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14802_3_lut (.I0(byte_transmit_counter_c[7]), .I1(n40145), 
            .I2(n24391), .I3(GND_net), .O(n18094));
    defparam i14802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14769_3_lut (.I0(byte_transmit_counter_c[6]), .I1(n40179), 
            .I2(n24391), .I3(GND_net), .O(n18093));
    defparam i14769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13054_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n17783));
    defparam i13054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13055_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n17784));
    defparam i13055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13056_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n17785));
    defparam i13056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.state_31__I_0_3574_i64_1_lut  (.I0(n15876), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2624 ));   // verilog/coms.v(204[5:16])
    defparam \FRAME_MATCHER.state_31__I_0_3574_i64_1_lut .LUT_INIT = 16'h5555;
    SB_LUT4 i13057_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n17786));
    defparam i13057_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13058_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n17787));
    defparam i13058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1055_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2][2] ), 
            .I2(n4348), .I3(GND_net), .O(n4359));
    defparam mux_1055_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13059_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n17788));
    defparam i13059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13060_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n17789));
    defparam i13060_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13061_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n17790));
    defparam i13061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_104_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4376));   // verilog/coms.v(151[7:23])
    defparam equal_104_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_119_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4375));   // verilog/coms.v(151[7:23])
    defparam equal_119_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_119_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4365));   // verilog/coms.v(151[7:23])
    defparam equal_119_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_125_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4377));   // verilog/coms.v(151[7:23])
    defparam equal_125_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_in_frame[15] [0]), .I1(n15414), 
            .I2(GND_net), .I3(GND_net), .O(n35200));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16631));
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1130 (.I0(n16631), .I1(n30861), .I2(n16537), 
            .I3(n15957), .O(n12_adj_4379));
    defparam i5_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_31_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4346));
    defparam select_343_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_30_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4345));
    defparam select_343_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_29_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4344));
    defparam select_343_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_28_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4343));
    defparam select_343_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_27_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4342));
    defparam select_343_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i6_4_lut_adj_1131 (.I0(n16869), .I1(n12_adj_4379), .I2(n35200), 
            .I3(\data_in_frame[19] [6]), .O(n34831));
    defparam i6_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i14559_3_lut (.I0(\data_out_frame[18]_c [2]), .I1(\displacement[18] ), 
            .I2(n13263), .I3(GND_net), .O(n17715));
    defparam i14559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1132 (.I0(n35131), .I1(n31006), .I2(n31298), 
            .I3(n15983), .O(n13));
    defparam i5_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1133 (.I0(n13), .I1(Kp_23__N_1535), .I2(n6_adj_4366), 
            .I3(n31386), .O(n34849));
    defparam i7_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15942));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1135 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[18] [3]), .I3(n15942), .O(n34775));
    defparam i3_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1136 (.I0(\data_in_frame[17] [4]), .I1(n36773), 
            .I2(GND_net), .I3(GND_net), .O(n15983));
    defparam i1_2_lut_adj_1136.LUT_INIT = 16'h9999;
    SB_LUT4 select_343_Select_26_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4341));
    defparam select_343_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i6_4_lut_adj_1137 (.I0(n35051), .I1(n34855), .I2(n31298), 
            .I3(\data_in_frame[17] [5]), .O(n14_adj_4380));
    defparam i6_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_25_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4340));
    defparam select_343_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i7_4_lut_adj_1138 (.I0(n35131), .I1(n14_adj_4380), .I2(n10_adj_4381), 
            .I3(\data_in_frame[19] [5]), .O(n30861));
    defparam i7_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_24_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4339));
    defparam select_343_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(n31273), .I1(n34775), .I2(GND_net), 
            .I3(GND_net), .O(n35091));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[21] [4]), .I1(\data_in_frame[21] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16570));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36400 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43238));
    defparam byte_transmit_counter_0__bdd_4_lut_36400.LUT_INIT = 16'he4aa;
    SB_LUT4 n43238_bdd_4_lut (.I0(n43238), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43241));
    defparam n43238_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_343_Select_23_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4338));
    defparam select_343_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_22_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4337));
    defparam select_343_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36395 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43232));
    defparam byte_transmit_counter_0__bdd_4_lut_36395.LUT_INIT = 16'he4aa;
    SB_LUT4 select_343_Select_21_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4336));
    defparam select_343_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1141 (.I0(n35029), .I1(n35785), .I2(\data_in_frame[18] [2]), 
            .I3(n35190), .O(n10_adj_4382));
    defparam i4_4_lut_adj_1141.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1142 (.I0(\data_in_frame[20] [5]), .I1(n10_adj_4382), 
            .I2(\data_in_frame[20] [3]), .I3(GND_net), .O(n30549));
    defparam i5_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_LUT4 n43232_bdd_4_lut (.I0(n43232), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43235));
    defparam n43232_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36390 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43226));
    defparam byte_transmit_counter_0__bdd_4_lut_36390.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(n30562), .I1(n35196), .I2(n16570), 
            .I3(n16188), .O(n35251));
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_20_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4335));
    defparam select_343_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 n43226_bdd_4_lut (.I0(n43226), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43229));
    defparam n43226_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_343_Select_19_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4334));
    defparam select_343_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36385 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18]_c [2]), .I2(\data_out_frame[19] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n43220));
    defparam byte_transmit_counter_0__bdd_4_lut_36385.LUT_INIT = 16'he4aa;
    SB_LUT4 n43220_bdd_4_lut (.I0(n43220), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n43223));
    defparam n43220_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35032));
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n38285), .I2(n38286), .I3(byte_transmit_counter[2]), .O(n43202));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43202_bdd_4_lut (.I0(n43202), .I1(n38283), .I2(n38282), .I3(byte_transmit_counter[2]), 
            .O(n43205));
    defparam n43202_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36367 (.I0(\byte_transmit_counter[1] ), 
            .I1(n19_adj_4374), .I2(n40133), .I3(byte_transmit_counter[2]), 
            .O(n43196));
    defparam byte_transmit_counter_1__bdd_4_lut_36367.LUT_INIT = 16'he4aa;
    SB_LUT4 n43196_bdd_4_lut (.I0(n43196), .I1(n17_adj_4373), .I2(n16_adj_4372), 
            .I3(byte_transmit_counter[2]), .O(n43199));
    defparam n43196_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_343_Select_18_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4332));
    defparam select_343_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_17_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4331));
    defparam select_343_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(n31298), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35190));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36362 (.I0(\byte_transmit_counter[1] ), 
            .I1(n19_adj_4371), .I2(n40113), .I3(byte_transmit_counter[2]), 
            .O(n43184));
    defparam byte_transmit_counter_1__bdd_4_lut_36362.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1146 (.I0(n37031), .I1(n35190), .I2(\data_in_frame[20] [2]), 
            .I3(GND_net), .O(n34852));
    defparam i2_3_lut_adj_1146.LUT_INIT = 16'h6969;
    SB_LUT4 select_343_Select_16_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4330));
    defparam select_343_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(n16537), .I1(n36773), .I2(GND_net), 
            .I3(GND_net), .O(n14247));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h9999;
    SB_LUT4 n43184_bdd_4_lut (.I0(n43184), .I1(n17_adj_4370), .I2(n16_adj_4369), 
            .I3(byte_transmit_counter[2]), .O(n43187));
    defparam n43184_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1148 (.I0(\data_in_frame[17] [5]), .I1(n34897), 
            .I2(\data_in_frame[17] [6]), .I3(n16537), .O(n31006));
    defparam i3_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1149 (.I0(\data_in_frame[20] [2]), .I1(n35038), 
            .I2(n31273), .I3(\data_in_frame[20] [3]), .O(Kp_23__N_1783));
    defparam i3_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_15_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4329));
    defparam select_343_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1150 (.I0(\data_in_frame[19] [7]), .I1(n14247), 
            .I2(\data_in_frame[18] [1]), .I3(n34852), .O(n10_adj_4383));
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i12668_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n17397));
    defparam i12668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(n34848), .I1(n34871), .I2(GND_net), 
            .I3(GND_net), .O(n16610));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1152 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4384));
    defparam i2_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1153 (.I0(n35003), .I1(\data_in_frame[12] [7]), 
            .I2(n16096), .I3(n30974), .O(n14_adj_4385));
    defparam i6_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_14_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4328));
    defparam select_343_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i7_4_lut_adj_1154 (.I0(\data_in_frame[15] [3]), .I1(n14_adj_4385), 
            .I2(n10_adj_4384), .I3(\data_in_frame[13] [1]), .O(n36773));
    defparam i7_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36353 (.I0(\byte_transmit_counter[1] ), 
            .I1(n38243), .I2(n38244), .I3(byte_transmit_counter[2]), .O(n43178));
    defparam byte_transmit_counter_1__bdd_4_lut_36353.LUT_INIT = 16'he4aa;
    SB_LUT4 select_343_Select_13_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4327));
    defparam select_343_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1155 (.I0(\data_in_frame[15] [5]), .I1(n35230), 
            .I2(n34955), .I3(\data_in_frame[13] [4]), .O(n10_adj_4368));
    defparam i4_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1156 (.I0(n16292), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[3] [1]), .I3(GND_net), .O(n15426));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1156.LUT_INIT = 16'h9696;
    SB_LUT4 i13015_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n17744));
    defparam i13015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18081_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(\data_in_frame[0] [2]), 
            .I3(rx_data[2]), .O(n17745));
    defparam i18081_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 select_343_Select_12_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4326));
    defparam select_343_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 data_in_frame_19__7__I_0_3516_2_lut (.I0(\data_in_frame[19] [7]), 
            .I1(\data_in_frame[19] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1535));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_19__7__I_0_3516_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_343_Select_11_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4325));
    defparam select_343_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(\data_in_frame[11] [3]), .I1(n31368), 
            .I2(n31060), .I3(GND_net), .O(n31327));
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1158 (.I0(n7_adj_4386), .I1(\data_in_frame[13] [6]), 
            .I2(n31327), .I3(n35094), .O(n14249));
    defparam i4_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35003));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_in_frame[13] [3]), .I1(n31094), 
            .I2(GND_net), .I3(GND_net), .O(n35230));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 select_343_Select_10_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4324));
    defparam select_343_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i13017_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n17746));
    defparam i13017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_343_Select_9_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4323));
    defparam select_343_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_8_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4322));
    defparam select_343_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_7_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4321));
    defparam select_343_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i6_4_lut_adj_1161 (.I0(n35230), .I1(n31060), .I2(n35003), 
            .I3(Kp_23__N_1189), .O(n14_adj_4387));
    defparam i6_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1162 (.I0(\data_in_frame[15] [4]), .I1(n14_adj_4387), 
            .I2(n10_adj_4388), .I3(\data_in_frame[8] [6]), .O(n16537));
    defparam i7_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i13018_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n17747));
    defparam i13018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1163 (.I0(\data_in_frame[17] [6]), .I1(n16537), 
            .I2(\data_in_frame[17] [7]), .I3(GND_net), .O(n34855));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[18] [2]), .I1(n6_adj_4366), .I2(n34855), 
            .I3(GND_net), .O(n37090));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_343_Select_6_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4320));
    defparam select_343_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(n14249), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16160));
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 select_343_Select_5_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4319));
    defparam select_343_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_4_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4318));
    defparam select_343_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_3_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4317));
    defparam select_343_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i3_4_lut_adj_1165 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[18] [7]), .I3(\data_in_frame[19] [1]), .O(n35069));
    defparam i3_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1166 (.I0(n34874), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[11] [2]), .I3(n35137), .O(n10_adj_4361));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 select_343_Select_2_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4316));
    defparam select_343_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_343_Select_1_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4310));
    defparam select_343_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1167 (.I0(\data_in_frame[13] [5]), .I1(n31030), 
            .I2(n31060), .I3(n6_adj_4367), .O(n37031));
    defparam i4_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16414));
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1169 (.I0(\data_in_frame[19] [2]), .I1(n30843), 
            .I2(\data_in_frame[19] [4]), .I3(GND_net), .O(n35048));
    defparam i2_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 select_343_Select_0_i3_2_lut_4_lut (.I0(n19503), .I1(n2060), 
            .I2(n81), .I3(\FRAME_MATCHER.i [0]), .O(n3_c));
    defparam select_343_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i36303_3_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n35375), .O(n36660));   // verilog/coms.v(126[12] 292[6])
    defparam i36303_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut_adj_1170 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n35375), .O(n17010));   // verilog/coms.v(126[12] 292[6])
    defparam i2_3_lut_4_lut_adj_1170.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_3_lut_adj_1171 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[1] ), .I3(GND_net), .O(n81));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_adj_1171.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1172 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state_31__N_2725 [3]), .I3(\FRAME_MATCHER.state[1] ), 
            .O(n34683));   // verilog/coms.v(126[12] 292[6])
    defparam i2_3_lut_4_lut_adj_1172.LUT_INIT = 16'h1000;
    SB_LUT4 i13150_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n17879));
    defparam i13150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n35016), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[8] [0]), .I3(n34984), .O(n15_adj_4389));
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i13151_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n17880));
    defparam i13151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1174 (.I0(n15_adj_4389), .I1(n4_adj_4390), .I2(n14_adj_4391), 
            .I3(n30543), .O(n36905));
    defparam i8_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(n36905), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n34871));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h9999;
    SB_LUT4 i13152_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n17881));
    defparam i13152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13153_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n17882));
    defparam i13153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1176 (.I0(n35179), .I1(n34906), .I2(n31283), 
            .I3(n35245), .O(n10_adj_4392));
    defparam i4_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1177 (.I0(n35022), .I1(n10_adj_4392), .I2(n16252), 
            .I3(GND_net), .O(n15435));
    defparam i5_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1178 (.I0(n16064), .I1(n35060), .I2(\data_in_frame[5] [3]), 
            .I3(GND_net), .O(n31283));
    defparam i2_3_lut_adj_1178.LUT_INIT = 16'h9696;
    SB_LUT4 n43178_bdd_4_lut (.I0(n43178), .I1(n38241), .I2(n38240), .I3(byte_transmit_counter[2]), 
            .O(n43181));
    defparam n43178_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13154_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n17883));
    defparam i13154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13155_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n17884));
    defparam i13155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13021_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n17750));
    defparam i13021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1179 (.I0(\data_in_frame[13] [6]), .I1(n34974), 
            .I2(\data_in_frame[14] [0]), .I3(n31283), .O(n12_adj_4393));
    defparam i5_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_LUT4 i13156_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n17885));
    defparam i13156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1180 (.I0(n15970), .I1(n12_adj_4393), .I2(n35173), 
            .I3(\data_in_frame[13] [7]), .O(n30999));
    defparam i6_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i13019_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n17748));
    defparam i13019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13157_3_lut_4_lut (.I0(n8_adj_4283), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n17886));
    defparam i13157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15957));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_15__7__I_0_3514_2_lut (.I0(\data_in_frame[15] [7]), 
            .I1(\data_in_frame[15] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_760));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_15__7__I_0_3514_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1182 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35185));
    defparam i1_2_lut_adj_1182.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1183 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [2]), 
            .I2(n35022), .I3(n16892), .O(n16_adj_4394));
    defparam i6_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i13020_3_lut_4_lut (.I0(n10_adj_4377), .I1(n34697), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n17749));
    defparam i13020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1184 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n35185), .I3(n30481), .O(n17_adj_4395));
    defparam i7_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1185 (.I0(n17_adj_4395), .I1(n30426), .I2(n16_adj_4394), 
            .I3(Kp_23__N_1276), .O(n36240));
    defparam i9_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_in_frame[19] [5]), .I1(n30999), .I2(n34871), 
            .I3(n31310), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1186 (.I0(Kp_23__N_760), .I1(\data_in_frame[16] [7]), 
            .I2(n15957), .I3(n31320), .O(n46));
    defparam i18_4_lut_adj_1186.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1187 (.I0(n31273), .I1(n36240), .I2(\data_in_frame[14] [1]), 
            .I3(n30525), .O(n47));
    defparam i19_4_lut_adj_1187.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_1188 (.I0(n35182), .I1(n35029), .I2(n35048), 
            .I3(\data_in_frame[19] [0]), .O(n45_adj_4396));
    defparam i17_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1189 (.I0(n35069), .I1(n35038), .I2(n35248), 
            .I3(\data_in_frame[20] [0]), .O(n44_adj_4397));
    defparam i16_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1190 (.I0(\data_in_frame[20] [6]), .I1(n34897), 
            .I2(\data_in_frame[21] [3]), .I3(Kp_23__N_1535), .O(n43_adj_4398));
    defparam i15_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n45_adj_4396), .I1(n47), .I2(n46), .I3(n48), 
            .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n15435), .I1(\data_in_frame[18] [6]), .I2(\data_in_frame[14] [7]), 
            .I3(n36773), .O(n49_adj_4399));
    defparam i21_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4399), .I1(n54), .I2(n43_adj_4398), 
            .I3(n44_adj_4397), .O(n35196));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1191 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[20] [2]), 
            .I2(\data_in_frame[20] [3]), .I3(GND_net), .O(n35269));
    defparam i2_3_lut_adj_1191.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15950));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1193 (.I0(n35137), .I1(n35209), .I2(n35108), 
            .I3(GND_net), .O(n30974));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_1193.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(n16716), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34796));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(n16706), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35209));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1196 (.I0(\data_in_frame[7] [3]), .I1(n35260), 
            .I2(n35221), .I3(n34987), .O(n36645));
    defparam i3_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1197 (.I0(n35160), .I1(n16716), .I2(\data_in_frame[7] [0]), 
            .I3(n16666), .O(n14_adj_4400));
    defparam i6_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1198 (.I0(\data_in_frame[9] [2]), .I1(n14_adj_4400), 
            .I2(n10_adj_4303), .I3(\data_in_frame[7] [1]), .O(n31368));
    defparam i7_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35115));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(\data_in_frame[9] [3]), .I1(n35221), 
            .I2(n15_adj_4401), .I3(n16716), .O(n10_adj_4402));
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n34675), 
            .I2(n10337), .I3(n3894), .O(n34));   // verilog/coms.v(126[12] 292[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 select_371_Select_2_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), 
            .I1(n34675), .I2(n3894), .I3(\FRAME_MATCHER.state_31__N_2661[2] ), 
            .O(n7));   // verilog/coms.v(126[12] 292[6])
    defparam select_371_Select_2_i7_3_lut_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(\FRAME_MATCHER.state[1] ), .I1(n34675), 
            .I2(n3894), .I3(GND_net), .O(n34681));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'h0808;
    SB_LUT4 i6_4_lut_adj_1202 (.I0(n35209), .I1(\data_in_frame[6] [7]), 
            .I2(n34796), .I3(n16641), .O(n14_adj_4404));   // verilog/coms.v(69[16:62])
    defparam i6_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1203 (.I0(\data_in_frame[9] [1]), .I1(n14_adj_4404), 
            .I2(n10_adj_4405), .I3(\data_in_frame[6] [0]), .O(n31094));   // verilog/coms.v(69[16:62])
    defparam i7_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(n31368), .I1(n36645), .I2(GND_net), 
            .I3(GND_net), .O(n15970));
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(n31094), .I1(n34974), .I2(GND_net), 
            .I3(GND_net), .O(n31030));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35108));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35173));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1208 (.I0(\FRAME_MATCHER.state [0]), .I1(n63_adj_4296), 
            .I2(n63_adj_4292), .I3(n63_adj_4285), .O(\FRAME_MATCHER.state_31__N_2661[0] ));
    defparam i3_4_lut_adj_1208.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35170));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\data_in_frame[9] [5]), .I1(n35781), 
            .I2(GND_net), .I3(GND_net), .O(n35060));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1211 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [6]), 
            .I2(n16430), .I3(GND_net), .O(n35105));   // verilog/coms.v(69[16:62])
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1212 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n35266));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1213 (.I0(\data_in_frame[3] [3]), .I1(n35212), 
            .I2(n35122), .I3(\data_in_frame[1] [2]), .O(n16252));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1214 (.I0(\data_in_frame[5] [5]), .I1(n31329), 
            .I2(\data_in_frame[5] [0]), .I3(\data_in_frame[5] [3]), .O(n28_adj_4406));
    defparam i12_4_lut_adj_1214.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4407));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31408_4_lut (.I0(n19_adj_4407), .I1(\data_out_frame[22] [7]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38238));
    defparam i31408_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33809_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n40641));   // verilog/coms.v(104[34:55])
    defparam i33809_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4408));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31409_3_lut (.I0(n43253), .I1(n38238), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38239));
    defparam i31409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31359_4_lut (.I0(n5_adj_4408), .I1(n40641), .I2(n40044), 
            .I3(\byte_transmit_counter[0] ), .O(n38189));
    defparam i31359_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31361_4_lut (.I0(n38189), .I1(n38239), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38191));
    defparam i31361_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10_4_lut_adj_1215 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(n35082), .I3(\data_in_frame[4] [0]), .O(n26_adj_4409));
    defparam i10_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4410));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33804_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40636));   // verilog/coms.v(104[34:55])
    defparam i33804_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4411));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31405_4_lut (.I0(n19_adj_4410), .I1(\data_out_frame[22] [6]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38235));
    defparam i31405_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11_4_lut_adj_1216 (.I0(n35781), .I1(n34987), .I2(n35105), 
            .I3(n34864), .O(n27_adj_4412));
    defparam i11_4_lut_adj_1216.LUT_INIT = 16'h9669;
    SB_LUT4 i31406_3_lut (.I0(n43247), .I1(n38235), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38236));
    defparam i31406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31389_4_lut (.I0(n5_adj_4411), .I1(n40636), .I2(n40044), 
            .I3(\byte_transmit_counter[0] ), .O(n38219));
    defparam i31389_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i9_4_lut_adj_1217 (.I0(n35212), .I1(\data_in_frame[5] [6]), 
            .I2(n16716), .I3(n14136), .O(n25_adj_4413));
    defparam i9_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1218 (.I0(n25_adj_4413), .I1(n27_adj_4412), .I2(n26_adj_4409), 
            .I3(n28_adj_4406), .O(n36911));
    defparam i15_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i31391_4_lut (.I0(n38219), .I1(n38236), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38221));
    defparam i31391_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i20_4_lut_adj_1219 (.I0(n34877), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[8] [7]), .O(n48_adj_4414));
    defparam i20_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i31390_3_lut (.I0(n43265), .I1(n43259), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38220));
    defparam i31390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1220 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[7] [2]), 
            .I2(n36911), .I3(n35266), .O(n46_adj_4415));
    defparam i18_4_lut_adj_1220.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1221 (.I0(n35173), .I1(n35108), .I2(n35167), 
            .I3(n35045), .O(n47_adj_4416));
    defparam i19_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4417));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40627));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4418));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31402_4_lut (.I0(n19_adj_4417), .I1(\data_out_frame[22] [5]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38232));
    defparam i31402_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31403_3_lut (.I0(n43241), .I1(n38232), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38233));
    defparam i31403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31386_4_lut (.I0(n5_adj_4418), .I1(\byte_transmit_counter[0] ), 
            .I2(n40044), .I3(n40627), .O(n38216));
    defparam i31386_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i17_4_lut_adj_1222 (.I0(\data_in_frame[11] [0]), .I1(n35060), 
            .I2(n35170), .I3(n34867), .O(n45_adj_4419));
    defparam i17_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1223 (.I0(\data_in_frame[6] [3]), .I1(n34906), 
            .I2(n35242), .I3(n15950), .O(n44_adj_4420));
    defparam i16_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1224 (.I0(n35115), .I1(n16178), .I2(\data_in_frame[12] [3]), 
            .I3(n30974), .O(n43_adj_4421));
    defparam i15_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i31388_4_lut (.I0(n38216), .I1(n38233), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38218));
    defparam i31388_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i26_4_lut_adj_1225 (.I0(n45_adj_4419), .I1(n47_adj_4416), .I2(n46_adj_4415), 
            .I3(n48_adj_4414), .O(n54_adj_4422));
    defparam i26_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i31387_3_lut (.I0(n43277), .I1(n43271), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38217));
    defparam i31387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_4_lut_adj_1226 (.I0(n16641), .I1(\data_in_frame[10] [1]), 
            .I2(n15426), .I3(\data_in_frame[10] [3]), .O(n49_adj_4423));
    defparam i21_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_1227 (.I0(n49_adj_4423), .I1(n54_adj_4422), .I2(n43_adj_4421), 
            .I3(n44_adj_4420), .O(n35245));
    defparam i27_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4424));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4425));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4426));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31399_4_lut (.I0(n19_adj_4424), .I1(\data_out_frame[22] [4]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38229));
    defparam i31399_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(n36645), .I1(n34974), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n30426));
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h6969;
    SB_LUT4 i31400_3_lut (.I0(n43235), .I1(n38229), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38230));
    defparam i31400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31383_3_lut (.I0(n5_adj_4426), .I1(n6_adj_4425), .I2(n40044), 
            .I3(GND_net), .O(n38213));
    defparam i31383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31385_4_lut (.I0(n38213), .I1(n38230), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38215));
    defparam i31385_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31384_3_lut (.I0(n43289), .I1(n43283), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38214));
    defparam i31384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4427));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4428));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4429));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31396_4_lut (.I0(n19_adj_4427), .I1(\data_out_frame[22] [3]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38226));
    defparam i31396_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31397_3_lut (.I0(n43229), .I1(n38226), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38227));
    defparam i31397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31380_3_lut (.I0(n5_adj_4429), .I1(n6_adj_4428), .I2(n40044), 
            .I3(GND_net), .O(n38210));
    defparam i31380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31382_4_lut (.I0(n38210), .I1(n38227), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38212));
    defparam i31382_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_3_lut_adj_1229 (.I0(n30426), .I1(n35245), .I2(\data_in_frame[12] [0]), 
            .I3(GND_net), .O(n35006));
    defparam i2_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i31381_3_lut (.I0(n43301), .I1(n43295), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38211));
    defparam i31381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4430));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31393_4_lut (.I0(n19_adj_4430), .I1(\data_out_frame[22] [2]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38223));
    defparam i31393_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4431));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha003;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4432));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31394_3_lut (.I0(n43223), .I1(n38223), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38224));
    defparam i31394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'heeee;
    SB_LUT4 i31377_3_lut (.I0(n5_adj_4432), .I1(n6_adj_4431), .I2(n40044), 
            .I3(GND_net), .O(n38207));
    defparam i31377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1231 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [0]), .O(n14_adj_4433));   // verilog/coms.v(126[12] 292[6])
    defparam i6_4_lut_adj_1231.LUT_INIT = 16'hfffe;
    SB_LUT4 i31379_4_lut (.I0(n38207), .I1(n38224), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38209));
    defparam i31379_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16892));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i33782_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40613));   // verilog/coms.v(104[34:55])
    defparam i33782_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4434));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\data_in_frame[10] [6]), .I1(Kp_23__N_1183), 
            .I2(GND_net), .I3(GND_net), .O(n34867));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 i31374_4_lut (.I0(n5_adj_4434), .I1(n40613), .I2(n40044), 
            .I3(\byte_transmit_counter[0] ), .O(n38204));
    defparam i31374_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31376_4_lut (.I0(n38204), .I1(n43187), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38206));
    defparam i31376_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36348 (.I0(\byte_transmit_counter[1] ), 
            .I1(n38249), .I2(n38250), .I3(byte_transmit_counter[2]), .O(n43172));
    defparam byte_transmit_counter_1__bdd_4_lut_36348.LUT_INIT = 16'he4aa;
    SB_LUT4 n43172_bdd_4_lut (.I0(n43172), .I1(n38247), .I2(n38246), .I3(byte_transmit_counter[2]), 
            .O(n43175));
    defparam n43172_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1234 (.I0(Kp_23__N_1276), .I1(\data_in_frame[8] [5]), 
            .I2(n35134), .I3(n6_adj_4435), .O(n34969));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4436));
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1236 (.I0(\FRAME_MATCHER.state_31__N_2725 [3]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n24684), .I3(\FRAME_MATCHER.state [2]), .O(n37203));
    defparam i3_4_lut_adj_1236.LUT_INIT = 16'h0040;
    SB_LUT4 i2_4_lut_adj_1237 (.I0(\FRAME_MATCHER.state [0]), .I1(n29), 
            .I2(n24684), .I3(\FRAME_MATCHER.state [2]), .O(n35855));
    defparam i2_4_lut_adj_1237.LUT_INIT = 16'hc800;
    SB_LUT4 i36290_4_lut (.I0(n35855), .I1(n37203), .I2(n24676), .I3(n6_adj_4436), 
            .O(n36824));
    defparam i36290_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i4_4_lut_adj_1238 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [1]), .I3(n34969), .O(n10_adj_4437));
    defparam i4_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1239 (.I0(n16354), .I1(\data_in_frame[6] [2]), 
            .I2(n16663), .I3(\data_in_frame[6] [3]), .O(Kp_23__N_1183));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1240 (.I0(Kp_23__N_1189), .I1(n35266), .I2(Kp_23__N_1186), 
            .I3(GND_net), .O(n34955));
    defparam i2_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1241 (.I0(\data_in_frame[10] [5]), .I1(Kp_23__N_1183), 
            .I2(\data_in_frame[8] [4]), .I3(n16096), .O(n16382));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1242 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4438));
    defparam i2_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1243 (.I0(\data_in_frame[13] [1]), .I1(n14_adj_4360), 
            .I2(n10_adj_4438), .I3(n34969), .O(n31386));
    defparam i7_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[17] [3]), .I1(n30625), 
            .I2(GND_net), .I3(GND_net), .O(n35051));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[14] [7]), .I1(n34981), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4439));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1246 (.I0(n30481), .I1(n31439), .I2(\data_in_frame[12] [7]), 
            .I3(n6_adj_4439), .O(n15414));
    defparam i4_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1055_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4348), .I3(GND_net), .O(n4349));
    defparam mux_1055_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1247 (.I0(n9), .I1(n14_adj_4433), .I2(\data_in_frame[0] [6]), 
            .I3(\data_in_frame[0] [7]), .O(n13355));   // verilog/coms.v(126[12] 292[6])
    defparam i7_4_lut_adj_1247.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1248 (.I0(\data_in_frame[22] [7]), .I1(\data_in_frame[22] [1]), 
            .I2(\data_in_frame[22] [2]), .I3(\data_in_frame[22] [3]), .O(n8_adj_4440));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1249 (.I0(\data_in_frame[22] [4]), .I1(n8_adj_4440), 
            .I2(\data_in_frame[22] [5]), .I3(\data_in_frame[22] [6]), .O(Kp_23__N_731));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1250 (.I0(n15414), .I1(n35051), .I2(\data_in_frame[15] [0]), 
            .I3(n31386), .O(n35248));
    defparam i1_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[22] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16869));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[10] [2]), .I1(n6_adj_4441), 
            .I2(GND_net), .I3(GND_net), .O(n34952));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1253 (.I0(n16273), .I1(n16503), .I2(\data_in_frame[10] [3]), 
            .I3(GND_net), .O(n30481));
    defparam i2_3_lut_adj_1253.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(n31394), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4442));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_in_frame[12] [4]), .I1(n30481), 
            .I2(GND_net), .I3(GND_net), .O(n31275));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[21] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16188));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1257 (.I0(\data_in_frame[14] [5]), .I1(n34845), 
            .I2(\data_in_frame[12] [3]), .I3(n31275), .O(n30843));
    defparam i3_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1258 (.I0(\data_in_frame[6] [1]), .I1(n16448), 
            .I2(n16033), .I3(GND_net), .O(n34877));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1258.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\FRAME_MATCHER.state [31]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4357));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1260 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[5] [6]), 
            .I2(n34806), .I3(n6_adj_4359), .O(n16503));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1261 (.I0(\data_in_frame[6] [2]), .I1(n34877), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n16096));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 i18880_2_lut (.I0(\FRAME_MATCHER.state [30]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23594));
    defparam i18880_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1262 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[6] [0]), 
            .I2(n16448), .I3(GND_net), .O(n34984));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\FRAME_MATCHER.state [29]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4355));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1264 (.I0(\data_in_frame[7] [7]), .I1(n34984), 
            .I2(n16053), .I3(GND_net), .O(n16273));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1264.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(\FRAME_MATCHER.state [28]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34219));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\FRAME_MATCHER.state [27]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4353));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\FRAME_MATCHER.state [26]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34217));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h8888;
    SB_LUT4 i18879_2_lut (.I0(\FRAME_MATCHER.state [25]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23592));
    defparam i18879_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\FRAME_MATCHER.state [24]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34221));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(n16096), .I1(n16503), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1276));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\FRAME_MATCHER.state [23]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4351));
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1271 (.I0(Kp_23__N_1276), .I1(n35167), .I2(n16273), 
            .I3(\data_in_frame[12] [5]), .O(n12_adj_4444));   // verilog/coms.v(73[16:43])
    defparam i5_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(\FRAME_MATCHER.state [22]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34187));
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1273 (.I0(n16252), .I1(n12_adj_4444), .I2(\data_in_frame[14] [6]), 
            .I3(n34952), .O(n34981));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\FRAME_MATCHER.state [21]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4349));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\FRAME_MATCHER.state [20]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34215));
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1276 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[20] [7]), 
            .I2(n34981), .I3(\data_in_frame[12] [4]), .O(n6_adj_4445));
    defparam i1_4_lut_adj_1276.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1277 (.I0(\FRAME_MATCHER.state [0]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n34603), .I3(n27212), .O(n19504));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1277.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\FRAME_MATCHER.state [19]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34213));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h8888;
    SB_LUT4 i18878_2_lut (.I0(\FRAME_MATCHER.state [18]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23590));
    defparam i18878_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\FRAME_MATCHER.state [17]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23588));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[10] [6]), .I1(Kp_23__N_1183), 
            .I2(\data_in_frame[8] [4]), .I3(\data_in_frame[11] [0]), .O(n10_adj_4388));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1280 (.I0(n1), .I1(n16053), .I2(n15_adj_4401), 
            .I3(n31392), .O(n28_adj_4446));   // verilog/coms.v(228[9:81])
    defparam i12_4_lut_adj_1280.LUT_INIT = 16'hfffb;
    SB_LUT4 i10_4_lut_adj_1281 (.I0(n16663), .I1(n16666), .I2(n16706), 
            .I3(n16716), .O(n26_adj_4447));   // verilog/coms.v(228[9:81])
    defparam i10_4_lut_adj_1281.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\FRAME_MATCHER.state [16]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34211));
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h8888;
    SB_LUT4 i28611_2_lut_3_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n34603), 
            .I2(n27212), .I3(GND_net), .O(n35375));
    defparam i28611_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(\data_in_frame[18] [5]), .I1(n30843), 
            .I2(n16188), .I3(n6_adj_4445), .O(n34997));
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\FRAME_MATCHER.state [15]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4347));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1285 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(n34793), .I3(\data_out_frame[11] [6]), .O(n35164));
    defparam i1_2_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\FRAME_MATCHER.state [14]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34209));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n34934));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\FRAME_MATCHER.state [13]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34207));
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16889));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n16482));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i18876_2_lut (.I0(\FRAME_MATCHER.state [12]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23586));
    defparam i18876_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[7] [4]), .I1(n34987), 
            .I2(GND_net), .I3(GND_net), .O(n30543));
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1292 (.I0(n16292), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[5] [3]), .O(n4_adj_4390));
    defparam i1_2_lut_3_lut_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[9] [4]), .I1(n35160), 
            .I2(GND_net), .I3(GND_net), .O(n35260));
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\FRAME_MATCHER.state [11]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34205));
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1295 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[7] [6]), .O(n6_adj_4448));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n16312));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i18875_2_lut (.I0(\FRAME_MATCHER.state [10]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23584));
    defparam i18875_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16064));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1298 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[7] [4]), .O(n34930));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\FRAME_MATCHER.state [9]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34203));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34834));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1301 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n34911));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1301.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\FRAME_MATCHER.state [8]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34201));
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n6_adj_4449));
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16178));
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1305 (.I0(\FRAME_MATCHER.state [7]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34199));
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1306 (.I0(\data_out_frame[7] [3]), .I1(n16072), 
            .I2(\data_out_frame[11] [5]), .I3(\data_out_frame[9] [4]), .O(n35203));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\FRAME_MATCHER.state [6]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34197));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1308 (.I0(\data_in_frame[9] [7]), .I1(n6_adj_4441), 
            .I2(n16053), .I3(\data_in_frame[7] [5]), .O(n12_adj_4450));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\FRAME_MATCHER.state [5]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n34195));
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1310 (.I0(n1211), .I1(n34), .I2(n15876), .I3(n10337), 
            .O(n4_adj_4443));
    defparam i2_4_lut_adj_1310.LUT_INIT = 16'hcecc;
    SB_LUT4 i6_4_lut_adj_1311 (.I0(n16229), .I1(n12_adj_4450), .I2(\data_in_frame[10] [1]), 
            .I3(n34834), .O(n34845));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1312 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n16499));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n6_adj_4451));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i18874_2_lut (.I0(\FRAME_MATCHER.state [4]), .I1(n4_adj_4443), 
            .I2(GND_net), .I3(GND_net), .O(n23582));
    defparam i18874_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(n16252), .I1(n4_adj_4390), .I2(GND_net), 
            .I3(GND_net), .O(n16229));
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1315 (.I0(n2957), .I1(\FRAME_MATCHER.i_31__N_2625 ), 
            .I2(n10337), .I3(GND_net), .O(n37));
    defparam i1_3_lut_adj_1315.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_3_lut_adj_1316 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n16124));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1317 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(n16020), .O(n35236));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(n10337), .I1(n2774), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4305));   // verilog/coms.v(154[6] 156[9])
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(n49), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n27214));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_in_frame[9] [5]), .I1(n31392), 
            .I2(GND_net), .I3(GND_net), .O(n35239));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n19503), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n34683), .I3(n27214), .O(n34193));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'hdc50;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[11] [2]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n16376));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n16404));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35242));
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1325 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(n10_adj_4452), .I3(\data_out_frame[13] [1]), .O(n34937));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(\data_out_frame[6] [6]), .I1(n35151), 
            .I2(\data_out_frame[8] [5]), .I3(n1336), .O(n34940));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 select_371_Select_1_i5_4_lut (.I0(n63_adj_4285), .I1(\FRAME_MATCHER.i_31__N_2625 ), 
            .I2(n2957), .I3(n92[1]), .O(n5_adj_4453));
    defparam select_371_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 i5_3_lut_4_lut_adj_1327 (.I0(n31273), .I1(n34775), .I2(n30861), 
            .I3(\data_in_frame[24] [1]), .O(n14_adj_4454));
    defparam i5_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1328 (.I0(n63), .I1(n29937), .I2(n5_adj_4453), 
            .I3(n1_adj_4455), .O(n43574));
    defparam i3_4_lut_adj_1328.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_4_lut_adj_1329 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[8] [7]), .O(n6_adj_4456));
    defparam i1_2_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1330 (.I0(\data_out_frame[6] [6]), .I1(n34934), 
            .I2(n16482), .I3(n35078), .O(n34809));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1331 (.I0(\data_out_frame[20] [5]), .I1(n35097), 
            .I2(n31342), .I3(GND_net), .O(n37115));
    defparam i2_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(n35035), .I1(n35193), .I2(GND_net), 
            .I3(GND_net), .O(n35194));
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(\data_in_frame[9] [6]), .I1(n30543), 
            .I2(\data_in_frame[7] [5]), .I3(\data_in_frame[11] [7]), .O(n34906));
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1334 (.I0(\data_out_frame[19] [1]), .I1(n31340), 
            .I2(n35224), .I3(n34966), .O(n36454));
    defparam i2_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1335 (.I0(\data_out_frame[14] [5]), .I1(n16060), 
            .I2(n34824), .I3(\data_out_frame[15] [0]), .O(n6_adj_4457));
    defparam i1_2_lut_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1336 (.I0(\data_out_frame[17] [2]), .I1(n36635), 
            .I2(n34966), .I3(\data_out_frame[19] [3]), .O(n36358));
    defparam i2_3_lut_4_lut_adj_1336.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(\data_out_frame[20] [4]), .I1(n16815), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4458));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1338 (.I0(n34755), .I1(\data_out_frame[16] [2]), 
            .I2(n35142), .I3(n6_adj_4458), .O(n35193));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n35072));
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1340 (.I0(n34886), .I1(n35142), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4459));
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1341 (.I0(\data_out_frame[16] [3]), .I1(n31306), 
            .I2(n35075), .I3(n6_adj_4459), .O(n31342));
    defparam i4_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1342 (.I0(n31281), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n35176));
    defparam i2_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1343 (.I0(n34991), .I1(n35176), .I2(n30432), 
            .I3(GND_net), .O(n31390));
    defparam i2_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1344 (.I0(n35239), .I1(n16229), .I2(n34845), 
            .I3(n16178), .O(n14_adj_4460));
    defparam i6_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1345 (.I0(\data_out_frame[20] [7]), .I1(n35035), 
            .I2(n35057), .I3(GND_net), .O(n7_adj_4461));
    defparam i2_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1346 (.I0(\data_out_frame[20] [2]), .I1(n37156), 
            .I2(\data_out_frame[18][1] ), .I3(n30432), .O(n35057));
    defparam i1_3_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n35075));
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1348 (.I0(n16593), .I1(n31281), .I2(\data_out_frame[16] [0]), 
            .I3(n6_adj_4302), .O(n37156));
    defparam i4_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1349 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_4460), 
            .I2(n10_adj_4304), .I3(n16064), .O(n34848));
    defparam i7_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1350 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[12] [0]), 
            .I2(n35016), .I3(\data_in_frame[14] [2]), .O(n18_adj_4462));
    defparam i7_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[18][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4463));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(n34755), .I1(n35075), .I2(n37156), 
            .I3(n6_adj_4463), .O(n35035));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1353 (.I0(\data_in_frame[3] [0]), .I1(n35122), 
            .I2(n34978), .I3(n6_adj_4363), .O(n31394));   // verilog/coms.v(68[16:69])
    defparam i2_3_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1354 (.I0(n16252), .I1(n4_adj_4390), .I2(n16_adj_4442), 
            .I3(n34987), .O(n27_adj_4464));   // verilog/coms.v(228[9:81])
    defparam i11_4_lut_adj_1354.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1355 (.I0(n16354), .I1(n6_adj_4441), .I2(n16033), 
            .I3(n16448), .O(n25_adj_4465));   // verilog/coms.v(228[9:81])
    defparam i9_4_lut_adj_1355.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1356 (.I0(n25_adj_4465), .I1(n27_adj_4464), .I2(n26_adj_4447), 
            .I3(n28_adj_4446), .O(n31_adj_4260));   // verilog/coms.v(228[9:81])
    defparam i15_4_lut_adj_1356.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[11] [6]), .I1(n16252), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4466));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1357 (.I0(n31_adj_4260), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n13355), .I3(GND_net), .O(n4348));
    defparam i2_3_lut_adj_1357.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(n35035), .I1(n35057), .I2(GND_net), 
            .I3(GND_net), .O(n34964));
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[10] [0]), .I3(GND_net), .O(n35016));
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1360 (.I0(\data_in_frame[3] [0]), .I1(n35122), 
            .I2(\data_in_frame[0] [4]), .I3(n34883), .O(n34900));   // verilog/coms.v(68[16:69])
    defparam i2_3_lut_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1361 (.I0(\data_out_frame[18] [5]), .I1(n34782), 
            .I2(n1765), .I3(n31306), .O(n35097));
    defparam i3_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1362 (.I0(n31342), .I1(n35193), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n34829));
    defparam i2_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1363 (.I0(\data_out_frame[20] [1]), .I1(n34829), 
            .I2(n35097), .I3(GND_net), .O(n8_adj_4467));
    defparam i3_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i13198_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n17927));
    defparam i13198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_4_lut_adj_1364 (.I0(n31390), .I1(n7_adj_4461), .I2(n36296), 
            .I3(n8_adj_4467), .O(n35055));
    defparam i2_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1365 (.I0(\data_in_frame[7] [2]), .I1(n18_adj_4462), 
            .I2(\data_in_frame[7] [6]), .I3(n35260), .O(n20_adj_4468));
    defparam i9_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1366 (.I0(n35239), .I1(n20_adj_4468), .I2(n16_adj_4466), 
            .I3(n16053), .O(n30525));
    defparam i10_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4469));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1368 (.I0(n35019), .I1(n16660), .I2(n35176), 
            .I3(n6_adj_4469), .O(n34994));
    defparam i4_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(n34994), .I1(n35055), .I2(GND_net), 
            .I3(GND_net), .O(n34972));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1370 (.I0(n30889), .I1(n35088), .I2(n34972), 
            .I3(n16130), .O(n37102));
    defparam i3_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1371 (.I0(n16404), .I1(n1336), .I2(n16753), .I3(n16857), 
            .O(n12_adj_4470));
    defparam i5_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1372 (.I0(n30525), .I1(n34848), .I2(\data_in_frame[16] [4]), 
            .I3(GND_net), .O(n30562));
    defparam i2_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1373 (.I0(\data_out_frame[17] [4]), .I1(n12_adj_4470), 
            .I2(n16736), .I3(\data_out_frame[13] [2]), .O(n35019));
    defparam i6_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1374 (.I0(\data_out_frame[19] [5]), .I1(n35019), 
            .I2(\data_out_frame[19] [4]), .I3(n31427), .O(n36919));
    defparam i3_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 select_371_Select_1_i1_3_lut_4_lut (.I0(n92[1]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n34675), .I3(n9001), .O(n1_adj_4455));
    defparam select_371_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'h2030;
    SB_LUT4 i3_4_lut_adj_1375 (.I0(n15974), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(\data_out_frame[15] [2]), 
            .O(n16857));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1376 (.I0(\data_in_frame[21] [4]), .I1(\data_in_frame[23] [7]), 
            .I2(\data_in_frame[17] [1]), .I3(\data_in_frame[21] [7]), .O(n28_adj_4471));
    defparam i12_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1377 (.I0(n34924), .I1(\data_out_frame[6] [3]), 
            .I2(n16857), .I3(n35148), .O(n10_adj_4472));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1378 (.I0(n16370), .I1(n10_adj_4472), .I2(n16401), 
            .I3(GND_net), .O(n30889));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1379 (.I0(\data_out_frame[17] [3]), .I1(n35257), 
            .I2(n35224), .I3(n30889), .O(n36643));
    defparam i3_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_out_frame[17] [2]), .I1(n36635), 
            .I2(GND_net), .I3(GND_net), .O(n31427));
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1381 (.I0(n31435), .I1(n16886), .I2(\data_out_frame[19] [2]), 
            .I3(GND_net), .O(n34966));
    defparam i2_3_lut_adj_1381.LUT_INIT = 16'h6969;
    SB_LUT4 i13205_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n17934));
    defparam i13205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13204_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n17933));
    defparam i13204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1382 (.I0(n34997), .I1(\data_in_frame[21] [6]), 
            .I2(n30562), .I3(\data_in_frame[19] [3]), .O(n26_adj_4473));
    defparam i10_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1383 (.I0(n16869), .I1(n35248), .I2(Kp_23__N_731), 
            .I3(\data_in_frame[20] [5]), .O(n27_adj_4474));
    defparam i11_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1384 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[14] [7]), .I3(n6_adj_4457), .O(n35224));
    defparam i4_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i13203_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n17932));
    defparam i13203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1385 (.I0(n16839), .I1(n16699), .I2(n16417), 
            .I3(\data_out_frame[14] [2]), .O(n34886));
    defparam i3_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(n16212), .I1(n34886), .I2(GND_net), 
            .I3(GND_net), .O(n1765));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1387 (.I0(n34921), .I1(n1765), .I2(\data_out_frame[19] [1]), 
            .I3(n35145), .O(n10_adj_4475));
    defparam i4_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1388 (.I0(\data_out_frame[18] [6]), .I1(n10_adj_4475), 
            .I2(n31340), .I3(GND_net), .O(n36072));
    defparam i5_3_lut_adj_1388.LUT_INIT = 16'h6969;
    SB_LUT4 i9_4_lut_adj_1389 (.I0(n35269), .I1(n35785), .I2(\data_in_frame[21] [0]), 
            .I3(n35196), .O(n25_adj_4476));
    defparam i9_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1390 (.I0(\data_out_frame[12] [5]), .I1(n15974), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4477));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1391 (.I0(n34746), .I1(n35072), .I2(n30562), 
            .I3(\data_in_frame[23] [4]), .O(n12_adj_4478));
    defparam i5_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1392 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(n31322), .I3(n6_adj_4477), .O(n16886));
    defparam i4_4_lut_adj_1392.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(n16299), .I1(n34903), .I2(GND_net), 
            .I3(GND_net), .O(n30491));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1394 (.I0(n34746), .I1(n30625), .I2(n16610), 
            .I3(n35069), .O(n10_adj_4479));
    defparam i4_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\data_out_frame[12] [4]), .I1(n30994), 
            .I2(GND_net), .I3(GND_net), .O(n31322));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h6666;
    SB_LUT4 i13202_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n17931));
    defparam i13202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1396 (.I0(n15422), .I1(n31322), .I2(n35233), 
            .I3(n34812), .O(n16_adj_4480));
    defparam i6_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1397 (.I0(\data_out_frame[12] [6]), .I1(n35188), 
            .I2(n35254), .I3(n16401), .O(n17_adj_4481));
    defparam i7_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i13201_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n17930));
    defparam i13201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1398 (.I0(n17_adj_4481), .I1(n30491), .I2(n16_adj_4480), 
            .I3(n15489), .O(n36635));
    defparam i9_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1399 (.I0(\data_in_frame[22] [3]), .I1(n30859), 
            .I2(Kp_23__N_1783), .I3(GND_net), .O(n8_adj_4482));
    defparam i3_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(\data_out_frame[12] [5]), .I1(n15489), 
            .I2(GND_net), .I3(GND_net), .O(n35148));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1401 (.I0(n16742), .I1(n16791), .I2(n34934), 
            .I3(n34759), .O(n35025));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1402 (.I0(n35148), .I1(n34762), .I2(\data_out_frame[13] [1]), 
            .I3(n35157), .O(n10_adj_4483));
    defparam i4_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1403 (.I0(n35078), .I1(n35025), .I2(n10_adj_4483), 
            .I3(\data_out_frame[13] [0]), .O(n35188));
    defparam i1_4_lut_adj_1403.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1404 (.I0(n16060), .I1(n34824), .I2(\data_out_frame[15] [0]), 
            .I3(GND_net), .O(n35118));
    defparam i2_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i13200_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n17929));
    defparam i13200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut_adj_1405 (.I0(\data_in_frame[21] [4]), .I1(n10_adj_4479), 
            .I2(\data_in_frame[23] [5]), .I3(GND_net), .O(n36985));
    defparam i5_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1406 (.I0(n30424), .I1(\data_out_frame[13] [5]), 
            .I2(n34790), .I3(n1713), .O(n35157));   // verilog/coms.v(83[17:63])
    defparam i3_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1407 (.I0(n35251), .I1(n30549), .I2(Kp_23__N_731), 
            .I3(GND_net), .O(n11));
    defparam i3_3_lut_adj_1407.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1408 (.I0(\data_out_frame[15] [1]), .I1(n34937), 
            .I2(n35157), .I3(n34940), .O(n35233));   // verilog/coms.v(83[17:63])
    defparam i3_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16791));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1410 (.I0(\data_out_frame[8] [6]), .I1(n1558), 
            .I2(n16875), .I3(n6_adj_4456), .O(n34903));
    defparam i4_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35145));
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1412 (.I0(\FRAME_MATCHER.state [3]), .I1(n10337), 
            .I2(n2774), .I3(n34), .O(n34053));
    defparam i1_3_lut_4_lut_adj_1412.LUT_INIT = 16'haa80;
    SB_LUT4 i5_4_lut_adj_1413 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[23] [2]), 
            .I2(\data_in_frame[18] [4]), .I3(n36905), .O(n14_adj_4484));
    defparam i5_4_lut_adj_1413.LUT_INIT = 16'h9669;
    SB_LUT4 i13199_3_lut_4_lut (.I0(n24351), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n17928));
    defparam i13199_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1414 (.I0(n36954), .I1(n34809), .I2(n35118), 
            .I3(n35188), .O(n18_adj_4485));
    defparam i7_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1415 (.I0(n35072), .I1(\data_in_frame[21] [1]), 
            .I2(n30843), .I3(n35032), .O(n15_adj_4486));
    defparam i6_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1416 (.I0(n35145), .I1(n34903), .I2(n35042), 
            .I3(n16324), .O(n19_adj_4487));
    defparam i8_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1417 (.I0(n19_adj_4487), .I1(n36635), .I2(n18_adj_4485), 
            .I3(n12), .O(n31340));
    defparam i10_4_lut_adj_1417.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1418 (.I0(\data_in_frame[22] [7]), .I1(\data_in_frame[22] [6]), 
            .I2(\data_in_frame[20] [4]), .I3(\data_in_frame[18] [3]), .O(n16_adj_4488));
    defparam i6_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35257));
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_out_frame[19] [1]), .I1(n31340), 
            .I2(GND_net), .I3(GND_net), .O(n35206));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1421 (.I0(\data_out_frame[19] [6]), .I1(n34771), 
            .I2(\data_out_frame[19] [5]), .I3(n16029), .O(n35088));
    defparam i3_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1422 (.I0(\data_in_frame[18] [2]), .I1(n30562), 
            .I2(n35032), .I3(n16160), .O(n17_adj_4489));
    defparam i7_4_lut_adj_1422.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1423 (.I0(\data_out_frame[19] [0]), .I1(n31381), 
            .I2(GND_net), .I3(GND_net), .O(n34921));
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1424 (.I0(n34793), .I1(n35154), .I2(\data_out_frame[11] [5]), 
            .I3(\data_out_frame[7] [5]), .O(n12_adj_4490));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1425 (.I0(\data_out_frame[12] [0]), .I1(n12_adj_4490), 
            .I2(n35236), .I3(n16742), .O(n16815));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1426 (.I0(n16889), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[23] [3]), .I3(n34997), .O(n10_adj_4491));
    defparam i4_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i35570_2_lut (.I0(n19260), .I1(\data_out_frame[18] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n42402));   // verilog/coms.v(95[12:26])
    defparam i35570_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1427 (.I0(n16815), .I1(n31421), .I2(\data_out_frame[18] [5]), 
            .I3(n42402), .O(n12_adj_4492));
    defparam i5_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1428 (.I0(n16324), .I1(n12_adj_4492), .I2(n34921), 
            .I3(\data_out_frame[16] [7]), .O(n36296));
    defparam i6_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1429 (.I0(n788), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n34675), .I3(n10337), .O(n49));
    defparam i1_3_lut_4_lut_adj_1429.LUT_INIT = 16'h1000;
    SB_LUT4 i9_4_lut_adj_1430 (.I0(n17_adj_4489), .I1(\data_in_frame[18] [4]), 
            .I2(n16_adj_4488), .I3(\data_in_frame[23] [0]), .O(n36936));
    defparam i9_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1431 (.I0(n35206), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[17] [5]), .I3(n35257), .O(n10_adj_4493));
    defparam i4_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1432 (.I0(n35088), .I1(n10_adj_4493), .I2(\data_out_frame[19] [2]), 
            .I3(GND_net), .O(n31421));
    defparam i5_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut (.I0(n15_adj_4401), .I1(n34900), .I2(n34978), 
            .I3(\data_in_frame[5] [0]), .O(n35160));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1433 (.I0(n16499), .I1(n34821), .I2(\data_out_frame[11] [1]), 
            .I3(n16376), .O(n1558));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1434 (.I0(n1558), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[13] [3]), .I3(GND_net), .O(n34771));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_1434.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[10] [4]), .I3(\data_in_frame[7] [6]), .O(n35167));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1436 (.I0(n16660), .I1(n16530), .I2(\data_out_frame[13] [5]), 
            .I3(GND_net), .O(n14_adj_4494));
    defparam i5_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1437 (.I0(n30859), .I1(\data_in_frame[21] [7]), 
            .I2(n34849), .I3(\data_in_frame[21] [6]), .O(n12_adj_4495));
    defparam i3_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1438 (.I0(n34948), .I1(\data_out_frame[18][0] ), 
            .I2(n16713), .I3(\data_out_frame[7] [2]), .O(n15_adj_4496));
    defparam i6_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1439 (.I0(n15_adj_4496), .I1(n16634), .I2(n14_adj_4494), 
            .I3(n16851), .O(n30432));
    defparam i8_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1440 (.I0(Kp_23__N_1783), .I1(n12_adj_4495), .I2(n30549), 
            .I3(Kp_23__N_731), .O(n15_adj_4497));
    defparam i6_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1441 (.I0(\data_out_frame[18][1] ), .I1(n30432), 
            .I2(GND_net), .I3(GND_net), .O(n35009));
    defparam i1_2_lut_adj_1441.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4498));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1443 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[6] [5]), .I3(n6_adj_4498), .O(n16370));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1444 (.I0(n16526), .I1(n16370), .I2(\data_out_frame[12] [7]), 
            .I3(\data_out_frame[10] [5]), .O(n10_adj_4452));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1445 (.I0(\data_out_frame[15] [3]), .I1(n34937), 
            .I2(GND_net), .I3(GND_net), .O(n16029));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1445.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34759));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1447 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16634));
    defparam i1_2_lut_adj_1447.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1448 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16875));
    defparam i1_2_lut_adj_1448.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1449 (.I0(\data_out_frame[13] [4]), .I1(n34759), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[15] [6]), .O(n16713));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1450 (.I0(n16713), .I1(n16376), .I2(\data_out_frame[16] [0]), 
            .I3(\data_out_frame[18]_c [2]), .O(n12_adj_4499));
    defparam i5_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1451 (.I0(\data_in_frame[24] [3]), .I1(\data_in_frame[22] [1]), 
            .I2(n34849), .I3(GND_net), .O(n8_adj_4500));
    defparam i3_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1452 (.I0(\data_out_frame[13] [7]), .I1(n12_adj_4499), 
            .I2(n35164), .I3(n16404), .O(n34755));
    defparam i6_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1453 (.I0(n15_adj_4497), .I1(n35251), .I2(n14_adj_4454), 
            .I3(n35269), .O(n37062));
    defparam i8_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16130));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1455 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16530));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1455.LUT_INIT = 16'h6666;
    SB_LUT4 i532_2_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1336));   // verilog/coms.v(69[16:27])
    defparam i532_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1456 (.I0(n16124), .I1(n16526), .I2(\data_out_frame[10] [5]), 
            .I3(GND_net), .O(n34812));
    defparam i2_3_lut_adj_1456.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_21__7__I_0_3518_rep_147_2_lut (.I0(\data_in_frame[21] [7]), 
            .I1(\data_in_frame[21] [6]), .I2(GND_net), .I3(GND_net), .O(n43807));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_21__7__I_0_3518_rep_147_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1457 (.I0(\data_in_frame[22] [7]), .I1(n16610), 
            .I2(\data_in_frame[18] [6]), .I3(n35091), .O(n10_adj_4501));
    defparam i4_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1458 (.I0(\data_in_frame[24] [2]), .I1(n34831), 
            .I2(n43807), .I3(\data_in_frame[22] [1]), .O(n37063));
    defparam i3_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1459 (.I0(n34812), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n34824));
    defparam i2_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1460 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16851));
    defparam i1_2_lut_adj_1460.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16753));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1462 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [2]), .I3(n6_adj_4451), .O(n35151));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1463 (.I0(n34852), .I1(n37090), .I2(\data_in_frame[20] [4]), 
            .I3(\data_in_frame[24] [6]), .O(n14_adj_4502));
    defparam i6_4_lut_adj_1463.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1464 (.I0(\data_in_frame[22] [2]), .I1(n30859), 
            .I2(\data_in_frame[22] [3]), .I3(n34849), .O(n4_adj_4503));
    defparam i1_4_lut_adj_1464.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1465 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n34821));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16839));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1467 (.I0(\data_in_frame[22] [5]), .I1(n31320), 
            .I2(n16414), .I3(\data_in_frame[22] [4]), .O(n13_adj_4504));
    defparam i5_4_lut_adj_1467.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34768));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1469 (.I0(\data_in_frame[12] [4]), .I1(n30481), 
            .I2(n10_adj_4437), .I3(n31439), .O(n30625));
    defparam i5_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1470 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[8] [3]), 
            .I2(n34768), .I3(n6_adj_4300), .O(n15974));
    defparam i4_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1471 (.I0(n15974), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16401));
    defparam i1_2_lut_adj_1471.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n41_adj_4362));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h5454;
    SB_LUT4 i1_4_lut_adj_1473 (.I0(n16631), .I1(n35182), .I2(n36905), 
            .I3(n31386), .O(n6_adj_4505));
    defparam i1_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1474 (.I0(\data_out_frame[6] [7]), .I1(n16482), 
            .I2(n16742), .I3(n16401), .O(n34762));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1475 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16526));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1476 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n35154));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_adj_1477 (.I0(n34762), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42_adj_4506));   // verilog/coms.v(71[16:27])
    defparam i4_2_lut_adj_1477.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[11] [7]), .I1(n34927), .I2(n16839), 
            .I3(n34821), .O(n60));   // verilog/coms.v(71[16:27])
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1478 (.I0(n31302), .I1(n35151), .I2(n34815), 
            .I3(\data_out_frame[9] [2]), .O(n58));   // verilog/coms.v(71[16:27])
    defparam i20_4_lut_adj_1478.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1479 (.I0(\data_in_frame[22] [5]), .I1(n30549), 
            .I2(\data_in_frame[22] [6]), .I3(GND_net), .O(n4_adj_4507));   // verilog/coms.v(83[17:28])
    defparam i1_3_lut_adj_1479.LUT_INIT = 16'h9696;
    SB_LUT4 i30_4_lut (.I0(n16851), .I1(n60), .I2(n42_adj_4506), .I3(n34824), 
            .O(n68));   // verilog/coms.v(71[16:27])
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut_adj_1480 (.I0(\data_out_frame[5] [4]), .I1(n16499), 
            .I2(n16526), .I3(\data_out_frame[6] [4]), .O(n64));   // verilog/coms.v(71[16:27])
    defparam i26_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1481 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[11] [3]), .I3(n16276), .O(n62));   // verilog/coms.v(71[16:27])
    defparam i24_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1482 (.I0(n25_adj_4476), .I1(n27_adj_4474), .I2(n26_adj_4473), 
            .I3(n28_adj_4471), .O(n36809));
    defparam i15_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1483 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [3]), 
            .I2(n34842), .I3(n34911), .O(n63_adj_4508));   // verilog/coms.v(71[16:27])
    defparam i25_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1484 (.I0(n34803), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[9] [3]), .I3(n16020), .O(n61));   // verilog/coms.v(71[16:27])
    defparam i23_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n16072), .I1(\data_out_frame[6] [7]), .I2(\data_out_frame[6] [6]), 
            .I3(n15886), .O(n66));   // verilog/coms.v(71[16:27])
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34_4_lut (.I0(n16124), .I1(n68), .I2(n58), .I3(\data_out_frame[8] [0]), 
            .O(n72));   // verilog/coms.v(71[16:27])
    defparam i34_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31330_4_lut (.I0(\data_in_frame[24] [4]), .I1(n13_adj_4504), 
            .I2(n4_adj_4503), .I3(n14_adj_4502), .O(n38096));
    defparam i31330_4_lut.LUT_INIT = 16'h1248;
    SB_LUT4 i6_4_lut_adj_1485 (.I0(\data_in_frame[19] [2]), .I1(n12_adj_4478), 
            .I2(n35200), .I3(\data_in_frame[21] [2]), .O(n36304));
    defparam i6_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1486 (.I0(\data_in_frame[24] [5]), .I1(n36985), 
            .I2(n8_adj_4482), .I3(\data_in_frame[22] [4]), .O(n22));
    defparam i6_4_lut_adj_1486.LUT_INIT = 16'hedde;
    SB_LUT4 i27_4_lut_adj_1487 (.I0(\data_out_frame[8] [2]), .I1(n34768), 
            .I2(n16016), .I3(\data_out_frame[6] [5]), .O(n65));   // verilog/coms.v(71[16:27])
    defparam i27_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n61), .I1(n63_adj_4508), .I2(n62), .I3(n64), 
            .O(n73));   // verilog/coms.v(71[16:27])
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i37_4_lut (.I0(n73), .I1(n65), .I2(n72), .I3(n66), .O(n30424));   // verilog/coms.v(71[16:27])
    defparam i37_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31353_4_lut (.I0(n38096), .I1(n36809), .I2(\data_in_frame[24] [7]), 
            .I3(n4_adj_4507), .O(n38120));
    defparam i31353_4_lut.LUT_INIT = 16'h0880;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35254));
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[13] [0]), 
            .I2(Kp_23__N_1186), .I3(GND_net), .O(n6_adj_4435));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1490 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[15] [1]), .I3(GND_net), .O(n34924));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1490.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(\data_in_frame[10] [6]), .I1(Kp_23__N_1183), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n35134));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16760));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1493 (.I0(\data_in_frame[23] [6]), .I1(n16570), 
            .I2(n35048), .I3(n6_adj_4505), .O(n36959));
    defparam i4_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(\data_in_frame[24] [0]), .I1(n34831), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4509));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1495 (.I0(n31094), .I1(n34974), .I2(n35094), 
            .I3(\data_in_frame[11] [3]), .O(n35045));
    defparam i2_3_lut_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1496 (.I0(\data_in_frame[11] [5]), .I1(n31368), 
            .I2(n36645), .I3(GND_net), .O(n35094));
    defparam i1_2_lut_3_lut_adj_1496.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1497 (.I0(\data_out_frame[12] [4]), .I1(n35263), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n34815));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1497.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1498 (.I0(n34815), .I1(n35215), .I2(\data_out_frame[12] [3]), 
            .I3(GND_net), .O(n16060));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1498.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1499 (.I0(n11), .I1(n34775), .I2(n30859), .I3(n34849), 
            .O(n14_adj_4510));
    defparam i6_4_lut_adj_1499.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1500 (.I0(n15_adj_4486), .I1(\data_in_frame[16] [6]), 
            .I2(n14_adj_4484), .I3(n31320), .O(n36997));
    defparam i8_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1501 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [6]), 
            .I2(n16430), .I3(\data_in_frame[6] [1]), .O(n10_adj_4405));   // verilog/coms.v(69[16:62])
    defparam i2_2_lut_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1502 (.I0(\data_out_frame[10] [3]), .I1(n15489), 
            .I2(n16060), .I3(GND_net), .O(n30545));
    defparam i2_3_lut_adj_1502.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16736));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1504 (.I0(\data_in_frame[17] [0]), .I1(n36936), 
            .I2(n10_adj_4491), .I3(n35785), .O(n18_adj_4511));
    defparam i2_4_lut_adj_1504.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35078));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1506 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(n10_adj_4402), .I3(n31392), .O(n34974));
    defparam i5_3_lut_4_lut_adj_1506.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1507 (.I0(n9_adj_4509), .I1(n16160), .I2(\data_in_frame[20] [4]), 
            .I3(n37090), .O(n13_adj_4512));
    defparam i5_4_lut_adj_1507.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16593));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1509 (.I0(\data_in_frame[22] [2]), .I1(n37062), 
            .I2(n8_adj_4500), .I3(n30861), .O(n20_adj_4513));
    defparam i4_4_lut_adj_1509.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_2_lut_3_lut_adj_1510 (.I0(\data_in_frame[9] [0]), .I1(n16716), 
            .I2(\data_in_frame[8] [7]), .I3(GND_net), .O(n35137));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1510.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1511 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(n34874), .I3(GND_net), .O(Kp_23__N_1189));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1511.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1512 (.I0(\data_out_frame[15] [2]), .I1(n34790), 
            .I2(n35203), .I3(n16593), .O(n32_adj_4514));
    defparam i12_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1513 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [4]), 
            .I2(n34948), .I3(\data_out_frame[14] [4]), .O(n31_adj_4515));
    defparam i11_4_lut_adj_1513.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1514 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [5]), 
            .I2(n16736), .I3(n30545), .O(n35));
    defparam i15_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i31332_4_lut (.I0(\data_in_frame[20] [5]), .I1(n37063), .I2(n10_adj_4501), 
            .I3(\data_in_frame[23] [1]), .O(n38098));
    defparam i31332_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i14_4_lut_adj_1515 (.I0(n36959), .I1(n38120), .I2(n22), .I3(n36304), 
            .O(n30));
    defparam i14_4_lut_adj_1515.LUT_INIT = 16'hfff7;
    SB_LUT4 i9_4_lut_adj_1516 (.I0(n13_adj_4512), .I1(n18_adj_4511), .I2(n36997), 
            .I3(n14_adj_4510), .O(n25_adj_4516));
    defparam i9_4_lut_adj_1516.LUT_INIT = 16'hefdf;
    SB_LUT4 i15_4_lut_adj_1517 (.I0(n25_adj_4516), .I1(n30), .I2(n38098), 
            .I3(n20_adj_4513), .O(n31));
    defparam i15_4_lut_adj_1517.LUT_INIT = 16'hffef;
    SB_LUT4 i14_4_lut_adj_1518 (.I0(n34924), .I1(\data_out_frame[14] [0]), 
            .I2(\data_out_frame[14] [3]), .I3(n16299), .O(n34_adj_4517));
    defparam i14_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i18_3_lut (.I0(n35), .I1(n31_adj_4515), .I2(n32_adj_4514), 
            .I3(GND_net), .O(n38_adj_4518));
    defparam i18_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4519));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[15] [7]), .I1(n35254), .I2(n30424), 
            .I3(n35154), .O(n33));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13094_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n17823));
    defparam i13094_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13095_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n17824));
    defparam i13095_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13183_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n17912));
    defparam i13183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1520 (.I0(n33), .I1(n6_adj_4519), .I2(n38_adj_4518), 
            .I3(n34_adj_4517), .O(n8_adj_4520));
    defparam i3_4_lut_adj_1520.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1521 (.I0(\data_out_frame[16] [1]), .I1(n16530), 
            .I2(n8_adj_4520), .I3(\data_out_frame[16] [2]), .O(n6_adj_4521));
    defparam i1_4_lut_adj_1521.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1522 (.I0(\data_out_frame[17] [1]), .I1(n16130), 
            .I2(\data_out_frame[17] [2]), .I3(n6_adj_4521), .O(n35042));
    defparam i4_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1523 (.I0(n16354), .I1(\data_in_frame[4] [4]), 
            .I2(n34749), .I3(GND_net), .O(n34874));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1524 (.I0(n35215), .I1(n35236), .I2(\data_out_frame[14] [3]), 
            .I3(n16103), .O(n12_adj_4522));   // verilog/coms.v(70[16:41])
    defparam i5_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1525 (.I0(\data_out_frame[12] [2]), .I1(n12_adj_4522), 
            .I2(n35263), .I3(\data_out_frame[12] [1]), .O(n16212));   // verilog/coms.v(70[16:41])
    defparam i6_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1526 (.I0(n16212), .I1(\data_out_frame[17] [0]), 
            .I2(n31381), .I3(n35042), .O(n10_adj_4301));
    defparam i4_4_lut_adj_1526.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1527 (.I0(n16530), .I1(\data_out_frame[18] [7]), 
            .I2(n34755), .I3(n16593), .O(n16_adj_4523));
    defparam i6_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(n36954), .I1(n16_adj_4523), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n18_adj_4524));
    defparam i8_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i7_4_lut_adj_1528 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(n35009), .I3(\data_out_frame[18] [3]), .O(n17_adj_4525));
    defparam i7_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i13182_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n17911));
    defparam i13182_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1529 (.I0(\data_out_frame[16] [0]), .I1(n35100), 
            .I2(n34991), .I3(n16212), .O(n37123));
    defparam i3_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i13096_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n17825));
    defparam i13096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1530 (.I0(n37123), .I1(n16886), .I2(n17_adj_4525), 
            .I3(n18_adj_4524), .O(n19260));
    defparam i11_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i13185_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n17914));
    defparam i13185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1531 (.I0(n19260), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4526));
    defparam i2_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1532 (.I0(n7_adj_4526), .I1(n31421), .I2(n31435), 
            .I3(n36296), .O(n36413));
    defparam i4_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i13097_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n17826));
    defparam i13097_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13098_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n17827));
    defparam i13098_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13184_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n17913));
    defparam i13184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13187_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n17916));
    defparam i13187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13186_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n17915));
    defparam i13186_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1533 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15886));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1533.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16020));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1535 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35111));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35218));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i13099_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n17828));
    defparam i13099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13189_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n17918));
    defparam i13189_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13188_3_lut_4_lut (.I0(n8_adj_4375), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n17917));
    defparam i13188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1537 (.I0(\data_out_frame[10] [0]), .I1(n35218), 
            .I2(n35111), .I3(n34930), .O(n16699));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1538 (.I0(\data_out_frame[10] [2]), .I1(n16312), 
            .I2(\data_out_frame[5] [7]), .I3(n6_adj_4448), .O(n30994));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1539 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34803));
    defparam i1_2_lut_adj_1539.LUT_INIT = 16'h6666;
    SB_LUT4 i13100_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n17829));
    defparam i13100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(n30994), .I1(n16699), .I2(GND_net), 
            .I3(GND_net), .O(n31302));
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1541 (.I0(n31030), .I1(n35094), .I2(\data_in_frame[11] [3]), 
            .I3(n35185), .O(n31310));
    defparam i1_2_lut_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i909_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1713));   // verilog/coms.v(83[17:28])
    defparam i909_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1542 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[10] [2]), .I3(n6_adj_4441), .O(n14_adj_4391));
    defparam i5_3_lut_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1543 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n34842));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1543.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1544 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16016));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1544.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1545 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16072));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i13177_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n17906));
    defparam i13177_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1546 (.I0(n16016), .I1(n34842), .I2(\data_out_frame[9] [5]), 
            .I3(GND_net), .O(n16103));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i13176_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n17905));
    defparam i13176_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13101_3_lut_4_lut (.I0(n8_adj_4364), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n17830));
    defparam i13101_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1547 (.I0(n16103), .I1(n16482), .I2(\data_out_frame[9] [4]), 
            .I3(GND_net), .O(n34793));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1548 (.I0(\data_out_frame[7] [2]), .I1(n34793), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n16417));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1548.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16276));
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1550 (.I0(\data_out_frame[6] [6]), .I1(n34934), 
            .I2(GND_net), .I3(GND_net), .O(n16794));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1550.LUT_INIT = 16'h6666;
    SB_LUT4 i13175_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n17904));
    defparam i13175_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13179_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n17908));
    defparam i13179_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1551 (.I0(\data_out_frame[18] [4]), .I1(n35164), 
            .I2(\data_out_frame[6] [7]), .I3(n16794), .O(n10_adj_4293));
    defparam i4_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i13178_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n17907));
    defparam i13178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1552 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(n37031), .I3(\data_in_frame[18] [4]), .O(n35029));
    defparam i2_3_lut_4_lut_adj_1552.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1553 (.I0(n31302), .I1(n34803), .I2(\data_out_frame[14] [4]), 
            .I3(GND_net), .O(n31414));
    defparam i2_3_lut_adj_1553.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1554 (.I0(n14249), .I1(\data_in_frame[16] [0]), 
            .I2(n37090), .I3(GND_net), .O(n35038));
    defparam i1_2_lut_3_lut_adj_1554.LUT_INIT = 16'h6969;
    SB_LUT4 i13181_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n17910));
    defparam i13181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1555 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n34782));
    defparam i2_3_lut_adj_1555.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16324));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(\data_out_frame[20] [7]), .I1(n35100), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4527));
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1558 (.I0(n16324), .I1(\data_out_frame[18] [6]), 
            .I2(n34782), .I3(n6_adj_4527), .O(n37121));
    defparam i4_4_lut_adj_1558.LUT_INIT = 16'h9669;
    SB_LUT4 i13180_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n17909));
    defparam i13180_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1559 (.I0(n14249), .I1(\data_in_frame[16] [0]), 
            .I2(n10_adj_4383), .I3(n31006), .O(n30859));
    defparam i5_3_lut_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1560 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[17] [4]), 
            .I2(n36773), .I3(GND_net), .O(n10_adj_4381));
    defparam i2_2_lut_3_lut_adj_1560.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1561 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[20] [0]), 
            .I2(n16537), .I3(n36773), .O(n35131));
    defparam i2_3_lut_4_lut_adj_1561.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36343 (.I0(\byte_transmit_counter[1] ), 
            .I1(n38255), .I2(n38256), .I3(byte_transmit_counter[2]), .O(n43166));
    defparam byte_transmit_counter_1__bdd_4_lut_36343.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1562 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n35122));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1562.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1563 (.I0(\FRAME_MATCHER.state [3]), .I1(n34603), 
            .I2(n27212), .I3(GND_net), .O(n19503));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_adj_1563.LUT_INIT = 16'hfefe;
    SB_LUT4 i13174_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n17903));
    defparam i13174_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13142_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n17871));
    defparam i13142_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1564 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[15] [7]), .I3(\data_in_frame[15] [6]), .O(n7_adj_4386));
    defparam i2_2_lut_3_lut_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i13076_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n17805));
    defparam i13076_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n43166_bdd_4_lut (.I0(n43166), .I1(n38253), .I2(n38252), .I3(byte_transmit_counter[2]), 
            .O(n43169));
    defparam n43166_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13077_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n17806));
    defparam i13077_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13070_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n17799));
    defparam i13070_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1565 (.I0(n29), .I1(n27212), .I2(n34603), .I3(n6_adj_4449), 
            .O(n36881));
    defparam i4_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i13071_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n17800));
    defparam i13071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13072_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n17801));
    defparam i13072_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13073_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n17802));
    defparam i13073_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13143_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n17872));
    defparam i13143_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13074_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n17803));
    defparam i13074_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13075_3_lut_4_lut (.I0(n24351), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n17804));
    defparam i13075_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19015_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15648), .I3(\FRAME_MATCHER.i [31]), .O(n2957));
    defparam i19015_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 equal_110_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4263));
    defparam equal_110_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i19625_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24351));
    defparam i19625_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13144_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n17873));
    defparam i13144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13062_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n17791));
    defparam i13062_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13063_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n17792));
    defparam i13063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13145_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n17874));
    defparam i13145_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13064_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n17793));
    defparam i13064_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13065_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n17794));
    defparam i13065_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13146_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n17875));
    defparam i13146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13066_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n17795));
    defparam i13066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13067_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n17796));
    defparam i13067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13147_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n17876));
    defparam i13147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13068_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n17797));
    defparam i13068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_107_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_4283));   // verilog/coms.v(151[7:23])
    defparam equal_107_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1566 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [7]), .O(n35215));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1566.LUT_INIT = 16'h6996;
    SB_LUT4 i13148_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n17877));
    defparam i13148_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1567 (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4296), 
            .I2(n63_adj_4292), .I3(n63_adj_4285), .O(\FRAME_MATCHER.state_31__N_2661[2] ));   // verilog/coms.v(141[7:84])
    defparam i1_2_lut_4_lut_adj_1567.LUT_INIT = 16'hb300;
    SB_LUT4 i13069_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n17798));
    defparam i13069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1568 (.I0(tx_transmit_N_3479), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3582[0]), .I3(GND_net), .O(n1211));   // verilog/coms.v(206[11:56])
    defparam i1_2_lut_3_lut_adj_1568.LUT_INIT = 16'hfefe;
    SB_LUT4 i19884_3_lut_4_lut (.I0(\byte_transmit_counter[1] ), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[3]), 
            .O(n24610));
    defparam i19884_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_4_lut_adj_1569 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n15731), .I3(\FRAME_MATCHER.i [2]), .O(n4_adj_4284));
    defparam i1_2_lut_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i13149_3_lut_4_lut (.I0(n10_adj_4378), .I1(n34697), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n17878));
    defparam i13149_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1570 (.I0(\FRAME_MATCHER.state [0]), .I1(n19503), 
            .I2(n31), .I3(GND_net), .O(n5_adj_4281));   // verilog/coms.v(126[12] 292[6])
    defparam i1_2_lut_3_lut_adj_1570.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38191), .I3(n43205), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_4_lut_adj_1571 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(n31129), .O(n34978));
    defparam i1_2_lut_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1572 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n14136));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1572.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38221), .I3(n38220), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_3_lut_adj_1573 (.I0(n16427), .I1(n6_adj_4363), .I2(n34749), 
            .I3(GND_net), .O(n16430));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 equal_1183_i15_2_lut_3_lut (.I0(n16427), .I1(n6_adj_4363), .I2(\data_in_frame[4] [6]), 
            .I3(GND_net), .O(n15_adj_4401));   // verilog/coms.v(74[16:43])
    defparam equal_1183_i15_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1574 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2][2] ), 
            .I2(\data_in_frame[4] [3]), .I3(GND_net), .O(n34864));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_3_lut_adj_1574.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1575 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2][2] ), 
            .I2(\data_in_frame[0] [0]), .I3(n4_c), .O(n34749));   // verilog/coms.v(163[9:87])
    defparam i2_3_lut_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i13197_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n17926));
    defparam i13197_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13196_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n17925));
    defparam i13196_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13195_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n17924));
    defparam i13195_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13194_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n17923));
    defparam i13194_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13193_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n17922));
    defparam i13193_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13192_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n17921));
    defparam i13192_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13191_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n17920));
    defparam i13191_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13190_3_lut_4_lut (.I0(n8_adj_4263), .I1(n34715), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n17919));
    defparam i13190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1576 (.I0(n34900), .I1(n34978), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n1));
    defparam i1_2_lut_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n6));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38218), .I3(n38217), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_4_lut_adj_1578 (.I0(\data_in_frame[2]_c [1]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[2][0] ), .I3(n35082), .O(n16354));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1579 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(n34806), .I3(GND_net), .O(n6_adj_4441));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1579.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38215), .I3(n38214), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13046_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n17775));
    defparam i13046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13047_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n17776));
    defparam i13047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13048_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n17777));
    defparam i13048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13049_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n17778));
    defparam i13049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38212), .I3(n38211), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_1055_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2]_c [1]), 
            .I2(n4348), .I3(GND_net), .O(n4358));
    defparam mux_1055_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38203), .I3(n43181), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13050_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n17779));
    defparam i13050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19665_3_lut_4_lut (.I0(n63), .I1(n15876), .I2(tx_active), 
            .I3(r_SM_Main_2__N_3582[0]), .O(n24391));
    defparam i19665_3_lut_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i2_3_lut_4_lut_adj_1580 (.I0(\FRAME_MATCHER.state [3]), .I1(n34603), 
            .I2(n27212), .I3(n81), .O(n63));   // verilog/coms.v(126[12] 292[6])
    defparam i2_3_lut_4_lut_adj_1580.LUT_INIT = 16'hfffd;
    SB_LUT4 i13051_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n17780));
    defparam i13051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13052_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n17781));
    defparam i13052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13053_3_lut_4_lut (.I0(n8_adj_4376), .I1(n34707), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n17782));
    defparam i13053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13102_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n17831));
    defparam i13102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38206), .I3(n43175), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38209), .I3(n43169), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1581 (.I0(n16299), .I1(\data_out_frame[6] [6]), 
            .I2(n34934), .I3(n35203), .O(n15422));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1582 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[8] [0]), .O(n35263));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_3_lut_4_lut_adj_1582.LUT_INIT = 16'h6996;
    SB_LUT4 i13103_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n17832));
    defparam i13103_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13104_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n17833));
    defparam i13104_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13105_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n17834));
    defparam i13105_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13106_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n17835));
    defparam i13106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13107_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n17836));
    defparam i13107_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13108_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n17837));
    defparam i13108_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13109_3_lut_4_lut (.I0(n8), .I1(n34723), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n17838));
    defparam i13109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1583 (.I0(n34603), .I1(n27212), .I2(n34683), 
            .I3(\FRAME_MATCHER.state [3]), .O(n13263));
    defparam i2_3_lut_4_lut_adj_1583.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_4_lut_adj_1584 (.I0(n34603), .I1(n27212), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(\FRAME_MATCHER.state [2]), .O(n24684));
    defparam i1_2_lut_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    uart_tx tx (.clk32MHz(clk32MHz), .n17314(n17314), .r_Bit_Index({r_Bit_Index}), 
            .n17311(n17311), .r_SM_Main({r_SM_Main}), .tx_data({tx_data}), 
            .GND_net(GND_net), .n17446(n17446), .n17412(n17412), .n17411(n17411), 
            .tx_active(tx_active), .n17410(n17410), .tx_o(tx_o), .VCC_net(VCC_net), 
            .\r_SM_Main_2__N_3582[0] (r_SM_Main_2__N_3582[0]), .\r_SM_Main_2__N_3579[1] (\r_SM_Main_2__N_3579[1] ), 
            .n17058(n17058), .n43694(n43694), .n4670(n4670), .n17189(n17189), 
            .n4(n4), .n3(n3), .n8936(n8936), .n10627(n10627), .tx_enable(tx_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n17338(n17338), .r_Bit_Index({r_Bit_Index_adj_11}), 
            .n17341(n17341), .n24450(n24450), .r_SM_Main({\r_SM_Main[2]_adj_7 , 
            \r_SM_Main[1]_adj_6 , Open_10}), .r_Rx_Data(r_Rx_Data), .PIN_13_N_105(PIN_13_N_105), 
            .GND_net(GND_net), .n40218(n40218), .n40217(n40217), .n17452(n17452), 
            .rx_data_ready(rx_data_ready), .n17462(n17462), .rx_data({rx_data}), 
            .n4(n4_adj_8), .n17429(n17429), .n17428(n17428), .n17427(n17427), 
            .n17426(n17426), .n17425(n17425), .n17403(n17403), .n17052(n17052), 
            .n17180(n17180), .n4648(n4648), .n17343(n17343), .n17342(n17342), 
            .VCC_net(VCC_net), .n43211(n43211), .n15734(n15734), .n15626(n15626), 
            .n23653(n23653), .n4_adj_1(n4_adj_9), .n4_adj_2(n4_adj_10)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, n17314, r_Bit_Index, n17311, r_SM_Main, 
            tx_data, GND_net, n17446, n17412, n17411, tx_active, 
            n17410, tx_o, VCC_net, \r_SM_Main_2__N_3582[0] , \r_SM_Main_2__N_3579[1] , 
            n17058, n43694, n4670, n17189, n4, n3, n8936, n10627, 
            tx_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n17314;
    output [2:0]r_Bit_Index;
    input n17311;
    output [2:0]r_SM_Main;
    input [7:0]tx_data;
    input GND_net;
    input n17446;
    input n17412;
    input n17411;
    output tx_active;
    input n17410;
    output tx_o;
    input VCC_net;
    input \r_SM_Main_2__N_3582[0] ;
    output \r_SM_Main_2__N_3579[1] ;
    output n17058;
    input n43694;
    output n4670;
    output n17189;
    output n4;
    output n3;
    output n8936;
    output n10627;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n17298;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n17295, n17292, n56, n17286, n17307, n17304, n17301, 
        n18035, n13253;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n26497, n17284, n17287, n17290, n17293, n10, n29969, 
        n38100, n63, n17296, n17443, n17441, n27869, n27868, n27867, 
        n27866, n27865, n17299, n27864, n17302, n27863, n17305, 
        n27862, n24134, n43214, n43217, n43190, n43193, o_Tx_Serial_N_3610;
    
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n17298));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n17295));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n17292));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n56));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n17286));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17314));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17311));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n17307));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17304));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n17301));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n18035));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut (.I0(n26497), .I1(n17284), .I2(GND_net), .I3(GND_net), 
            .O(n17286));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_994 (.I0(n26497), .I1(n17287), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_995 (.I0(n26497), .I1(n17290), .I2(GND_net), 
            .I3(GND_net), .O(n17292));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_996 (.I0(n26497), .I1(n17293), .I2(GND_net), 
            .I3(GND_net), .O(n17295));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[5]), 
            .I3(r_Clock_Count[1]), .O(n10));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[4]), .I1(n10), .I2(r_Clock_Count[3]), 
            .I3(GND_net), .O(n29969));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i31334_3_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[8]), 
            .I2(n29969), .I3(GND_net), .O(n38100));
    defparam i31334_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_997 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n63));   // verilog/uart_tx.v(31[16:25])
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n63), .I2(n38100), .I3(r_Clock_Count[7]), 
            .O(n26497));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut.LUT_INIT = 16'haaae;
    SB_LUT4 i1_2_lut_adj_998 (.I0(n26497), .I1(n17296), .I2(GND_net), 
            .I3(GND_net), .O(n17298));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h8888;
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n17443));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17446));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut_adj_999 (.I0(n26497), .I1(n17441), .I2(GND_net), 
            .I3(GND_net), .O(n17443));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h8888;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n17412));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n17411));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n17410));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13253), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[8]), 
            .I2(r_SM_Main[2]), .I3(n27869), .O(n17284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_59_9_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[7]), 
            .I2(r_SM_Main[2]), .I3(n27868), .O(n17287)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_9 (.CI(n27868), .I0(r_Clock_Count[7]), .I1(r_SM_Main[2]), 
            .CO(n27869));
    SB_LUT4 add_59_8_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[6]), 
            .I2(r_SM_Main[2]), .I3(n27867), .O(n17290)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_8 (.CI(n27867), .I0(r_Clock_Count[6]), .I1(r_SM_Main[2]), 
            .CO(n27868));
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(r_SM_Main[2]), .I3(n27866), .O(n17293)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n27866), .I0(r_Clock_Count[5]), .I1(r_SM_Main[2]), 
            .CO(n27867));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(r_SM_Main[2]), .I3(n27865), .O(n17296)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n27865), .I0(r_Clock_Count[4]), .I1(r_SM_Main[2]), 
            .CO(n27866));
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(r_SM_Main[2]), .I3(n27864), .O(n17299)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_5 (.CI(n27864), .I0(r_Clock_Count[3]), .I1(r_SM_Main[2]), 
            .CO(n27865));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(r_SM_Main[2]), .I3(n27863), .O(n17302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n27863), .I0(r_Clock_Count[2]), .I1(r_SM_Main[2]), 
            .CO(n27864));
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(r_SM_Main[2]), .I3(n27862), .O(n17305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n27862), .I0(r_Clock_Count[1]), .I1(r_SM_Main[2]), 
            .CO(n27863));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(r_SM_Main[2]), .I3(VCC_net), .O(n17441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(r_SM_Main[2]), 
            .CO(n27862));
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3582[0] ), 
            .I3(r_SM_Main[1]), .O(n13253));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3579[1] ), .O(n17058));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n43694));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut_adj_1000 (.I0(n26497), .I1(n17299), .I2(GND_net), 
            .I3(GND_net), .O(n17301));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(n26497), .I1(n17302), .I2(GND_net), 
            .I3(GND_net), .O(n17304));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(n26497), .I1(n17305), .I2(GND_net), 
            .I3(GND_net), .O(n17307));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h8888;
    SB_LUT4 i1299_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4670));   // verilog/uart_tx.v(98[36:51])
    defparam i1299_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24134));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n29969), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3579[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12460_3_lut (.I0(n17058), .I1(n24134), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17189));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12460_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n43214));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43214_bdd_4_lut (.I0(n43214), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n43217));
    defparam n43214_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_36376 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n43190));
    defparam r_Bit_Index_0__bdd_4_lut_36376.LUT_INIT = 16'he4aa;
    SB_LUT4 n43190_bdd_4_lut (.I0(n43190), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n43193));
    defparam n43190_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1003 (.I0(\r_SM_Main_2__N_3579[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_adj_1003.LUT_INIT = 16'h008f;
    SB_LUT4 i13306_3_lut_4_lut (.I0(\r_SM_Main_2__N_3579[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n18035));
    defparam i13306_3_lut_4_lut.LUT_INIT = 16'h0078;
    SB_LUT4 i1999836_i1_3_lut (.I0(n43193), .I1(n43217), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3610));
    defparam i1999836_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3610), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i4284_2_lut (.I0(\r_SM_Main_2__N_3582[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n8936));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i4284_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5955_4_lut (.I0(\r_SM_Main_2__N_3582[0] ), .I1(n24134), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3579[1] ), .O(n10627));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5955_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n17338, r_Bit_Index, n17341, n24450, r_SM_Main, 
            r_Rx_Data, PIN_13_N_105, GND_net, n40218, n40217, n17452, 
            rx_data_ready, n17462, rx_data, n4, n17429, n17428, 
            n17427, n17426, n17425, n17403, n17052, n17180, n4648, 
            n17343, n17342, VCC_net, n43211, n15734, n15626, n23653, 
            n4_adj_1, n4_adj_2) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n17338;
    output [2:0]r_Bit_Index;
    input n17341;
    input n24450;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input PIN_13_N_105;
    input GND_net;
    output n40218;
    output n40217;
    input n17452;
    output rx_data_ready;
    input n17462;
    output [7:0]rx_data;
    output n4;
    input n17429;
    input n17428;
    input n17427;
    input n17426;
    input n17425;
    input n17403;
    output n17052;
    output n17180;
    output n4648;
    input n17343;
    input n17342;
    input VCC_net;
    output n43211;
    output n15734;
    output n15626;
    output n23653;
    output n4_adj_1;
    output n4_adj_2;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n17274;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n45, n17268, n17265, n17283, n17280, n17277, n35310, 
        r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3508;
    
    wire n34673;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n34702, n34731, n24382, n37230, n19380, n36891, n34657, 
        n6, n19399, n6_adj_4254, n2588;
    wire [31:0]n194;
    
    wire n34271, n24484, n16980, n27861, n27860, n27859, n27858, 
        n27857, n27856, n27855, n40176, n43208;
    
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n17274));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n45));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n17268));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n17265));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n17283));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17280));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n17277));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17338));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17341));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n24450));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n35310));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3508[2]), 
            .R(n34673));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n34702));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_989 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n34731));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut (.I0(n24382), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[5]), .O(n37230));
    defparam i3_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2_4_lut (.I0(n19380), .I1(n34731), .I2(r_Clock_Count[5]), 
            .I3(n24382), .O(n36891));
    defparam i2_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut (.I0(n36891), .I1(n37230), .I2(n34702), .I3(r_SM_Main[2]), 
            .O(n34657));
    defparam i1_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_adj_990 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19380));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_990.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_991 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[2]), 
            .I3(n6), .O(n24382));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_2_lut (.I0(n19399), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4254));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_992 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4254), 
            .I3(r_Rx_Data), .O(n2588));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hbaaa;
    SB_LUT4 i28549_4_lut (.I0(r_Clock_Count[0]), .I1(n194[0]), .I2(n2588), 
            .I3(n34657), .O(n35310));
    defparam i28549_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i33764_2_lut (.I0(r_SM_Main_2__N_3508[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n40218));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33764_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33807_3_lut (.I0(r_SM_Main_c[0]), .I1(n19399), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n40217));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33807_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17452));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n34271));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n17462));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_139_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_139_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17429));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17428));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17427));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17426));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17425));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n17403));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24484));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i12451_3_lut (.I0(n17052), .I1(r_SM_Main[1]), .I2(n24484), 
            .I3(GND_net), .O(n17180));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12451_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1277_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4648));   // verilog/uart_rx.v(102[36:51])
    defparam i1277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3508[2]), 
            .I3(r_SM_Main_c[0]), .O(n16980));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n16980), 
            .I3(rx_data_ready), .O(n34271));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i36282_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_c[0]), 
            .I3(GND_net), .O(n34673));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36282_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17343));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17342));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n27861), .O(n194[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n27860), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n27860), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n27861));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n27859), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n27859), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n27860));
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n27858), .O(n194[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_6 (.CI(n27858), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n27859));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n27857), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n27857), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n27858));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27856), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n27856), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27857));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27855), .O(n194[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n27855), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27856));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n27855));
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(r_SM_Main_2__N_3508[2]), .I1(r_SM_Main[1]), 
            .I2(n40176), .I3(r_SM_Main_c[0]), .O(n43208));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 n43208_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n19399), 
            .I3(n43208), .O(n43211));   // verilog/uart_rx.v(30[17:26])
    defparam n43208_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_SM_Main_2__N_3508[2]), .I1(n34731), .I2(r_SM_Main_c[0]), 
            .I3(r_Bit_Index[0]), .O(n15734));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_993 (.I0(r_SM_Main_2__N_3508[2]), .I1(n34731), 
            .I2(r_SM_Main_c[0]), .I3(r_Bit_Index[0]), .O(n15626));
    defparam i1_2_lut_4_lut_adj_993.LUT_INIT = 16'hfffd;
    SB_LUT4 i18939_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23653));
    defparam i18939_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_135_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_135_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_137_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_137_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_3508[2]), .O(n17052));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0301;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(r_Clock_Count[5]), .I3(n24382), .O(r_SM_Main_2__N_3508[2]));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i33683_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(r_SM_Main_2__N_3508[2]), .O(n40176));   // verilog/uart_rx.v(36[17:26])
    defparam i33683_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12536_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[7]), 
            .I3(r_Clock_Count[7]), .O(n17265));
    defparam i12536_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i1_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[5]), .I3(r_Clock_Count[5]), 
            .O(n45));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12545_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[4]), 
            .I3(r_Clock_Count[4]), .O(n17274));
    defparam i12545_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12539_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[6]), 
            .I3(r_Clock_Count[6]), .O(n17268));
    defparam i12539_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12554_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[1]), 
            .I3(r_Clock_Count[1]), .O(n17283));
    defparam i12554_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12551_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[2]), 
            .I3(r_Clock_Count[2]), .O(n17280));
    defparam i12551_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12548_4_lut_4_lut (.I0(n2588), .I1(n34657), .I2(n194[3]), 
            .I3(r_Clock_Count[3]), .O(n17277));
    defparam i12548_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(n24382), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[6]), .O(n19399));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffb;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n18003, encoder1_position, clk32MHz, 
            n18004, n18005, n18006, n18007, n18008, n18009, n18010, 
            n18011, n18012, n18001, n18002, n17999, n18000, n17997, 
            n17998, n17995, n17996, n17993, n17994, n17990, n17991, 
            n17992, data_o, GND_net, n2944, count_enable, n17401, 
            n18036, PIN_6_c_1, reg_B, n35775, n17413, PIN_7_c_0) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18003;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n18004;
    input n18005;
    input n18006;
    input n18007;
    input n18008;
    input n18009;
    input n18010;
    input n18011;
    input n18012;
    input n18001;
    input n18002;
    input n17999;
    input n18000;
    input n17997;
    input n17998;
    input n17995;
    input n17996;
    input n17993;
    input n17994;
    input n17990;
    input n17991;
    input n17992;
    output [1:0]data_o;
    input GND_net;
    output [23:0]n2944;
    output count_enable;
    input n17401;
    input n18036;
    input PIN_6_c_1;
    output [1:0]reg_B;
    output n35775;
    input n17413;
    input PIN_7_c_0;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, count_direction, n2931, n27961, n27960, 
        n27959, n27958, n27957, n27956, n27955, n27954, n27953, 
        n27952, n27951, n27950, n27949, n27948, n27947, n27946, 
        n27945, n27944, n27943, n27942, n27941, n27940, n27939, 
        n27938;
    
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18003));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18004));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18005));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18006));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18007));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18008));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18009));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18010));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18011));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18012));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18001));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18002));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n17999));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18000));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n17997));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n17998));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n17995));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n17996));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n17993));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n17994));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n17990));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n17991));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n17992));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_608_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2931), 
            .I3(n27961), .O(n2944[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_608_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2931), 
            .I3(n27960), .O(n2944[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_24 (.CI(n27960), .I0(encoder1_position[22]), .I1(n2931), 
            .CO(n27961));
    SB_LUT4 add_608_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2931), 
            .I3(n27959), .O(n2944[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_23 (.CI(n27959), .I0(encoder1_position[21]), .I1(n2931), 
            .CO(n27960));
    SB_LUT4 add_608_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2931), 
            .I3(n27958), .O(n2944[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_22 (.CI(n27958), .I0(encoder1_position[20]), .I1(n2931), 
            .CO(n27959));
    SB_LUT4 add_608_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2931), 
            .I3(n27957), .O(n2944[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_21 (.CI(n27957), .I0(encoder1_position[19]), .I1(n2931), 
            .CO(n27958));
    SB_LUT4 add_608_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2931), 
            .I3(n27956), .O(n2944[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_20 (.CI(n27956), .I0(encoder1_position[18]), .I1(n2931), 
            .CO(n27957));
    SB_LUT4 add_608_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2931), 
            .I3(n27955), .O(n2944[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_19 (.CI(n27955), .I0(encoder1_position[17]), .I1(n2931), 
            .CO(n27956));
    SB_LUT4 add_608_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2931), 
            .I3(n27954), .O(n2944[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_18 (.CI(n27954), .I0(encoder1_position[16]), .I1(n2931), 
            .CO(n27955));
    SB_LUT4 add_608_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2931), 
            .I3(n27953), .O(n2944[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_17 (.CI(n27953), .I0(encoder1_position[15]), .I1(n2931), 
            .CO(n27954));
    SB_LUT4 add_608_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2931), 
            .I3(n27952), .O(n2944[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_16 (.CI(n27952), .I0(encoder1_position[14]), .I1(n2931), 
            .CO(n27953));
    SB_LUT4 add_608_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2931), 
            .I3(n27951), .O(n2944[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_15 (.CI(n27951), .I0(encoder1_position[13]), .I1(n2931), 
            .CO(n27952));
    SB_LUT4 add_608_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2931), 
            .I3(n27950), .O(n2944[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_14 (.CI(n27950), .I0(encoder1_position[12]), .I1(n2931), 
            .CO(n27951));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17401));   // quad.v(35[10] 41[6])
    SB_LUT4 add_608_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2931), 
            .I3(n27949), .O(n2944[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_13 (.CI(n27949), .I0(encoder1_position[11]), .I1(n2931), 
            .CO(n27950));
    SB_LUT4 add_608_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2931), 
            .I3(n27948), .O(n2944[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_12 (.CI(n27948), .I0(encoder1_position[10]), .I1(n2931), 
            .CO(n27949));
    SB_LUT4 add_608_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2931), 
            .I3(n27947), .O(n2944[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_11 (.CI(n27947), .I0(encoder1_position[9]), .I1(n2931), 
            .CO(n27948));
    SB_LUT4 add_608_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2931), 
            .I3(n27946), .O(n2944[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_10 (.CI(n27946), .I0(encoder1_position[8]), .I1(n2931), 
            .CO(n27947));
    SB_LUT4 add_608_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2931), 
            .I3(n27945), .O(n2944[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_9 (.CI(n27945), .I0(encoder1_position[7]), .I1(n2931), 
            .CO(n27946));
    SB_LUT4 add_608_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2931), 
            .I3(n27944), .O(n2944[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_8 (.CI(n27944), .I0(encoder1_position[6]), .I1(n2931), 
            .CO(n27945));
    SB_LUT4 add_608_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2931), 
            .I3(n27943), .O(n2944[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_7 (.CI(n27943), .I0(encoder1_position[5]), .I1(n2931), 
            .CO(n27944));
    SB_LUT4 add_608_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2931), 
            .I3(n27942), .O(n2944[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_6 (.CI(n27942), .I0(encoder1_position[4]), .I1(n2931), 
            .CO(n27943));
    SB_LUT4 add_608_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2931), 
            .I3(n27941), .O(n2944[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_5 (.CI(n27941), .I0(encoder1_position[3]), .I1(n2931), 
            .CO(n27942));
    SB_LUT4 add_608_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2931), 
            .I3(n27940), .O(n2944[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_4 (.CI(n27940), .I0(encoder1_position[2]), .I1(n2931), 
            .CO(n27941));
    SB_LUT4 add_608_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2931), 
            .I3(n27939), .O(n2944[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_3 (.CI(n27939), .I0(encoder1_position[1]), .I1(n2931), 
            .CO(n27940));
    SB_LUT4 add_608_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n27938), .O(n2944[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_608_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_608_2 (.CI(n27938), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n27939));
    SB_CARRY add_608_1 (.CI(GND_net), .I0(n2931), .I1(n2931), .CO(n27938));
    SB_LUT4 i919_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2931));   // quad.v(37[5] 40[8])
    defparam i919_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n18036(n18036), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_6_c_1(PIN_6_c_1), .reg_B({reg_B}), .n35775(n35775), .GND_net(GND_net), 
            .n17413(n17413), .PIN_7_c_0(PIN_7_c_0)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n18036, data_o, clk32MHz, PIN_6_c_1, reg_B, 
            n35775, GND_net, n17413, PIN_7_c_0) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18036;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_6_c_1;
    output [1:0]reg_B;
    output n35775;
    input GND_net;
    input n17413;
    input PIN_7_c_0;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3818, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18036));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_6_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1190__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n35775));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17413));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_7_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n35775), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22771_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22771_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1190__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1190__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22780_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22780_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22773_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22773_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n17983, encoder0_position, clk32MHz, 
            n17984, n17985, n17986, n17987, n17988, n17975, n17976, 
            n17977, n17978, n17979, n17980, n17981, n17982, n17971, 
            n17972, n17973, n17974, n17966, n17967, n17968, n17969, 
            n17970, data_o, count_enable, n17399, n2994, GND_net, 
            n18020, reg_B, n35976, PIN_2_c_0, n17402, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17983;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n17984;
    input n17985;
    input n17986;
    input n17987;
    input n17988;
    input n17975;
    input n17976;
    input n17977;
    input n17978;
    input n17979;
    input n17980;
    input n17981;
    input n17982;
    input n17971;
    input n17972;
    input n17973;
    input n17974;
    input n17966;
    input n17967;
    input n17968;
    input n17969;
    input n17970;
    output [1:0]data_o;
    output count_enable;
    input n17399;
    output [23:0]n2994;
    input GND_net;
    input n18020;
    output [1:0]reg_B;
    output n35976;
    input PIN_2_c_0;
    input n17402;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2990, n27937, n27936, n27935, n27934, 
        n27933, n27932, n27931, n27930, n27929, n27928, n27927, 
        n27926, n27925, n27924, n27923, n27922, n27921, n27920, 
        n27919, n27918, n27917, n27916, n27915, count_direction, 
        n27914;
    
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n17983));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n17984));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n17985));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n17986));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n17987));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n17988));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n17975));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n17976));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n17977));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n17978));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n17979));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n17980));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n17981));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n17982));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n17971));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n17972));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n17973));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n17974));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n17966));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n17967));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n17968));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n17969));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n17970));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17399));   // quad.v(35[10] 41[6])
    SB_LUT4 add_634_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2990), 
            .I3(n27937), .O(n2994[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_634_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2990), 
            .I3(n27936), .O(n2994[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_24 (.CI(n27936), .I0(encoder0_position[22]), .I1(n2990), 
            .CO(n27937));
    SB_LUT4 add_634_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2990), 
            .I3(n27935), .O(n2994[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_23 (.CI(n27935), .I0(encoder0_position[21]), .I1(n2990), 
            .CO(n27936));
    SB_LUT4 add_634_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2990), 
            .I3(n27934), .O(n2994[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_22 (.CI(n27934), .I0(encoder0_position[20]), .I1(n2990), 
            .CO(n27935));
    SB_LUT4 add_634_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2990), 
            .I3(n27933), .O(n2994[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_21 (.CI(n27933), .I0(encoder0_position[19]), .I1(n2990), 
            .CO(n27934));
    SB_LUT4 add_634_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2990), 
            .I3(n27932), .O(n2994[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_20 (.CI(n27932), .I0(encoder0_position[18]), .I1(n2990), 
            .CO(n27933));
    SB_LUT4 add_634_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2990), 
            .I3(n27931), .O(n2994[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_19 (.CI(n27931), .I0(encoder0_position[17]), .I1(n2990), 
            .CO(n27932));
    SB_LUT4 add_634_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2990), 
            .I3(n27930), .O(n2994[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_18 (.CI(n27930), .I0(encoder0_position[16]), .I1(n2990), 
            .CO(n27931));
    SB_LUT4 add_634_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2990), 
            .I3(n27929), .O(n2994[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_17 (.CI(n27929), .I0(encoder0_position[15]), .I1(n2990), 
            .CO(n27930));
    SB_LUT4 add_634_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2990), 
            .I3(n27928), .O(n2994[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_16 (.CI(n27928), .I0(encoder0_position[14]), .I1(n2990), 
            .CO(n27929));
    SB_LUT4 add_634_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2990), 
            .I3(n27927), .O(n2994[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_15 (.CI(n27927), .I0(encoder0_position[13]), .I1(n2990), 
            .CO(n27928));
    SB_LUT4 add_634_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2990), 
            .I3(n27926), .O(n2994[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_14 (.CI(n27926), .I0(encoder0_position[12]), .I1(n2990), 
            .CO(n27927));
    SB_LUT4 add_634_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2990), 
            .I3(n27925), .O(n2994[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_13 (.CI(n27925), .I0(encoder0_position[11]), .I1(n2990), 
            .CO(n27926));
    SB_LUT4 add_634_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2990), 
            .I3(n27924), .O(n2994[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_12 (.CI(n27924), .I0(encoder0_position[10]), .I1(n2990), 
            .CO(n27925));
    SB_LUT4 add_634_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2990), 
            .I3(n27923), .O(n2994[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_11 (.CI(n27923), .I0(encoder0_position[9]), .I1(n2990), 
            .CO(n27924));
    SB_LUT4 add_634_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2990), 
            .I3(n27922), .O(n2994[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_10 (.CI(n27922), .I0(encoder0_position[8]), .I1(n2990), 
            .CO(n27923));
    SB_LUT4 add_634_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2990), 
            .I3(n27921), .O(n2994[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_9 (.CI(n27921), .I0(encoder0_position[7]), .I1(n2990), 
            .CO(n27922));
    SB_LUT4 add_634_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2990), 
            .I3(n27920), .O(n2994[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_8 (.CI(n27920), .I0(encoder0_position[6]), .I1(n2990), 
            .CO(n27921));
    SB_LUT4 add_634_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2990), 
            .I3(n27919), .O(n2994[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_7 (.CI(n27919), .I0(encoder0_position[5]), .I1(n2990), 
            .CO(n27920));
    SB_LUT4 add_634_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2990), 
            .I3(n27918), .O(n2994[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_6 (.CI(n27918), .I0(encoder0_position[4]), .I1(n2990), 
            .CO(n27919));
    SB_LUT4 add_634_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2990), 
            .I3(n27917), .O(n2994[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_5 (.CI(n27917), .I0(encoder0_position[3]), .I1(n2990), 
            .CO(n27918));
    SB_LUT4 add_634_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2990), 
            .I3(n27916), .O(n2994[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_4 (.CI(n27916), .I0(encoder0_position[2]), .I1(n2990), 
            .CO(n27917));
    SB_LUT4 add_634_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2990), 
            .I3(n27915), .O(n2994[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_3 (.CI(n27915), .I0(encoder0_position[1]), .I1(n2990), 
            .CO(n27916));
    SB_LUT4 add_634_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27914), .O(n2994[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_634_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_634_2 (.CI(n27914), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27915));
    SB_CARRY add_634_1 (.CI(GND_net), .I0(n2990), .I1(n2990), .CO(n27914));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i906_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2990));   // quad.v(37[5] 40[8])
    defparam i906_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n18020(n18020), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .n35976(n35976), .GND_net(GND_net), 
            .PIN_2_c_0(PIN_2_c_0), .n17402(n17402), .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18020, data_o, clk32MHz, reg_B, n35976, 
            GND_net, PIN_2_c_0, n17402, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18020;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    output n35976;
    input GND_net;
    input PIN_2_c_0;
    input n17402;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3818, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18020));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1189__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n35976));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17402));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n35976), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22749_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22749_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1189__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1189__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3818));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i22758_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22758_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22751_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22751_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (duty, GND_net, PWMLimit, \Kp[15] , \Kp[3] , \Kp[4] , 
            \Kp[5] , \Kp[1] , \Kp[0] , \Kp[6] , \Kp[7] , \Kp[2] , 
            \Kp[8] , \Kp[10] , clk32MHz, \Kp[9] , \Kp[11] , \Kp[12] , 
            \Kp[13] , \Kp[14] , VCC_net, n25, IntegralLimit, \Ki[3] , 
            \Ki[2] , \Ki[0] , \Ki[1] , n43164, setpoint, \Ki[4] , 
            \Ki[5] , \Ki[6] , motor_state, \Ki[7] , \Ki[8] , \Ki[9] , 
            \Ki[10] , \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] ) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]duty;
    input GND_net;
    input [23:0]PWMLimit;
    input \Kp[15] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[2] ;
    input \Kp[8] ;
    input \Kp[10] ;
    input clk32MHz;
    input \Kp[9] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input VCC_net;
    input n25;
    input [23:0]IntegralLimit;
    input \Ki[3] ;
    input \Ki[2] ;
    input \Ki[0] ;
    input \Ki[1] ;
    output n43164;
    input [23:0]setpoint;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input [23:0]motor_state;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n12, n35, n30, n13, n11, n9, n40780, n41381, n19, 
        n17, n15, n41371, n29457;
    wire [13:0]n7966;
    
    wire n463, n29458;
    wire [14:0]n7949;
    
    wire n390, n29456;
    wire [23:0]duty_23__N_3737;
    wire [23:0]n3050;
    wire [23:0]n3075;
    
    wire n27913, n25_c, n23, n21, n42203, n31, n29, n27, n41735, 
        n37, n33, n42289, n317, n29455, n27912, n27911, n244, 
        n29454, n171, n29453, n6, n41903, n29_adj_3825, n98, n41904;
    wire [15:0]n7931;
    
    wire n29452, n1117, n29451, n27910, n16, n45, n24, n43, 
        n40741, n40650, n8, n40610, n41635, n41166, n4, n41901, 
        n41902, n40726, n40696, n10, n40674, n42193, n41168, n42360, 
        n42361, n39, n42326, n41, n40656, n42112, n41174, n42259, 
        duty_23__N_3761;
    wire [23:0]duty_23__N_3614;
    wire [23:0]n1;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n1114, n241;
    wire [47:0]n155;
    
    wire n256, n314, n27909, n387, n1044, n29450, n95, n26, 
        n460, n533, n971, n29449, n27908, n898, n29448, n825, 
        n29447, n752, n29446, n679, n29445, n606, n29444, n168, 
        n29443, n27907, n29442, n737, n47, n28007;
    wire [23:0]n257;
    
    wire n28006, n29441, n29440, n28005, n28004, n27906, n28003, 
        n28002, n29439, n28001;
    wire [23:0]\PID_CONTROLLER.err_23__N_3638 ;
    
    wire n29438, n28000;
    wire [16:0]n7912;
    
    wire n29437, n29436, n27905;
    wire [23:0]n28;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    
    wire n28598, n29435, n28597, n28596, n28595, n28594, n28593, 
        n1041, n29434, n27999, n28592, n968, n29433, n27904, n27998, 
        n895, n29432, n27903, n27997, n810, n28591, n28590, n883, 
        n28589, n28588, n28587, n28586, n28585, n822, n29431, 
        n28584, n28583, n28582, n28581, n28580, n28579, n749, 
        n29430, n676, n29429, n27996, n28578, n28577, n603, n29428, 
        n28576, n530, n29427, n27902, n27901, n457, n29426, n27900, 
        n384, n29425, n311, n29424, n27899, n238, n29423, n27898, 
        n27995, n165, n29422, n27994, n27897, n23_adj_3835, n92, 
        n27896, n27993, n27895, n27992, n27991, n27990, n27989, 
        n27894;
    wire [17:0]n7892;
    
    wire n29421, n29420, n27893, n27988, n29419, n1111, n29418, 
        n1038, n29417, n27987, n965, n29416, n27892, n27986, n892, 
        n29415, n819, n29414, n746, n29413, n27985, n27891, n40150, 
        n673, n29412;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3713 ;
    wire [23:0]n1_adj_4252;
    
    wire n27984, n45_adj_3845, n27983, n43_adj_3847, n27982, n600, 
        n29411, n41_adj_3849, n27981, n527, n29410, n454, n29409, 
        n381, n29408, n308, n29407, n235, n29406, n162, n29405, 
        n20_adj_3851, n89;
    wire [18:0]n7871;
    
    wire n29404, n39_adj_3852, n27980, n29403, n37_adj_3854, n27979, 
        n29402, n29401, n1108, n29400, n1035, n29399, n35_adj_3856, 
        n27978, n962, n29398, n889, n29397, n33_adj_3858, n27977, 
        n816, n29396, n31_adj_3860, n27976, n29_adj_3862, n27975, 
        n27_adj_3864, n27974, n743, n29395, n25_adj_3866, n27973, 
        n670, n29394, n597, n29393, n524, n29392, n451, n29391, 
        n378, n29390, n305, n29389, n232, n29388, n159, n29387, 
        n17_adj_3868, n86;
    wire [19:0]n7849;
    
    wire n29386, n29385, n29384, n29383, n23_adj_3869, n27972, n29382, 
        n1105, n29381, n21_adj_3871, n27971, n1032, n29380, n959, 
        n29379, n886, n29378, n19_adj_3873, n27970, n813, n29377, 
        n740, n29376, n667, n29375, n594, n29374, n521, n29373, 
        n448, n29372, n375, n29371, n17_adj_3875, n27969, n302, 
        n29370, n229, n29369, n156, n29368, n15_adj_3877, n27968, 
        n14_adj_3879, n83;
    wire [20:0]n7826;
    
    wire n29367, n29366, n13_adj_3880, n27967, n11_adj_3882, n27966, 
        n29365, \PID_CONTROLLER.integral_23__N_3710 , n29364, n29363, 
        n29362, n1102, n29361, n1029, n29360, n9_adj_3884, n27965, 
        n7_adj_3886, n27964, n5_adj_3888, n27963, n956, n3_adj_3891, 
        n27962, n41_adj_3893, n39_adj_3894, n45_adj_3895, n43_adj_3896, 
        n37_adj_3897, n35_adj_3898, n29_adj_3899, n31_adj_3900, n23_adj_3901, 
        n25_adj_3902, n9_adj_3903, n17_adj_3904, n19_adj_3905, n21_adj_3906, 
        n33_adj_3907, n11_adj_3908, n13_adj_3909, n15_adj_3910, n27_adj_3911, 
        n40577, n40518, n12_adj_3912, n10_adj_3913, n30_adj_3914, 
        n40606, n41297, n41287, n42159, n41647, n42261, n16_adj_3915, 
        n6_adj_3916, n41897, n41898, n8_adj_3917, n24_adj_3918, n40433, 
        n40425, n41637, n41176, n4_adj_3919, n41645, n41646, n40485, 
        n40479, n42265, n41178, n42388, n42389, n42363, n40435, 
        n42116, n40, n42118, n40206;
    wire [0:0]n6255;
    
    wire n29359, n29358, n29357, n29356, n664, n29355, n591, n29354, 
        n518, n29353, n445, n29352, n372, n29351, n299, n29350, 
        n226, n29349, n153, n29348, n11_adj_3920, n80;
    wire [21:0]n7802;
    
    wire n29347, n29346, n23909, n4_adj_3921;
    wire [3:0]n8378;
    
    wire n6_adj_3922, n17_adj_3923, n536;
    wire [4:0]n8371;
    
    wire n9_adj_3924, n609, n11_adj_3925, n27618, n682, n755, n828, 
        n901, n40579, n974, n1047, n40465, n1120, n44118, n101, 
        n41563, n32, n174, n247, n320, n41557, n393, n44100, 
        n466, n41553, n539, n612, n41551, n685, n758, n44094, 
        n40822, n831, n904, n40836, n16_adj_3926, n40782, n8_adj_3927, 
        n24_adj_3928, n40889, n977, n1050, n41465, n41453, n104_adj_3929, 
        n35_adj_3930, n177, n250, n42231, n41773, n42293, n323, 
        n396, n469, n542, n40999, n44087, n615, n41539, n44082, 
        n12_adj_3931, n40941, n44105, n10_adj_3932, n688, n30_adj_3933, 
        n761, n42041, n834, n907, n980, n27695;
    wire [1:0]n8389;
    
    wire n4_adj_3934, n107_adj_3935, n40956, n38, n180, n44085, 
        n253, n41821, n326, n399, n472, n44111, n545, n42243, 
        n44076, n618, n691, n764, n42348, n44073, n837, n16_adj_3936, 
        n910, n110_adj_3937;
    wire [2:0]n8384;
    
    wire n40891, n62, n131, n204, n41_adj_3938, n183_adj_3939, n4_adj_3940, 
        n256_adj_3941, n329, n24_adj_3942, n402, n475, n6_adj_3943, 
        n41915, n41916, n548, n40898, n621, n8_adj_3944, n44071, 
        n41631, n694, n767, n41146, n840, n4_adj_3945, n113_adj_3946, 
        n41907, n41908, n12_adj_3947, n44, n40808, n186_adj_3948, 
        n10_adj_3949, n259_adj_3950, n30_adj_3951, n332, n40814, n42191, 
        n405, n478, n551, n41158, n624, n42358, n42359, n697, 
        n42328, n6_adj_3952, n770, n116_adj_3953, n47_adj_3954, n41909, 
        n189, n262_adj_3955, n41910, n335, n40788, n408, n481, 
        n554, n41633, n627, n700, n41156, n40790, n119_adj_3956, 
        n50, n192, n265_adj_3957, n42110, n338, n41164, n42257, 
        n411, n4_adj_3958, n484, n41913, n557, n41914, n630, n122_adj_3959, 
        n53, n40943, n42187, n41148, n195, n42356, n42357, n77, 
        n8_adj_3960, n42330, n40904, n150, n42108, n41154, \PID_CONTROLLER.integral_23__N_3712 , 
        n223, n296, n42255, n268_adj_3961, n369, n442, n515, n29345;
    wire [23:0]n1_adj_4253;
    
    wire n29344, n341, n414, n487, n560, n125_adj_3964, n56, n198, 
        n271_adj_3965, n588, n344, n29343, n417, n6_adj_3967;
    wire [3:0]n8081;
    wire [4:0]n8074;
    
    wire n29342, n29341, n4_adj_3970;
    wire [2:0]n8087;
    wire [1:0]n8092;
    
    wire n490, n12_adj_3971, n8_adj_3972, n11_adj_3973, n6_adj_3974, 
        n29340, n27550, n1096, n29339, n1023, n29338, n950, n29337;
    wire [5:0]n8363;
    
    wire n35988, n490_adj_3975, n29790, n417_adj_3976, n29789, n344_adj_3977, 
        n29788, n271_adj_3978, n29787, n198_adj_3979, n29786, n56_adj_3980, 
        n125_adj_3981;
    wire [6:0]n8354;
    
    wire n560_adj_3982, n29785, n487_adj_3983, n29784, n414_adj_3984, 
        n29783, n341_adj_3985, n29782, n268_adj_3986, n29781, n195_adj_3987, 
        n29780, n53_adj_3988, n122_adj_3989;
    wire [7:0]n8344;
    
    wire n630_adj_3990, n29779, n557_adj_3991, n29778, n484_adj_3992, 
        n29777, n877, n29336, n411_adj_3993, n29776, n18_adj_3994, 
        n804, n29335, n338_adj_3995, n29775, n265_adj_3996, n29774, 
        n192_adj_3997, n29773, n731, n29334, n50_adj_3998, n119_adj_3999, 
        n658, n29333, n585, n29332;
    wire [8:0]n8333;
    
    wire n700_adj_4000, n29772, n627_adj_4001, n29771, n554_adj_4002, 
        n29770, n481_adj_4003, n29769, n408_adj_4004, n29768, n335_adj_4005, 
        n29767, n262_adj_4006, n29766, n189_adj_4007, n29765, n47_adj_4008, 
        n116_adj_4009;
    wire [9:0]n8321;
    
    wire n770_adj_4010, n29764, n697_adj_4011, n29763, n624_adj_4012, 
        n29762, n551_adj_4013, n29761, n478_adj_4014, n29760, n405_adj_4015, 
        n29759, n332_adj_4016, n29758, n512, n29331, n259_adj_4017, 
        n29757, n186_adj_4018, n29756, n44_adj_4019, n113_adj_4020;
    wire [10:0]n8308;
    
    wire n840_adj_4021, n29755, n767_adj_4022, n29754, n694_adj_4023, 
        n29753, n621_adj_4024, n29752, n548_adj_4025, n29751, n13_adj_4026, 
        n475_adj_4027, n29750, n402_adj_4028, n29749, n329_adj_4029, 
        n29748, n256_adj_4030, n29747, n183_adj_4031, n29746, n41_adj_4032, 
        n110_adj_4033, n4_adj_4034, n36490;
    wire [11:0]n8294;
    
    wire n910_adj_4035, n29745, n837_adj_4036, n29744, n764_adj_4037, 
        n29743, n691_adj_4038, n29742, n618_adj_4039, n29741, n545_adj_4040, 
        n29740, n472_adj_4041, n29739, n439, n29330, n399_adj_4042, 
        n29738, n326_adj_4043, n29737, n253_adj_4044, n29736, n180_adj_4045, 
        n29735, n38_adj_4046, n107_adj_4047;
    wire [12:0]n8279;
    
    wire n980_adj_4048, n29734, n77_adj_4049, n8_adj_4050, n907_adj_4051, 
        n29733, n834_adj_4052, n29732, n761_adj_4053, n29731, n688_adj_4054, 
        n29730, n615_adj_4055, n29729, n542_adj_4056, n29728, n469_adj_4057, 
        n29727, n396_adj_4058, n29726, n323_adj_4059, n29725, n250_adj_4060, 
        n29724, n177_adj_4061, n29723, n35_adj_4062, n104_adj_4063;
    wire [13:0]n8263;
    
    wire n1050_adj_4064, n29722, n977_adj_4065, n29721, n366, n29329, 
        n293, n29328, n904_adj_4066, n29720, n831_adj_4068, n29719, 
        n758_adj_4069, n29718, n685_adj_4070, n29717, n612_adj_4071, 
        n29716, n539_adj_4072, n29715, n466_adj_4073, n29714, n393_adj_4074, 
        n29713, n320_adj_4075, n29712, n247_adj_4076, n29711, n220, 
        n29327, n174_adj_4077, n29710, n32_adj_4078, n101_adj_4079;
    wire [14:0]n8246;
    
    wire n1120_adj_4080, n29709, n1047_adj_4081, n29708, n974_adj_4082, 
        n29707, n901_adj_4083, n29706, n828_adj_4084, n29705, n755_adj_4085, 
        n29704, n147, n29326, n682_adj_4086, n29703, n609_adj_4087, 
        n29702, n536_adj_4088, n29701, n463_adj_4089, n29700, n390_adj_4090, 
        n29699, n317_adj_4091, n29698, n244_adj_4092, n29697, n171_adj_4093, 
        n29696, n5_adj_4094, n74, n29_adj_4095, n98_adj_4096;
    wire [15:0]n8228;
    
    wire n29695, n1117_adj_4097, n29694, n29325, n1044_adj_4098, n29693, 
        n971_adj_4099, n29692, n898_adj_4100, n29691, n825_adj_4101, 
        n29690, n752_adj_4102, n29689, n679_adj_4103, n29688, n606_adj_4104, 
        n29687, n533_adj_4105, n29686, n460_adj_4106, n29685, n387_adj_4107, 
        n29684, n29324, n314_adj_4108, n29683, n241_adj_4109, n29682, 
        n168_adj_4110, n29681, n26_adj_4111, n95_adj_4112;
    wire [16:0]n8209;
    
    wire n29680, n29679, n1114_adj_4113, n29678, n1041_adj_4114, n29677, 
        n968_adj_4115, n29676, n895_adj_4116, n29675, n822_adj_4117, 
        n29674, n749_adj_4118, n29673, n676_adj_4119, n29672, n603_adj_4120, 
        n29671, n29323, n530_adj_4121, n29670, n457_adj_4122, n29669, 
        n384_adj_4123, n29668, n311_adj_4124, n29667, n238_adj_4125, 
        n29666, n165_adj_4126, n29665, n150_adj_4127, n23_adj_4128, 
        n92_adj_4129, n223_adj_4130, n296_adj_4131;
    wire [17:0]n8189;
    
    wire n29664, n29663, n29662, n1111_adj_4132, n29661, n1038_adj_4133, 
        n29660, n965_adj_4134, n29659, n892_adj_4135, n29658, n369_adj_4136, 
        n819_adj_4137, n29657, n746_adj_4138, n29656, n673_adj_4139, 
        n29655, n600_adj_4140, n29654, n527_adj_4141, n29653, n454_adj_4142, 
        n29652, n442_adj_4143, n381_adj_4144, n29651, n308_adj_4145, 
        n29650, n235_adj_4146, n29649, n162_adj_4147, n29648, n20_adj_4148, 
        n89_adj_4149;
    wire [18:0]n8168;
    
    wire n29647, n27491, n29646, n29645, n29644, n27525, n1108_adj_4150, 
        n29643, n1035_adj_4151, n29642, n962_adj_4152, n29641, n889_adj_4153, 
        n29640, n816_adj_4154, n29639, n743_adj_4155, n29638, n29322, 
        n670_adj_4156, n29637, n597_adj_4157, n29636, n524_adj_4158, 
        n29635, n451_adj_4159, n29634, n378_adj_4160, n29633, n305_adj_4161, 
        n29632, n232_adj_4162, n29631, n159_adj_4163, n29630, n17_adj_4164, 
        n86_adj_4165;
    wire [19:0]n8146;
    
    wire n29629, n29628, n29627, n29626, n29625, n1105_adj_4166, 
        n29624, n1032_adj_4167, n29623, n959_adj_4168, n29622, n29321, 
        n886_adj_4169, n29621, n813_adj_4170, n29620, n740_adj_4171, 
        n29619, n667_adj_4172, n29618, n594_adj_4173, n29617, n521_adj_4174, 
        n29616, n29320, n448_adj_4175, n29615, n375_adj_4176, n29614, 
        n302_adj_4177, n29613, n229_adj_4178, n29612, n156_adj_4179, 
        n29611, n14_adj_4180, n83_adj_4181;
    wire [20:0]n8123;
    
    wire n29610, n29609, n29608, n29607, n29606, n29605, n1102_adj_4182, 
        n29604, n1029_adj_4183, n29603, n956_adj_4184, n29602, n883_adj_4185, 
        n29601, n810_adj_4186, n29600, n737_adj_4187, n29599, n664_adj_4188, 
        n29598, n591_adj_4189, n29597, n29319, n518_adj_4190, n29596, 
        n445_adj_4191, n29595, n372_adj_4192, n29594, n299_adj_4193, 
        n29593, n226_adj_4194, n29592, n153_adj_4195, n29591, n11_adj_4196, 
        n80_adj_4197;
    wire [21:0]n8099;
    
    wire n29590, n29589, n29588, n29587, n29586, n1099, n29318, 
        n29585, n29584, n29583, n1096_adj_4198, n29582, n28083, 
        n1023_adj_4201, n29581, n950_adj_4202, n29580, n28082, n877_adj_4204, 
        n29579, n1026, n29317, n804_adj_4207, n29578, n731_adj_4208, 
        n29577, n28081, n28080, n658_adj_4211, n29576, n585_adj_4213, 
        n29575, n28079, n512_adj_4215, n29574, n439_adj_4216, n29573, 
        n4_adj_4217, n366_adj_4219, n29572, n28078, n293_adj_4221, 
        n29571, n28077, n28076, n28075, n28074, n953, n29316, 
        n28073, n220_adj_4227, n29570, n147_adj_4228, n29569, n28072, 
        n880, n29315, n28071, n5_adj_4231, n74_adj_4232, n29568, 
        n28070, n29567, n29566, n29565, n807, n29314, n734, n29313, 
        n29564, n29563, n29562, n1099_adj_4234, n29561, n1026_adj_4235, 
        n29560, n953_adj_4236, n29559, n880_adj_4237, n29558, n807_adj_4238, 
        n29557, n734_adj_4239, n29556, n661, n29555, n588_adj_4240, 
        n29554, n661_adj_4241, n29312, n28069, n27448, n28068, n515_adj_4244, 
        n29553, n28067, n28066, n29552, n29551, n29550, n29549, 
        n29548, n28065;
    wire [5:0]n8066;
    
    wire n29547, n28064, n28063, n29546, n29545, n29311, n28062, 
        n29544, n29543, n28061;
    wire [6:0]n8057;
    
    wire n29542, n29541, n29540, n29539, n29310, n29309, n29308, 
        n29538, n29307, n29306, n29305, n29537;
    wire [7:0]n8047;
    
    wire n29536, n29535, n29534, n29533, n29532, n29531, n29530;
    wire [8:0]n8036;
    
    wire n29529, n29528, n29527, n29526, n29525, n29524, n29523, 
        n29522;
    wire [9:0]n8024;
    
    wire n29521, n29520, n29519, n29518, n29517, n29516, n29515, 
        n29514, n29513;
    wire [10:0]n8011;
    
    wire n29512, n29511, n29510, n29509, n29508, n29507, n29506, 
        n29505, n29504, n29503;
    wire [11:0]n7997;
    
    wire n29502, n29501, n29500, n29499, n29498, n29497, n29496, 
        n29495, n29494, n29493, n29492;
    wire [12:0]n7982;
    
    wire n29491, n29490, n29489, n29488, n29487, n29486, n29485, 
        n29484, n29483, n29482, n29481, n29480, n29479, n29478, 
        n29477, n29476, n29475, n29474, n29473, n29472, n29471, 
        n29470, n29469, n29468, n29467, n29466, n29465, n29464, 
        n29463, n29462, n29461, n29460, n29459, n12_adj_4246, n8_adj_4247, 
        n11_adj_4248, n6_adj_4249, n27720, n18_adj_4250, n13_adj_4251;
    
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(duty[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34549_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n40780), 
            .O(n41381));
    defparam i34549_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34539_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n41381), 
            .O(n41371));
    defparam i34539_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3735_7 (.CI(n29457), .I0(n7966[4]), .I1(n463), .CO(n29458));
    SB_LUT4 add_3735_6_lut (.I0(GND_net), .I1(n7966[3]), .I2(n390), .I3(n29456), 
            .O(n7949[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_25_lut (.I0(GND_net), .I1(n3050[23]), .I2(n3075[23]), 
            .I3(n27913), .O(duty_23__N_3737[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35371_4_lut (.I0(n25_c), .I1(n23), .I2(n21), .I3(n41371), 
            .O(n42203));
    defparam i35371_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3735_6 (.CI(n29456), .I0(n7966[3]), .I1(n390), .CO(n29457));
    SB_LUT4 i34903_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n42203), 
            .O(n41735));
    defparam i34903_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35457_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n41735), 
            .O(n42289));
    defparam i35457_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3735_5_lut (.I0(GND_net), .I1(n7966[2]), .I2(n317), .I3(n29455), 
            .O(n7949[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_24_lut (.I0(GND_net), .I1(n3050[22]), .I2(n3075[22]), 
            .I3(n27912), .O(duty_23__N_3737[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_24 (.CI(n27912), .I0(n3050[22]), .I1(n3075[22]), 
            .CO(n27913));
    SB_CARRY add_3735_5 (.CI(n29455), .I0(n7966[2]), .I1(n317), .CO(n29456));
    SB_LUT4 add_642_23_lut (.I0(GND_net), .I1(n3050[21]), .I2(n3075[21]), 
            .I3(n27911), .O(duty_23__N_3737[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_23 (.CI(n27911), .I0(n3050[21]), .I1(n3075[21]), 
            .CO(n27912));
    SB_LUT4 add_3735_4_lut (.I0(GND_net), .I1(n7966[1]), .I2(n244), .I3(n29454), 
            .O(n7949[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_4 (.CI(n29454), .I0(n7966[1]), .I1(n244), .CO(n29455));
    SB_LUT4 add_3735_3_lut (.I0(GND_net), .I1(n7966[0]), .I2(n171), .I3(n29453), 
            .O(n7949[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_3 (.CI(n29453), .I0(n7966[0]), .I1(n171), .CO(n29454));
    SB_LUT4 i35071_3_lut (.I0(n6), .I1(duty[10]), .I2(n21), .I3(GND_net), 
            .O(n41903));   // verilog/motorControl.v(44[10:25])
    defparam i35071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3735_2_lut (.I0(GND_net), .I1(n29_adj_3825), .I2(n98), 
            .I3(GND_net), .O(n7949[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_2 (.CI(GND_net), .I0(n29_adj_3825), .I1(n98), .CO(n29453));
    SB_LUT4 i35072_3_lut (.I0(n41903), .I1(duty[11]), .I2(n23), .I3(GND_net), 
            .O(n41904));   // verilog/motorControl.v(44[10:25])
    defparam i35072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3734_17_lut (.I0(GND_net), .I1(n7949[14]), .I2(GND_net), 
            .I3(n29452), .O(n7931[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3734_16_lut (.I0(GND_net), .I1(n7949[13]), .I2(n1117), 
            .I3(n29451), .O(n7931[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_22_lut (.I0(GND_net), .I1(n3050[20]), .I2(n3075[20]), 
            .I3(n27910), .O(duty_23__N_3737[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(duty[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33818_4_lut (.I0(n43), .I1(n25_c), .I2(n23), .I3(n40741), 
            .O(n40650));
    defparam i33818_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34803_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n40610), 
            .O(n41635));   // verilog/motorControl.v(44[10:25])
    defparam i34803_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34334_3_lut (.I0(n41904), .I1(duty[12]), .I2(n25_c), .I3(GND_net), 
            .O(n41166));   // verilog/motorControl.v(44[10:25])
    defparam i34334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35069_3_lut (.I0(n4), .I1(duty[13]), .I2(n27), .I3(GND_net), 
            .O(n41901));   // verilog/motorControl.v(44[10:25])
    defparam i35069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35070_3_lut (.I0(n41901), .I1(duty[14]), .I2(n29), .I3(GND_net), 
            .O(n41902));   // verilog/motorControl.v(44[10:25])
    defparam i35070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33864_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n40726), 
            .O(n40696));
    defparam i33864_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35361_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n40674), 
            .O(n42193));   // verilog/motorControl.v(44[10:25])
    defparam i35361_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34336_3_lut (.I0(n41902), .I1(duty[15]), .I2(n31), .I3(GND_net), 
            .O(n41168));   // verilog/motorControl.v(44[10:25])
    defparam i34336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35528_4_lut (.I0(n41168), .I1(n42193), .I2(n35), .I3(n40696), 
            .O(n42360));   // verilog/motorControl.v(44[10:25])
    defparam i35528_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35529_3_lut (.I0(n42360), .I1(duty[18]), .I2(n37), .I3(GND_net), 
            .O(n42361));   // verilog/motorControl.v(44[10:25])
    defparam i35529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35494_3_lut (.I0(n42361), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n42326));   // verilog/motorControl.v(44[10:25])
    defparam i35494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33824_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n42289), 
            .O(n40656));
    defparam i33824_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35280_4_lut (.I0(n41166), .I1(n41635), .I2(n45), .I3(n40650), 
            .O(n42112));   // verilog/motorControl.v(44[10:25])
    defparam i35280_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34342_3_lut (.I0(n42326), .I1(duty[20]), .I2(n41), .I3(GND_net), 
            .O(n41174));   // verilog/motorControl.v(44[10:25])
    defparam i34342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35427_4_lut (.I0(n41174), .I1(n42112), .I2(n45), .I3(n40656), 
            .O(n42259));   // verilog/motorControl.v(44[10:25])
    defparam i35427_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35428_3_lut (.I0(n42259), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3761));   // verilog/motorControl.v(44[10:25])
    defparam i35428_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3737[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256), 
            .I3(GND_net), .O(n3075[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_640_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256), 
            .I3(GND_net), .O(n3075[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3734_16 (.CI(n29451), .I0(n7949[13]), .I1(n1117), .CO(n29452));
    SB_CARRY add_642_22 (.CI(n27910), .I0(n3050[20]), .I1(n3075[20]), 
            .CO(n27911));
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_642_21_lut (.I0(GND_net), .I1(n3050[19]), .I2(n3075[19]), 
            .I3(n27909), .O(duty_23__N_3737[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3734_15_lut (.I0(GND_net), .I1(n7949[12]), .I2(n1044), 
            .I3(n29450), .O(n7931[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256), 
            .I3(GND_net), .O(n3075[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3734_15 (.CI(n29450), .I0(n7949[12]), .I1(n1044), .CO(n29451));
    SB_LUT4 add_3734_14_lut (.I0(GND_net), .I1(n7949[11]), .I2(n971), 
            .I3(n29449), .O(n7931[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_21 (.CI(n27909), .I0(n3050[19]), .I1(n3075[19]), 
            .CO(n27910));
    SB_LUT4 add_642_20_lut (.I0(GND_net), .I1(n3050[18]), .I2(n3075[18]), 
            .I3(n27908), .O(duty_23__N_3737[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_14 (.CI(n29449), .I0(n7949[11]), .I1(n971), .CO(n29450));
    SB_CARRY add_642_20 (.CI(n27908), .I0(n3050[18]), .I1(n3075[18]), 
            .CO(n27909));
    SB_LUT4 add_3734_13_lut (.I0(GND_net), .I1(n7949[10]), .I2(n898), 
            .I3(n29448), .O(n7931[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_13 (.CI(n29448), .I0(n7949[10]), .I1(n898), .CO(n29449));
    SB_LUT4 add_3734_12_lut (.I0(GND_net), .I1(n7949[9]), .I2(n825), .I3(n29447), 
            .O(n7931[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_12 (.CI(n29447), .I0(n7949[9]), .I1(n825), .CO(n29448));
    SB_LUT4 add_3734_11_lut (.I0(GND_net), .I1(n7949[8]), .I2(n752), .I3(n29446), 
            .O(n7931[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_11 (.CI(n29446), .I0(n7949[8]), .I1(n752), .CO(n29447));
    SB_LUT4 add_3734_10_lut (.I0(GND_net), .I1(n7949[7]), .I2(n679), .I3(n29445), 
            .O(n7931[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_10 (.CI(n29445), .I0(n7949[7]), .I1(n679), .CO(n29446));
    SB_LUT4 add_3734_9_lut (.I0(GND_net), .I1(n7949[6]), .I2(n606), .I3(n29444), 
            .O(n7931[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_9 (.CI(n29444), .I0(n7949[6]), .I1(n606), .CO(n29445));
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3734_8_lut (.I0(GND_net), .I1(n7949[5]), .I2(n533), .I3(n29443), 
            .O(n7931[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3734_8 (.CI(n29443), .I0(n7949[5]), .I1(n533), .CO(n29444));
    SB_LUT4 add_642_19_lut (.I0(GND_net), .I1(n3050[17]), .I2(n3075[17]), 
            .I3(n27907), .O(duty_23__N_3737[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3734_7_lut (.I0(GND_net), .I1(n7949[4]), .I2(n460), .I3(n29442), 
            .O(n7931[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3734_7 (.CI(n29442), .I0(n7949[4]), .I1(n460), .CO(n29443));
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1[23]), 
            .I3(n28007), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n28006), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3734_6_lut (.I0(GND_net), .I1(n7949[3]), .I2(n387), .I3(n29441), 
            .O(n7931[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3734_6 (.CI(n29441), .I0(n7949[3]), .I1(n387), .CO(n29442));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28006), .I0(GND_net), .I1(n1[22]), 
            .CO(n28007));
    SB_LUT4 add_3734_5_lut (.I0(GND_net), .I1(n7949[2]), .I2(n314), .I3(n29440), 
            .O(n7931[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n28005), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28005), .I0(GND_net), .I1(n1[21]), 
            .CO(n28006));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n28004), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_19 (.CI(n27907), .I0(n3050[17]), .I1(n3075[17]), 
            .CO(n27908));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28004), .I0(GND_net), .I1(n1[20]), 
            .CO(n28005));
    SB_LUT4 add_642_18_lut (.I0(GND_net), .I1(n3050[16]), .I2(n3075[16]), 
            .I3(n27906), .O(duty_23__N_3737[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n28003), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28003), .I0(GND_net), .I1(n1[19]), 
            .CO(n28004));
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_642_18 (.CI(n27906), .I0(n3050[16]), .I1(n3075[16]), 
            .CO(n27907));
    SB_CARRY add_3734_5 (.CI(n29440), .I0(n7949[2]), .I1(n314), .CO(n29441));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n28002), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28002), .I0(GND_net), .I1(n1[18]), 
            .CO(n28003));
    SB_LUT4 add_3734_4_lut (.I0(GND_net), .I1(n7949[1]), .I2(n241), .I3(n29439), 
            .O(n7931[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n28001), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3614[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28001), .I0(GND_net), .I1(n1[17]), 
            .CO(n28002));
    SB_CARRY add_3734_4 (.CI(n29439), .I0(n7949[1]), .I1(n241), .CO(n29440));
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3734_3_lut (.I0(GND_net), .I1(n7949[0]), .I2(n168), .I3(n29438), 
            .O(n7931[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n28000), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3734_3 (.CI(n29438), .I0(n7949[0]), .I1(n168), .CO(n29439));
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28000), .I0(GND_net), .I1(n1[16]), 
            .CO(n28001));
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3734_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7931[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3734_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33909_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n40741));
    defparam i33909_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3734_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n29438));
    SB_LUT4 i33894_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n40726));
    defparam i33894_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3733_18_lut (.I0(GND_net), .I1(n7931[15]), .I2(GND_net), 
            .I3(n29437), .O(n7912[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3733_17_lut (.I0(GND_net), .I1(n7931[14]), .I2(GND_net), 
            .I3(n29436), .O(n7912[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_17_lut (.I0(GND_net), .I1(n3050[15]), .I2(n3075[15]), 
            .I3(n27905), .O(duty_23__N_3737[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n28598), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_17 (.CI(n29436), .I0(n7931[14]), .I1(GND_net), .CO(n29437));
    SB_LUT4 add_3733_16_lut (.I0(GND_net), .I1(n7931[13]), .I2(n1114), 
            .I3(n29435), .O(n7912[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n28597), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_24  (.CI(n28597), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n28598));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n28596), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_23  (.CI(n28596), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n28597));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n28595), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_22  (.CI(n28595), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n28596));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n28594), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_21  (.CI(n28594), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n28595));
    SB_CARRY add_3733_16 (.CI(n29435), .I0(n7931[13]), .I1(n1114), .CO(n29436));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n28593), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_20  (.CI(n28593), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n28594));
    SB_LUT4 add_3733_15_lut (.I0(GND_net), .I1(n7931[12]), .I2(n1041), 
            .I3(n29434), .O(n7912[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n27999), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_17 (.CI(n27905), .I0(n3050[15]), .I1(n3075[15]), 
            .CO(n27906));
    SB_CARRY add_3733_15 (.CI(n29434), .I0(n7931[12]), .I1(n1041), .CO(n29435));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n28592), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3733_14_lut (.I0(GND_net), .I1(n7931[11]), .I2(n968), 
            .I3(n29433), .O(n7912[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_16_lut (.I0(GND_net), .I1(n3050[14]), .I2(n3075[14]), 
            .I3(n27904), .O(duty_23__N_3737[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n27999), .I0(GND_net), .I1(n1[15]), 
            .CO(n28000));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n27998), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3733_14 (.CI(n29433), .I0(n7931[11]), .I1(n968), .CO(n29434));
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256), 
            .I3(GND_net), .O(n3075[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3733_13_lut (.I0(GND_net), .I1(n7931[10]), .I2(n895), 
            .I3(n29432), .O(n7912[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_16 (.CI(n27904), .I0(n3050[14]), .I1(n3075[14]), 
            .CO(n27905));
    SB_LUT4 add_642_15_lut (.I0(GND_net), .I1(n3050[13]), .I2(n3075[13]), 
            .I3(n27903), .O(duty_23__N_3737[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_640_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256), 
            .I3(GND_net), .O(n3075[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n27998), .I0(GND_net), .I1(n1[14]), 
            .CO(n27999));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n27997), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n27997), .I0(GND_net), .I1(n1[13]), 
            .CO(n27998));
    SB_CARRY add_3733_13 (.CI(n29432), .I0(n7931[10]), .I1(n895), .CO(n29433));
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_19  (.CI(n28592), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n28593));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n28591), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_18  (.CI(n28591), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n28592));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n28590), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_17  (.CI(n28590), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n28591));
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n28589), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_16  (.CI(n28589), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n28590));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n28588), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_15  (.CI(n28588), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n28589));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n28587), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_14  (.CI(n28587), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n28588));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n28586), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_13  (.CI(n28586), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n28587));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n28585), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3733_12_lut (.I0(GND_net), .I1(n7931[9]), .I2(n822), .I3(n29431), 
            .O(n7912[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_12  (.CI(n28585), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n28586));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n28584), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_12 (.CI(n29431), .I0(n7931[9]), .I1(n822), .CO(n29432));
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_11  (.CI(n28584), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n28585));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n28583), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_10  (.CI(n28583), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n28584));
    SB_CARRY add_642_15 (.CI(n27903), .I0(n3050[13]), .I1(n3075[13]), 
            .CO(n27904));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n28582), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_9  (.CI(n28582), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n28583));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n28581), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_8  (.CI(n28581), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n28582));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n28580), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_7  (.CI(n28580), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n28581));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n28579), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3733_11_lut (.I0(GND_net), .I1(n7931[8]), .I2(n749), .I3(n29430), 
            .O(n7912[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_6  (.CI(n28579), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n28580));
    SB_CARRY add_3733_11 (.CI(n29430), .I0(n7931[8]), .I1(n749), .CO(n29431));
    SB_LUT4 add_3733_10_lut (.I0(GND_net), .I1(n7931[7]), .I2(n676), .I3(n29429), 
            .O(n7912[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n27996), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n28578), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_10 (.CI(n29429), .I0(n7931[7]), .I1(n676), .CO(n29430));
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_5  (.CI(n28578), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n28579));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n28577), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_4  (.CI(n28577), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n28578));
    SB_LUT4 add_3733_9_lut (.I0(GND_net), .I1(n7931[6]), .I2(n603), .I3(n29428), 
            .O(n7912[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_9 (.CI(n29428), .I0(n7931[6]), .I1(n603), .CO(n29429));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n28576), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_3  (.CI(n28576), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n28577));
    SB_LUT4 \PID_CONTROLLER.integral_1188_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1188_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1188_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n28576));
    SB_LUT4 add_3733_8_lut (.I0(GND_net), .I1(n7931[5]), .I2(n530), .I3(n29427), 
            .O(n7912[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_8 (.CI(n29427), .I0(n7931[5]), .I1(n530), .CO(n29428));
    SB_LUT4 add_642_14_lut (.I0(GND_net), .I1(n3050[12]), .I2(n3075[12]), 
            .I3(n27902), .O(duty_23__N_3737[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_14 (.CI(n27902), .I0(n3050[12]), .I1(n3075[12]), 
            .CO(n27903));
    SB_LUT4 add_642_13_lut (.I0(GND_net), .I1(n3050[11]), .I2(n3075[11]), 
            .I3(n27901), .O(duty_23__N_3737[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3733_7_lut (.I0(GND_net), .I1(n7931[4]), .I2(n457), .I3(n29426), 
            .O(n7912[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_13 (.CI(n27901), .I0(n3050[11]), .I1(n3075[11]), 
            .CO(n27902));
    SB_LUT4 add_642_12_lut (.I0(GND_net), .I1(n3050[10]), .I2(n3075[10]), 
            .I3(n27900), .O(duty_23__N_3737[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_7 (.CI(n29426), .I0(n7931[4]), .I1(n457), .CO(n29427));
    SB_LUT4 add_3733_6_lut (.I0(GND_net), .I1(n7931[3]), .I2(n384), .I3(n29425), 
            .O(n7912[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_12 (.CI(n27900), .I0(n3050[10]), .I1(n3075[10]), 
            .CO(n27901));
    SB_CARRY add_3733_6 (.CI(n29425), .I0(n7931[3]), .I1(n384), .CO(n29426));
    SB_CARRY unary_minus_16_add_3_14 (.CI(n27996), .I0(GND_net), .I1(n1[12]), 
            .CO(n27997));
    SB_LUT4 add_3733_5_lut (.I0(GND_net), .I1(n7931[2]), .I2(n311), .I3(n29424), 
            .O(n7912[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_11_lut (.I0(GND_net), .I1(n3050[9]), .I2(n3075[9]), 
            .I3(n27899), .O(duty_23__N_3737[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_5 (.CI(n29424), .I0(n7931[2]), .I1(n311), .CO(n29425));
    SB_LUT4 add_3733_4_lut (.I0(GND_net), .I1(n7931[1]), .I2(n238), .I3(n29423), 
            .O(n7912[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_11 (.CI(n27899), .I0(n3050[9]), .I1(n3075[9]), .CO(n27900));
    SB_CARRY add_3733_4 (.CI(n29423), .I0(n7931[1]), .I1(n238), .CO(n29424));
    SB_LUT4 add_642_10_lut (.I0(GND_net), .I1(n3050[8]), .I2(n3075[8]), 
            .I3(n27898), .O(duty_23__N_3737[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n27995), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n27995), .I0(GND_net), .I1(n1[11]), 
            .CO(n27996));
    SB_CARRY add_642_10 (.CI(n27898), .I0(n3050[8]), .I1(n3075[8]), .CO(n27899));
    SB_LUT4 add_3733_3_lut (.I0(GND_net), .I1(n7931[0]), .I2(n165), .I3(n29422), 
            .O(n7912[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3733_3 (.CI(n29422), .I0(n7931[0]), .I1(n165), .CO(n29423));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n27994), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_9_lut (.I0(GND_net), .I1(n3050[7]), .I2(n3075[7]), 
            .I3(n27897), .O(duty_23__N_3737[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n27994), .I0(GND_net), .I1(n1[10]), 
            .CO(n27995));
    SB_LUT4 add_3733_2_lut (.I0(GND_net), .I1(n23_adj_3835), .I2(n92), 
            .I3(GND_net), .O(n7912[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3733_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_9 (.CI(n27897), .I0(n3050[7]), .I1(n3075[7]), .CO(n27898));
    SB_LUT4 add_642_8_lut (.I0(GND_net), .I1(n3050[6]), .I2(n3075[6]), 
            .I3(n27896), .O(duty_23__N_3737[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_8 (.CI(n27896), .I0(n3050[6]), .I1(n3075[6]), .CO(n27897));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n27993), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_7_lut (.I0(GND_net), .I1(n3050[5]), .I2(n3075[5]), 
            .I3(n27895), .O(duty_23__N_3737[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n27993), .I0(GND_net), .I1(n1[9]), 
            .CO(n27994));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n27992), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_7 (.CI(n27895), .I0(n3050[5]), .I1(n3075[5]), .CO(n27896));
    SB_CARRY add_3733_2 (.CI(GND_net), .I0(n23_adj_3835), .I1(n92), .CO(n29422));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n27992), .I0(GND_net), .I1(n1[8]), 
            .CO(n27993));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n27991), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n27991), .I0(GND_net), .I1(n1[7]), 
            .CO(n27992));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n27990), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n27990), .I0(GND_net), .I1(n1[6]), 
            .CO(n27991));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n27989), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_6_lut (.I0(GND_net), .I1(n3050[4]), .I2(n3075[4]), 
            .I3(n27894), .O(duty_23__N_3737[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n27989), .I0(GND_net), .I1(n1[5]), 
            .CO(n27990));
    SB_CARRY add_642_6 (.CI(n27894), .I0(n3050[4]), .I1(n3075[4]), .CO(n27895));
    SB_LUT4 add_3732_19_lut (.I0(GND_net), .I1(n7912[16]), .I2(GND_net), 
            .I3(n29421), .O(n7892[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_18_lut (.I0(GND_net), .I1(n7912[15]), .I2(GND_net), 
            .I3(n29420), .O(n7892[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_18 (.CI(n29420), .I0(n7912[15]), .I1(GND_net), .CO(n29421));
    SB_LUT4 add_642_5_lut (.I0(GND_net), .I1(n3050[3]), .I2(n3075[3]), 
            .I3(n27893), .O(duty_23__N_3737[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n27988), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_17_lut (.I0(GND_net), .I1(n7912[14]), .I2(GND_net), 
            .I3(n29419), .O(n7892[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_5 (.CI(n27893), .I0(n3050[3]), .I1(n3075[3]), .CO(n27894));
    SB_CARRY add_3732_17 (.CI(n29419), .I0(n7912[14]), .I1(GND_net), .CO(n29420));
    SB_LUT4 add_3732_16_lut (.I0(GND_net), .I1(n7912[13]), .I2(n1111), 
            .I3(n29418), .O(n7892[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n27988), .I0(GND_net), .I1(n1[4]), 
            .CO(n27989));
    SB_CARRY add_3732_16 (.CI(n29418), .I0(n7912[13]), .I1(n1111), .CO(n29419));
    SB_LUT4 add_3732_15_lut (.I0(GND_net), .I1(n7912[12]), .I2(n1038), 
            .I3(n29417), .O(n7892[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_15 (.CI(n29417), .I0(n7912[12]), .I1(n1038), .CO(n29418));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n27987), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n27987), .I0(GND_net), .I1(n1[3]), 
            .CO(n27988));
    SB_LUT4 add_3732_14_lut (.I0(GND_net), .I1(n7912[11]), .I2(n965), 
            .I3(n29416), .O(n7892[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_14 (.CI(n29416), .I0(n7912[11]), .I1(n965), .CO(n29417));
    SB_LUT4 add_642_4_lut (.I0(GND_net), .I1(n3050[2]), .I2(n3075[2]), 
            .I3(n27892), .O(duty_23__N_3737[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n27986), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3732_13_lut (.I0(GND_net), .I1(n7912[10]), .I2(n892), 
            .I3(n29415), .O(n7892[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_4 (.CI(n27892), .I0(n3050[2]), .I1(n3075[2]), .CO(n27893));
    SB_CARRY add_3732_13 (.CI(n29415), .I0(n7912[10]), .I1(n892), .CO(n29416));
    SB_LUT4 add_3732_12_lut (.I0(GND_net), .I1(n7912[9]), .I2(n819), .I3(n29414), 
            .O(n7892[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_12 (.CI(n29414), .I0(n7912[9]), .I1(n819), .CO(n29415));
    SB_LUT4 add_3732_11_lut (.I0(GND_net), .I1(n7912[8]), .I2(n746), .I3(n29413), 
            .O(n7892[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n27986), .I0(GND_net), .I1(n1[2]), 
            .CO(n27987));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n27985), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_642_3_lut (.I0(GND_net), .I1(n3050[1]), .I2(n3075[1]), 
            .I3(n27891), .O(duty_23__N_3737[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n27985), .I0(GND_net), .I1(n1[1]), 
            .CO(n27986));
    SB_CARRY add_3732_11 (.CI(n29413), .I0(n7912[8]), .I1(n746), .CO(n29414));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n40150)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3732_10_lut (.I0(GND_net), .I1(n7912[7]), .I2(n673), .I3(n29412), 
            .O(n7892[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_642_3 (.CI(n27891), .I0(n3050[1]), .I1(n3075[1]), .CO(n27892));
    SB_CARRY add_3732_10 (.CI(n29412), .I0(n7912[7]), .I1(n673), .CO(n29413));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n27985));
    SB_LUT4 add_642_2_lut (.I0(GND_net), .I1(n3050[0]), .I2(n3075[0]), 
            .I3(GND_net), .O(duty_23__N_3737[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_642_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4252[23]), 
            .I3(n27984), .O(\PID_CONTROLLER.integral_23__N_3713 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4252[22]), .I3(n27983), .O(n45_adj_3845)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n27983), .I0(GND_net), .I1(n1_adj_4252[22]), 
            .CO(n27984));
    SB_CARRY add_642_2 (.CI(GND_net), .I0(n3050[0]), .I1(n3075[0]), .CO(n27891));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4252[21]), .I3(n27982), .O(n43_adj_3847)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3732_9_lut (.I0(GND_net), .I1(n7912[6]), .I2(n600), .I3(n29411), 
            .O(n7892[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_9 (.CI(n29411), .I0(n7912[6]), .I1(n600), .CO(n29412));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n27982), .I0(GND_net), .I1(n1_adj_4252[21]), 
            .CO(n27983));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4252[20]), .I3(n27981), .O(n41_adj_3849)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3732_8_lut (.I0(GND_net), .I1(n7912[5]), .I2(n527), .I3(n29410), 
            .O(n7892[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_8 (.CI(n29410), .I0(n7912[5]), .I1(n527), .CO(n29411));
    SB_LUT4 add_3732_7_lut (.I0(GND_net), .I1(n7912[4]), .I2(n454), .I3(n29409), 
            .O(n7892[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n27981), .I0(GND_net), .I1(n1_adj_4252[20]), 
            .CO(n27982));
    SB_CARRY add_3732_7 (.CI(n29409), .I0(n7912[4]), .I1(n454), .CO(n29410));
    SB_LUT4 add_3732_6_lut (.I0(GND_net), .I1(n7912[3]), .I2(n381), .I3(n29408), 
            .O(n7892[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_6 (.CI(n29408), .I0(n7912[3]), .I1(n381), .CO(n29409));
    SB_LUT4 add_3732_5_lut (.I0(GND_net), .I1(n7912[2]), .I2(n308), .I3(n29407), 
            .O(n7892[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_5 (.CI(n29407), .I0(n7912[2]), .I1(n308), .CO(n29408));
    SB_LUT4 add_3732_4_lut (.I0(GND_net), .I1(n7912[1]), .I2(n235), .I3(n29406), 
            .O(n7892[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_4 (.CI(n29406), .I0(n7912[1]), .I1(n235), .CO(n29407));
    SB_LUT4 add_3732_3_lut (.I0(GND_net), .I1(n7912[0]), .I2(n162), .I3(n29405), 
            .O(n7892[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_3 (.CI(n29405), .I0(n7912[0]), .I1(n162), .CO(n29406));
    SB_LUT4 add_3732_2_lut (.I0(GND_net), .I1(n20_adj_3851), .I2(n89), 
            .I3(GND_net), .O(n7892[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3732_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3732_2 (.CI(GND_net), .I0(n20_adj_3851), .I1(n89), .CO(n29405));
    SB_LUT4 add_3731_20_lut (.I0(GND_net), .I1(n7892[17]), .I2(GND_net), 
            .I3(n29404), .O(n7871[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4252[19]), .I3(n27980), .O(n39_adj_3852)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n27980), .I0(GND_net), .I1(n1_adj_4252[19]), 
            .CO(n27981));
    SB_LUT4 add_3731_19_lut (.I0(GND_net), .I1(n7892[16]), .I2(GND_net), 
            .I3(n29403), .O(n7871[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4252[18]), .I3(n27979), .O(n37_adj_3854)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3731_19 (.CI(n29403), .I0(n7892[16]), .I1(GND_net), .CO(n29404));
    SB_LUT4 add_3731_18_lut (.I0(GND_net), .I1(n7892[15]), .I2(GND_net), 
            .I3(n29402), .O(n7871[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_18 (.CI(n29402), .I0(n7892[15]), .I1(GND_net), .CO(n29403));
    SB_LUT4 add_3731_17_lut (.I0(GND_net), .I1(n7892[14]), .I2(GND_net), 
            .I3(n29401), .O(n7871[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_17 (.CI(n29401), .I0(n7892[14]), .I1(GND_net), .CO(n29402));
    SB_LUT4 add_3731_16_lut (.I0(GND_net), .I1(n7892[13]), .I2(n1108), 
            .I3(n29400), .O(n7871[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_16 (.CI(n29400), .I0(n7892[13]), .I1(n1108), .CO(n29401));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n27979), .I0(GND_net), .I1(n1_adj_4252[18]), 
            .CO(n27980));
    SB_LUT4 add_3731_15_lut (.I0(GND_net), .I1(n7892[12]), .I2(n1035), 
            .I3(n29399), .O(n7871[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_15 (.CI(n29399), .I0(n7892[12]), .I1(n1035), .CO(n29400));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4252[17]), .I3(n27978), .O(n35_adj_3856)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3731_14_lut (.I0(GND_net), .I1(n7892[11]), .I2(n962), 
            .I3(n29398), .O(n7871[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_14 (.CI(n29398), .I0(n7892[11]), .I1(n962), .CO(n29399));
    SB_LUT4 add_3731_13_lut (.I0(GND_net), .I1(n7892[10]), .I2(n889), 
            .I3(n29397), .O(n7871[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_13 (.CI(n29397), .I0(n7892[10]), .I1(n889), .CO(n29398));
    SB_CARRY unary_minus_5_add_3_19 (.CI(n27978), .I0(GND_net), .I1(n1_adj_4252[17]), 
            .CO(n27979));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4252[16]), .I3(n27977), .O(n33_adj_3858)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3731_12_lut (.I0(GND_net), .I1(n7892[9]), .I2(n816), .I3(n29396), 
            .O(n7871[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n27977), .I0(GND_net), .I1(n1_adj_4252[16]), 
            .CO(n27978));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4252[15]), .I3(n27976), .O(n31_adj_3860)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n27976), .I0(GND_net), .I1(n1_adj_4252[15]), 
            .CO(n27977));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4252[14]), .I3(n27975), .O(n29_adj_3862)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n27975), .I0(GND_net), .I1(n1_adj_4252[14]), 
            .CO(n27976));
    SB_CARRY add_3731_12 (.CI(n29396), .I0(n7892[9]), .I1(n816), .CO(n29397));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4252[13]), .I3(n27974), .O(n27_adj_3864)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3731_11_lut (.I0(GND_net), .I1(n7892[8]), .I2(n743), .I3(n29395), 
            .O(n7871[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n27974), .I0(GND_net), .I1(n1_adj_4252[13]), 
            .CO(n27975));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4252[12]), .I3(n27973), .O(n25_adj_3866)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3731_11 (.CI(n29395), .I0(n7892[8]), .I1(n743), .CO(n29396));
    SB_LUT4 add_3731_10_lut (.I0(GND_net), .I1(n7892[7]), .I2(n670), .I3(n29394), 
            .O(n7871[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n27973), .I0(GND_net), .I1(n1_adj_4252[12]), 
            .CO(n27974));
    SB_CARRY add_3731_10 (.CI(n29394), .I0(n7892[7]), .I1(n670), .CO(n29395));
    SB_LUT4 add_3731_9_lut (.I0(GND_net), .I1(n7892[6]), .I2(n597), .I3(n29393), 
            .O(n7871[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_9 (.CI(n29393), .I0(n7892[6]), .I1(n597), .CO(n29394));
    SB_LUT4 add_3731_8_lut (.I0(GND_net), .I1(n7892[5]), .I2(n524), .I3(n29392), 
            .O(n7871[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_8 (.CI(n29392), .I0(n7892[5]), .I1(n524), .CO(n29393));
    SB_LUT4 add_3731_7_lut (.I0(GND_net), .I1(n7892[4]), .I2(n451), .I3(n29391), 
            .O(n7871[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_7 (.CI(n29391), .I0(n7892[4]), .I1(n451), .CO(n29392));
    SB_LUT4 add_3731_6_lut (.I0(GND_net), .I1(n7892[3]), .I2(n378), .I3(n29390), 
            .O(n7871[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_6 (.CI(n29390), .I0(n7892[3]), .I1(n378), .CO(n29391));
    SB_LUT4 add_3731_5_lut (.I0(GND_net), .I1(n7892[2]), .I2(n305), .I3(n29389), 
            .O(n7871[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_5 (.CI(n29389), .I0(n7892[2]), .I1(n305), .CO(n29390));
    SB_LUT4 add_3731_4_lut (.I0(GND_net), .I1(n7892[1]), .I2(n232), .I3(n29388), 
            .O(n7871[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_4 (.CI(n29388), .I0(n7892[1]), .I1(n232), .CO(n29389));
    SB_LUT4 add_3731_3_lut (.I0(GND_net), .I1(n7892[0]), .I2(n159), .I3(n29387), 
            .O(n7871[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_3 (.CI(n29387), .I0(n7892[0]), .I1(n159), .CO(n29388));
    SB_LUT4 add_3731_2_lut (.I0(GND_net), .I1(n17_adj_3868), .I2(n86), 
            .I3(GND_net), .O(n7871[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3731_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3731_2 (.CI(GND_net), .I0(n17_adj_3868), .I1(n86), .CO(n29387));
    SB_LUT4 add_3730_21_lut (.I0(GND_net), .I1(n7871[18]), .I2(GND_net), 
            .I3(n29386), .O(n7849[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3730_20_lut (.I0(GND_net), .I1(n7871[17]), .I2(GND_net), 
            .I3(n29385), .O(n7849[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_20 (.CI(n29385), .I0(n7871[17]), .I1(GND_net), .CO(n29386));
    SB_LUT4 add_3730_19_lut (.I0(GND_net), .I1(n7871[16]), .I2(GND_net), 
            .I3(n29384), .O(n7849[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_19 (.CI(n29384), .I0(n7871[16]), .I1(GND_net), .CO(n29385));
    SB_LUT4 add_3730_18_lut (.I0(GND_net), .I1(n7871[15]), .I2(GND_net), 
            .I3(n29383), .O(n7849[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4252[11]), .I3(n27972), .O(n23_adj_3869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3730_18 (.CI(n29383), .I0(n7871[15]), .I1(GND_net), .CO(n29384));
    SB_LUT4 add_3730_17_lut (.I0(GND_net), .I1(n7871[14]), .I2(GND_net), 
            .I3(n29382), .O(n7849[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_17 (.CI(n29382), .I0(n7871[14]), .I1(GND_net), .CO(n29383));
    SB_LUT4 add_3730_16_lut (.I0(GND_net), .I1(n7871[13]), .I2(n1105), 
            .I3(n29381), .O(n7849[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n27972), .I0(GND_net), .I1(n1_adj_4252[11]), 
            .CO(n27973));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4252[10]), .I3(n27971), .O(n21_adj_3871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3730_16 (.CI(n29381), .I0(n7871[13]), .I1(n1105), .CO(n29382));
    SB_LUT4 add_3730_15_lut (.I0(GND_net), .I1(n7871[12]), .I2(n1032), 
            .I3(n29380), .O(n7849[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_640_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256), 
            .I3(GND_net), .O(n3075[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3730_15 (.CI(n29380), .I0(n7871[12]), .I1(n1032), .CO(n29381));
    SB_LUT4 add_3730_14_lut (.I0(GND_net), .I1(n7871[11]), .I2(n959), 
            .I3(n29379), .O(n7849[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_14 (.CI(n29379), .I0(n7871[11]), .I1(n959), .CO(n29380));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n27971), .I0(GND_net), .I1(n1_adj_4252[10]), 
            .CO(n27972));
    SB_LUT4 add_3730_13_lut (.I0(GND_net), .I1(n7871[10]), .I2(n886), 
            .I3(n29378), .O(n7849[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4252[9]), .I3(n27970), .O(n19_adj_3873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3730_13 (.CI(n29378), .I0(n7871[10]), .I1(n886), .CO(n29379));
    SB_LUT4 add_3730_12_lut (.I0(GND_net), .I1(n7871[9]), .I2(n813), .I3(n29377), 
            .O(n7849[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_12 (.CI(n29377), .I0(n7871[9]), .I1(n813), .CO(n29378));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n27970), .I0(GND_net), .I1(n1_adj_4252[9]), 
            .CO(n27971));
    SB_LUT4 add_3730_11_lut (.I0(GND_net), .I1(n7871[8]), .I2(n740), .I3(n29376), 
            .O(n7849[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_11 (.CI(n29376), .I0(n7871[8]), .I1(n740), .CO(n29377));
    SB_LUT4 add_3730_10_lut (.I0(GND_net), .I1(n7871[7]), .I2(n667), .I3(n29375), 
            .O(n7849[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_10 (.CI(n29375), .I0(n7871[7]), .I1(n667), .CO(n29376));
    SB_LUT4 add_3730_9_lut (.I0(GND_net), .I1(n7871[6]), .I2(n594), .I3(n29374), 
            .O(n7849[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_9 (.CI(n29374), .I0(n7871[6]), .I1(n594), .CO(n29375));
    SB_LUT4 add_3730_8_lut (.I0(GND_net), .I1(n7871[5]), .I2(n521), .I3(n29373), 
            .O(n7849[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_8 (.CI(n29373), .I0(n7871[5]), .I1(n521), .CO(n29374));
    SB_LUT4 add_3730_7_lut (.I0(GND_net), .I1(n7871[4]), .I2(n448), .I3(n29372), 
            .O(n7849[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_7 (.CI(n29372), .I0(n7871[4]), .I1(n448), .CO(n29373));
    SB_LUT4 add_3730_6_lut (.I0(GND_net), .I1(n7871[3]), .I2(n375), .I3(n29371), 
            .O(n7849[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4252[8]), .I3(n27969), .O(n17_adj_3875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3730_6 (.CI(n29371), .I0(n7871[3]), .I1(n375), .CO(n29372));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n27969), .I0(GND_net), .I1(n1_adj_4252[8]), 
            .CO(n27970));
    SB_LUT4 add_3730_5_lut (.I0(GND_net), .I1(n7871[2]), .I2(n302), .I3(n29370), 
            .O(n7849[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_5 (.CI(n29370), .I0(n7871[2]), .I1(n302), .CO(n29371));
    SB_LUT4 add_3730_4_lut (.I0(GND_net), .I1(n7871[1]), .I2(n229), .I3(n29369), 
            .O(n7849[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_4 (.CI(n29369), .I0(n7871[1]), .I1(n229), .CO(n29370));
    SB_LUT4 add_3730_3_lut (.I0(GND_net), .I1(n7871[0]), .I2(n156), .I3(n29368), 
            .O(n7849[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_3 (.CI(n29368), .I0(n7871[0]), .I1(n156), .CO(n29369));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4252[7]), .I3(n27968), .O(n15_adj_3877)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3730_2_lut (.I0(GND_net), .I1(n14_adj_3879), .I2(n83), 
            .I3(GND_net), .O(n7849[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3730_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3730_2 (.CI(GND_net), .I0(n14_adj_3879), .I1(n83), .CO(n29368));
    SB_LUT4 add_3729_22_lut (.I0(GND_net), .I1(n7849[19]), .I2(GND_net), 
            .I3(n29367), .O(n7826[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3729_21_lut (.I0(GND_net), .I1(n7849[18]), .I2(GND_net), 
            .I3(n29366), .O(n7826[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_21 (.CI(n29366), .I0(n7849[18]), .I1(GND_net), .CO(n29367));
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n27968), .I0(GND_net), .I1(n1_adj_4252[7]), 
            .CO(n27969));
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3825));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4252[6]), .I3(n27967), .O(n13_adj_3880)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n27967), .I0(GND_net), .I1(n1_adj_4252[6]), 
            .CO(n27968));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4252[5]), .I3(n27966), .O(n11_adj_3882)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3729_20_lut (.I0(GND_net), .I1(n7849[17]), .I2(GND_net), 
            .I3(n29365), .O(n7826[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_20 (.CI(n29365), .I0(n7849[17]), .I1(GND_net), .CO(n29366));
    SB_DFFE \PID_CONTROLLER.integral_1188__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[0]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256), 
            .I3(GND_net), .O(n3075[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_640_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256), 
            .I3(GND_net), .O(n3075[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3729_19_lut (.I0(GND_net), .I1(n7849[16]), .I2(GND_net), 
            .I3(n29364), .O(n7826[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_19 (.CI(n29364), .I0(n7849[16]), .I1(GND_net), .CO(n29365));
    SB_LUT4 add_3729_18_lut (.I0(GND_net), .I1(n7849[15]), .I2(GND_net), 
            .I3(n29363), .O(n7826[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_18 (.CI(n29363), .I0(n7849[15]), .I1(GND_net), .CO(n29364));
    SB_LUT4 add_3729_17_lut (.I0(GND_net), .I1(n7849[14]), .I2(GND_net), 
            .I3(n29362), .O(n7826[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_17 (.CI(n29362), .I0(n7849[14]), .I1(GND_net), .CO(n29363));
    SB_LUT4 add_3729_16_lut (.I0(GND_net), .I1(n7849[13]), .I2(n1102), 
            .I3(n29361), .O(n7826[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_16 (.CI(n29361), .I0(n7849[13]), .I1(n1102), .CO(n29362));
    SB_LUT4 add_3729_15_lut (.I0(GND_net), .I1(n7849[12]), .I2(n1029), 
            .I3(n29360), .O(n7826[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_15 (.CI(n29360), .I0(n7849[12]), .I1(n1029), .CO(n29361));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n27966), .I0(GND_net), .I1(n1_adj_4252[5]), 
            .CO(n27967));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4252[4]), .I3(n27965), .O(n9_adj_3884)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n27965), .I0(GND_net), .I1(n1_adj_4252[4]), 
            .CO(n27966));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4252[3]), .I3(n27964), .O(n7_adj_3886)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n27964), .I0(GND_net), .I1(n1_adj_4252[3]), 
            .CO(n27965));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4252[2]), .I3(n27963), .O(n5_adj_3888)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n27963), .I0(GND_net), .I1(n1_adj_4252[2]), 
            .CO(n27964));
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4252[1]), .I3(n27962), .O(n3_adj_3891)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n27962), .I0(GND_net), .I1(n1_adj_4252[1]), 
            .CO(n27963));
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3893));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3894));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3895));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3896));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3897));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3898));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3899));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3900));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3901));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3902));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3903));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3904));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3905));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3906));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3907));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3908));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3909));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3910));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3911));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33746_4_lut (.I0(n21_adj_3906), .I1(n19_adj_3905), .I2(n17_adj_3904), 
            .I3(n9_adj_3903), .O(n40577));
    defparam i33746_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33688_4_lut (.I0(n27_adj_3911), .I1(n15_adj_3910), .I2(n13_adj_3909), 
            .I3(n11_adj_3908), .O(n40518));
    defparam i33688_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3907), 
            .I3(GND_net), .O(n12_adj_3912));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3909), 
            .I3(GND_net), .O(n10_adj_3913));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_3912), .I1(n257[17]), .I2(n35_adj_3898), 
            .I3(GND_net), .O(n30_adj_3914));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34465_4_lut (.I0(n13_adj_3909), .I1(n11_adj_3908), .I2(n9_adj_3903), 
            .I3(n40606), .O(n41297));
    defparam i34465_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34455_4_lut (.I0(n19_adj_3905), .I1(n17_adj_3904), .I2(n15_adj_3910), 
            .I3(n41297), .O(n41287));
    defparam i34455_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35327_4_lut (.I0(n25_adj_3902), .I1(n23_adj_3901), .I2(n21_adj_3906), 
            .I3(n41287), .O(n42159));
    defparam i35327_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34815_4_lut (.I0(n31_adj_3900), .I1(n29_adj_3899), .I2(n27_adj_3911), 
            .I3(n42159), .O(n41647));
    defparam i34815_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35429_4_lut (.I0(n37_adj_3897), .I1(n35_adj_3898), .I2(n33_adj_3907), 
            .I3(n41647), .O(n42261));
    defparam i35429_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_3896), 
            .I3(GND_net), .O(n16_adj_3915));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35065_3_lut (.I0(n6_adj_3916), .I1(n257[10]), .I2(n21_adj_3906), 
            .I3(GND_net), .O(n41897));   // verilog/motorControl.v(46[19:35])
    defparam i35065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35066_3_lut (.I0(n41897), .I1(n257[11]), .I2(n23_adj_3901), 
            .I3(GND_net), .O(n41898));   // verilog/motorControl.v(46[19:35])
    defparam i35066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3904), 
            .I3(GND_net), .O(n8_adj_3917));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_3915), .I1(n257[22]), .I2(n45_adj_3895), 
            .I3(GND_net), .O(n24_adj_3918));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33603_4_lut (.I0(n43_adj_3896), .I1(n25_adj_3902), .I2(n23_adj_3901), 
            .I3(n40577), .O(n40433));
    defparam i33603_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34805_4_lut (.I0(n24_adj_3918), .I1(n8_adj_3917), .I2(n45_adj_3895), 
            .I3(n40425), .O(n41637));   // verilog/motorControl.v(46[19:35])
    defparam i34805_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34344_3_lut (.I0(n41898), .I1(n257[12]), .I2(n25_adj_3902), 
            .I3(GND_net), .O(n41176));   // verilog/motorControl.v(46[19:35])
    defparam i34344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n40150), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_3919));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34813_3_lut (.I0(n4_adj_3919), .I1(n257[13]), .I2(n27_adj_3911), 
            .I3(GND_net), .O(n41645));   // verilog/motorControl.v(46[19:35])
    defparam i34813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34814_3_lut (.I0(n41645), .I1(n257[14]), .I2(n29_adj_3899), 
            .I3(GND_net), .O(n41646));   // verilog/motorControl.v(46[19:35])
    defparam i34814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33655_4_lut (.I0(n33_adj_3907), .I1(n31_adj_3900), .I2(n29_adj_3899), 
            .I3(n40518), .O(n40485));
    defparam i33655_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35433_4_lut (.I0(n30_adj_3914), .I1(n10_adj_3913), .I2(n35_adj_3898), 
            .I3(n40479), .O(n42265));   // verilog/motorControl.v(46[19:35])
    defparam i35433_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34346_3_lut (.I0(n41646), .I1(n257[15]), .I2(n31_adj_3900), 
            .I3(GND_net), .O(n41178));   // verilog/motorControl.v(46[19:35])
    defparam i34346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35556_4_lut (.I0(n41178), .I1(n42265), .I2(n35_adj_3898), 
            .I3(n40485), .O(n42388));   // verilog/motorControl.v(46[19:35])
    defparam i35556_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35557_3_lut (.I0(n42388), .I1(n257[18]), .I2(n37_adj_3897), 
            .I3(GND_net), .O(n42389));   // verilog/motorControl.v(46[19:35])
    defparam i35557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35531_3_lut (.I0(n42389), .I1(n257[19]), .I2(n39_adj_3894), 
            .I3(GND_net), .O(n42363));   // verilog/motorControl.v(46[19:35])
    defparam i35531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33605_4_lut (.I0(n43_adj_3896), .I1(n41_adj_3893), .I2(n39_adj_3894), 
            .I3(n42261), .O(n40435));
    defparam i33605_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35284_4_lut (.I0(n41176), .I1(n41637), .I2(n45_adj_3895), 
            .I3(n40433), .O(n42116));   // verilog/motorControl.v(46[19:35])
    defparam i35284_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35490_3_lut (.I0(n42363), .I1(n257[20]), .I2(n41_adj_3893), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(46[19:35])
    defparam i35490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35286_4_lut (.I0(n40), .I1(n42116), .I2(n45_adj_3895), .I3(n40435), 
            .O(n42118));   // verilog/motorControl.v(46[19:35])
    defparam i35286_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35287_3_lut (.I0(n42118), .I1(duty[23]), .I2(n47), .I3(GND_net), 
            .O(n256));   // verilog/motorControl.v(46[19:35])
    defparam i35287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_640_i24_3_lut (.I0(n40206), .I1(PWMLimit[23]), .I2(n256), 
            .I3(GND_net), .O(n3075[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i19211_2_lut (.I0(n6255[0]), .I1(n256), .I2(GND_net), .I3(GND_net), 
            .O(n3050[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i19211_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4252[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3713 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4252[0]), 
            .CO(n27962));
    SB_LUT4 add_3729_14_lut (.I0(GND_net), .I1(n7849[11]), .I2(n956), 
            .I3(n29359), .O(n7826[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_14 (.CI(n29359), .I0(n7849[11]), .I1(n956), .CO(n29360));
    SB_LUT4 add_3729_13_lut (.I0(GND_net), .I1(n7849[10]), .I2(n883), 
            .I3(n29358), .O(n7826[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_13 (.CI(n29358), .I0(n7849[10]), .I1(n883), .CO(n29359));
    SB_LUT4 add_3729_12_lut (.I0(GND_net), .I1(n7849[9]), .I2(n810), .I3(n29357), 
            .O(n7826[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_12 (.CI(n29357), .I0(n7849[9]), .I1(n810), .CO(n29358));
    SB_LUT4 add_3729_11_lut (.I0(GND_net), .I1(n7849[8]), .I2(n737), .I3(n29356), 
            .O(n7826[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_11 (.CI(n29356), .I0(n7849[8]), .I1(n737), .CO(n29357));
    SB_LUT4 add_3729_10_lut (.I0(GND_net), .I1(n7849[7]), .I2(n664), .I3(n29355), 
            .O(n7826[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_10 (.CI(n29355), .I0(n7849[7]), .I1(n664), .CO(n29356));
    SB_LUT4 add_3729_9_lut (.I0(GND_net), .I1(n7849[6]), .I2(n591), .I3(n29354), 
            .O(n7826[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_9 (.CI(n29354), .I0(n7849[6]), .I1(n591), .CO(n29355));
    SB_LUT4 add_3729_8_lut (.I0(GND_net), .I1(n7849[5]), .I2(n518), .I3(n29353), 
            .O(n7826[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_8 (.CI(n29353), .I0(n7849[5]), .I1(n518), .CO(n29354));
    SB_LUT4 add_3729_7_lut (.I0(GND_net), .I1(n7849[4]), .I2(n445), .I3(n29352), 
            .O(n7826[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_7 (.CI(n29352), .I0(n7849[4]), .I1(n445), .CO(n29353));
    SB_LUT4 add_3729_6_lut (.I0(GND_net), .I1(n7849[3]), .I2(n372), .I3(n29351), 
            .O(n7826[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_6 (.CI(n29351), .I0(n7849[3]), .I1(n372), .CO(n29352));
    SB_LUT4 add_3729_5_lut (.I0(GND_net), .I1(n7849[2]), .I2(n299), .I3(n29350), 
            .O(n7826[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_5 (.CI(n29350), .I0(n7849[2]), .I1(n299), .CO(n29351));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3614[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_3729_4_lut (.I0(GND_net), .I1(n7849[1]), .I2(n226), .I3(n29349), 
            .O(n7826[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_4 (.CI(n29349), .I0(n7849[1]), .I1(n226), .CO(n29350));
    SB_LUT4 add_3729_3_lut (.I0(GND_net), .I1(n7849[0]), .I2(n153), .I3(n29348), 
            .O(n7826[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3614[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3614[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3614[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3614[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3614[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3614[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3614[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3614[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3614[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3614[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3614[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3614[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3614[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3614[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3614[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3614[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3614[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3614[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3614[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3614[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3614[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3614[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3638 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_3729_3 (.CI(n29348), .I0(n7849[0]), .I1(n153), .CO(n29349));
    SB_LUT4 add_3729_2_lut (.I0(GND_net), .I1(n11_adj_3920), .I2(n80), 
            .I3(GND_net), .O(n7826[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3729_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3729_2 (.CI(GND_net), .I0(n11_adj_3920), .I1(n80), .CO(n29348));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7802[21]), 
            .I2(GND_net), .I3(n29347), .O(n6255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n23909), .I1(n7802[20]), .I2(GND_net), 
            .I3(n29346), .O(n3050[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22967_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_3921), .I3(n8378[1]), .O(n6_adj_3922));   // verilog/motorControl.v(42[26:37])
    defparam i22967_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_3923));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8378[1]), .I3(n4_adj_3921), .O(n8371[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_3924));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_3925));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_973 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8378[0]), .I3(n27618), .O(n8371[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_973.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33748_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n40579));
    defparam i33748_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22959_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n27618), .I3(n8378[0]), .O(n4_adj_3921));   // verilog/motorControl.v(42[26:37])
    defparam i22959_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i33635_3_lut (.I0(n11_adj_3925), .I1(n9_adj_3924), .I2(n40579), 
            .I3(GND_net), .O(n40465));
    defparam i33635_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_458_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n44118));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_458_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34731_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44118), 
            .I2(IntegralLimit[7]), .I3(n40465), .O(n41563));
    defparam i34731_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34725_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3923), 
            .I2(IntegralLimit[9]), .I3(n41563), .O(n41557));
    defparam i34725_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_440_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n44100));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_440_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34721_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3923), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3924), .O(n41553));
    defparam i34721_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i22948_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n27618));   // verilog/motorControl.v(42[26:37])
    defparam i22948_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34719_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44100), 
            .I2(IntegralLimit[11]), .I3(n41553), .O(n41551));
    defparam i34719_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_434_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n44094));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_434_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33990_4_lut (.I0(n27_adj_3864), .I1(n15_adj_3877), .I2(n13_adj_3880), 
            .I3(n11_adj_3882), .O(n40822));
    defparam i33990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i22946_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n8371[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22946_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34004_4_lut (.I0(n21_adj_3871), .I1(n19_adj_3873), .I2(n17_adj_3875), 
            .I3(n9_adj_3884), .O(n40836));
    defparam i34004_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_3847), .I3(GND_net), 
            .O(n16_adj_3926));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i33950_2_lut (.I0(n43_adj_3847), .I1(n19_adj_3873), .I2(GND_net), 
            .I3(GND_net), .O(n40782));
    defparam i33950_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3875), .I3(GND_net), 
            .O(n8_adj_3927));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_3926), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_3845), .I3(GND_net), 
            .O(n24_adj_3928));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34057_2_lut (.I0(n7_adj_3886), .I1(n5_adj_3888), .I2(GND_net), 
            .I3(GND_net), .O(n40889));
    defparam i34057_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34633_4_lut (.I0(n13_adj_3880), .I1(n11_adj_3882), .I2(n9_adj_3884), 
            .I3(n40889), .O(n41465));
    defparam i34633_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34621_4_lut (.I0(n19_adj_3873), .I1(n17_adj_3875), .I2(n15_adj_3877), 
            .I3(n41465), .O(n41453));
    defparam i34621_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3929));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3930));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35399_4_lut (.I0(n25_adj_3866), .I1(n23_adj_3869), .I2(n21_adj_3871), 
            .I3(n41453), .O(n42231));
    defparam i35399_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34941_4_lut (.I0(n31_adj_3860), .I1(n29_adj_3862), .I2(n27_adj_3864), 
            .I3(n42231), .O(n41773));
    defparam i34941_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35461_4_lut (.I0(n37_adj_3854), .I1(n35_adj_3856), .I2(n33_adj_3858), 
            .I3(n41773), .O(n42293));
    defparam i35461_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34167_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44118), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3925), .O(n40999));
    defparam i34167_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_427_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n44087));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_427_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34707_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n44087), 
            .I2(IntegralLimit[14]), .I3(n40999), .O(n41539));
    defparam i34707_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_422_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n44082));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_422_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_3931));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34109_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n40941));
    defparam i34109_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_445_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n44105));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_445_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3932));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_3931), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_3933));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35209_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44100), 
            .I2(IntegralLimit[11]), .I3(n41557), .O(n42041));
    defparam i35209_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23029_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n27695), .I3(n8389[0]), .O(n4_adj_3934));   // verilog/motorControl.v(42[26:37])
    defparam i23029_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3935));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34124_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n44094), 
            .I2(IntegralLimit[13]), .I3(n42041), .O(n40956));
    defparam i34124_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_425_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n44085));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_425_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34989_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n44085), 
            .I2(IntegralLimit[15]), .I3(n40956), .O(n41821));
    defparam i34989_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_451_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n44111));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_451_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35411_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n44111), 
            .I2(IntegralLimit[17]), .I3(n41821), .O(n42243));
    defparam i35411_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_416_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n44076));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_416_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35516_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n44076), 
            .I2(IntegralLimit[19]), .I3(n42243), .O(n42348));
    defparam i35516_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_413_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n44073));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_413_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3936));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3937));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_974 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n8389[0]), .I3(n27695), .O(n8384[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_974.LUT_INIT = 16'h8778;
    SB_LUT4 i34059_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n40891));
    defparam i34059_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(n62), .I1(n131), .I2(n8384[0]), 
            .I3(n204), .O(n8378[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3938));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3939));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22998_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n8384[0]), 
            .O(n4_adj_3940));   // verilog/motorControl.v(42[26:37])
    defparam i22998_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3941));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23016_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8384[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23016_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3936), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3942));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3943));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35083_3_lut (.I0(n6_adj_3943), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n41915));   // verilog/motorControl.v(39[10:34])
    defparam i35083_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35084_3_lut (.I0(n41915), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n41916));   // verilog/motorControl.v(39[10:34])
    defparam i35084_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i23018_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n27695));   // verilog/motorControl.v(42[26:37])
    defparam i23018_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34066_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n44094), 
            .I2(IntegralLimit[21]), .I3(n41551), .O(n40898));
    defparam i34066_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34799_4_lut (.I0(n24_adj_3942), .I1(n8_adj_3944), .I2(n44071), 
            .I3(n40891), .O(n41631));   // verilog/motorControl.v(39[10:34])
    defparam i34799_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34314_3_lut (.I0(n41916), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n41146));   // verilog/motorControl.v(39[10:34])
    defparam i34314_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3713 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_3891), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_3945));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3946));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35075_3_lut (.I0(n4_adj_3945), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_3864), .I3(GND_net), .O(n41907));   // verilog/motorControl.v(39[38:63])
    defparam i35075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35076_3_lut (.I0(n41907), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_3862), .I3(GND_net), .O(n41908));   // verilog/motorControl.v(39[38:63])
    defparam i35076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_3858), .I3(GND_net), 
            .O(n12_adj_3947));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33976_2_lut (.I0(n33_adj_3858), .I1(n15_adj_3877), .I2(GND_net), 
            .I3(GND_net), .O(n40808));
    defparam i33976_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3948));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3880), .I3(GND_net), 
            .O(n10_adj_3949));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3950));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3947), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_3856), .I3(GND_net), 
            .O(n30_adj_3951));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33982_4_lut (.I0(n33_adj_3858), .I1(n31_adj_3860), .I2(n29_adj_3862), 
            .I3(n40822), .O(n40814));
    defparam i33982_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35359_4_lut (.I0(n30_adj_3951), .I1(n10_adj_3949), .I2(n35_adj_3856), 
            .I3(n40808), .O(n42191));   // verilog/motorControl.v(39[38:63])
    defparam i35359_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34326_3_lut (.I0(n41908), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_3860), .I3(GND_net), .O(n41158));   // verilog/motorControl.v(39[38:63])
    defparam i34326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35526_4_lut (.I0(n41158), .I1(n42191), .I2(n35_adj_3856), 
            .I3(n40814), .O(n42358));   // verilog/motorControl.v(39[38:63])
    defparam i35526_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35527_3_lut (.I0(n42358), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_3854), .I3(GND_net), .O(n42359));   // verilog/motorControl.v(39[38:63])
    defparam i35527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35496_3_lut (.I0(n42359), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_3852), .I3(GND_net), .O(n42328));   // verilog/motorControl.v(39[38:63])
    defparam i35496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_3886), .I3(GND_net), 
            .O(n6_adj_3952));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3953));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3954));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35077_3_lut (.I0(n6_adj_3952), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_3871), .I3(GND_net), .O(n41909));   // verilog/motorControl.v(39[38:63])
    defparam i35077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3955));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35078_3_lut (.I0(n41909), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_3869), .I3(GND_net), .O(n41910));   // verilog/motorControl.v(39[38:63])
    defparam i35078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33956_4_lut (.I0(n43_adj_3847), .I1(n25_adj_3866), .I2(n23_adj_3869), 
            .I3(n40836), .O(n40788));
    defparam i33956_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34801_4_lut (.I0(n24_adj_3928), .I1(n8_adj_3927), .I2(n45_adj_3845), 
            .I3(n40782), .O(n41633));   // verilog/motorControl.v(39[38:63])
    defparam i34801_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34324_3_lut (.I0(n41910), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_3866), .I3(GND_net), .O(n41156));   // verilog/motorControl.v(39[38:63])
    defparam i34324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33958_4_lut (.I0(n43_adj_3847), .I1(n41_adj_3849), .I2(n39_adj_3852), 
            .I3(n42293), .O(n40790));
    defparam i33958_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3956));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3957));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35278_4_lut (.I0(n41156), .I1(n41633), .I2(n45_adj_3845), 
            .I3(n40788), .O(n42110));   // verilog/motorControl.v(39[38:63])
    defparam i35278_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34332_3_lut (.I0(n42328), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_3849), .I3(GND_net), .O(n41164));   // verilog/motorControl.v(39[38:63])
    defparam i34332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35425_4_lut (.I0(n41164), .I1(n42110), .I2(n45_adj_3845), 
            .I3(n40790), .O(n42257));   // verilog/motorControl.v(39[38:63])
    defparam i35425_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3958));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35081_3_lut (.I0(n4_adj_3958), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n41913));   // verilog/motorControl.v(39[10:34])
    defparam i35081_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35082_3_lut (.I0(n41913), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n41914));   // verilog/motorControl.v(39[10:34])
    defparam i35082_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3959));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34111_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n44082), 
            .I2(IntegralLimit[16]), .I3(n41539), .O(n40943));
    defparam i34111_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35355_4_lut (.I0(n30_adj_3933), .I1(n10_adj_3932), .I2(n44105), 
            .I3(n40941), .O(n42187));   // verilog/motorControl.v(39[10:34])
    defparam i35355_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34316_3_lut (.I0(n41914), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n41148));   // verilog/motorControl.v(39[10:34])
    defparam i34316_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35524_4_lut (.I0(n41148), .I1(n42187), .I2(n44105), .I3(n40943), 
            .O(n42356));   // verilog/motorControl.v(39[10:34])
    defparam i35524_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35525_3_lut (.I0(n42356), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n42357));   // verilog/motorControl.v(39[10:34])
    defparam i35525_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3960));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35498_3_lut (.I0(n42357), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n42330));   // verilog/motorControl.v(39[10:34])
    defparam i35498_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34072_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n44073), 
            .I2(IntegralLimit[21]), .I3(n42348), .O(n40904));
    defparam i34072_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_411_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n44071));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_411_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35276_4_lut (.I0(n41146), .I1(n41631), .I2(n44071), .I3(n40898), 
            .O(n42108));   // verilog/motorControl.v(39[10:34])
    defparam i35276_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34322_3_lut (.I0(n42330), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n41154));   // verilog/motorControl.v(39[10:34])
    defparam i34322_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35426_3_lut (.I0(n42257), .I1(\PID_CONTROLLER.integral_23__N_3713 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3712 ));   // verilog/motorControl.v(39[38:63])
    defparam i35426_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35423_4_lut (.I0(n41154), .I1(n42108), .I2(n44071), .I3(n40904), 
            .O(n42255));   // verilog/motorControl.v(39[10:34])
    defparam i35423_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3961));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_967_4_lut  (.I0(n42255), .I1(\PID_CONTROLLER.integral_23__N_3712 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3710 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_967_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_23 (.CI(n29346), .I0(n7802[20]), .I1(GND_net), 
            .CO(n29347));
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n23909), .I1(n7802[19]), .I2(GND_net), 
            .I3(n29345), .O(n3050[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36334_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43164));   // verilog/motorControl.v(37[14] 56[8])
    defparam i36334_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_22 (.CI(n29345), .I0(n7802[19]), .I1(GND_net), 
            .CO(n29346));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n23909), .I1(n7802[18]), .I2(GND_net), 
            .I3(n29344), .O(n3050[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_21 (.CI(n29344), .I0(n7802[18]), .I1(GND_net), 
            .CO(n29345));
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3964));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3965));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n23909), .I1(n7802[17]), .I2(GND_net), 
            .I3(n29343), .O(n3050[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_20 (.CI(n29343), .I0(n7802[17]), .I1(GND_net), 
            .CO(n29344));
    SB_LUT4 i2_4_lut (.I0(n6_adj_3967), .I1(\Kp[4] ), .I2(n8081[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8074[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n23909), .I1(n7802[16]), .I2(GND_net), 
            .I3(n29342), .O(n3050[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_19 (.CI(n29342), .I0(n7802[16]), .I1(GND_net), 
            .CO(n29343));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n23909), .I1(n7802[15]), .I2(GND_net), 
            .I3(n29341), .O(n3050[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_18 (.CI(n29341), .I0(n7802[15]), .I1(GND_net), 
            .CO(n29342));
    SB_LUT4 i2_4_lut_adj_976 (.I0(n4_adj_3970), .I1(\Kp[3] ), .I2(n8087[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8081[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_976.LUT_INIT = 16'h965a;
    SB_LUT4 i22879_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8092[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22879_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_977 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_3971));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_977.LUT_INIT = 16'h9c50;
    SB_DFFE \PID_CONTROLLER.integral_1188__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[1]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1188__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3710 ), .D(n28[23]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 i22815_4_lut (.I0(n8081[2]), .I1(\Kp[4] ), .I2(n6_adj_3967), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_3972));   // verilog/motorControl.v(42[17:23])
    defparam i22815_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_3973));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22846_4_lut (.I0(n8087[1]), .I1(\Kp[3] ), .I2(n4_adj_3970), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_3974));   // verilog/motorControl.v(42[17:23])
    defparam i22846_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n23909), .I1(n7802[14]), .I2(GND_net), 
            .I3(n29340), .O(n3050[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_17 (.CI(n29340), .I0(n7802[14]), .I1(GND_net), 
            .CO(n29341));
    SB_LUT4 i22881_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n27550));   // verilog/motorControl.v(42[17:23])
    defparam i22881_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n23909), .I1(n7802[13]), .I2(n1096), 
            .I3(n29339), .O(n3050[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_16 (.CI(n29339), .I0(n7802[13]), .I1(n1096), 
            .CO(n29340));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n23909), .I1(n7802[12]), .I2(n1023), 
            .I3(n29338), .O(n3050[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_15 (.CI(n29338), .I0(n7802[12]), .I1(n1023), 
            .CO(n29339));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n23909), .I1(n7802[11]), .I2(n950), 
            .I3(n29337), .O(n3050[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3766_7_lut (.I0(GND_net), .I1(n35988), .I2(n490_adj_3975), 
            .I3(n29790), .O(n8363[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n29337), .I0(n7802[11]), .I1(n950), 
            .CO(n29338));
    SB_LUT4 add_3766_6_lut (.I0(GND_net), .I1(n8371[3]), .I2(n417_adj_3976), 
            .I3(n29789), .O(n8363[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3766_6 (.CI(n29789), .I0(n8371[3]), .I1(n417_adj_3976), 
            .CO(n29790));
    SB_LUT4 add_3766_5_lut (.I0(GND_net), .I1(n8371[2]), .I2(n344_adj_3977), 
            .I3(n29788), .O(n8363[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3766_5 (.CI(n29788), .I0(n8371[2]), .I1(n344_adj_3977), 
            .CO(n29789));
    SB_LUT4 add_3766_4_lut (.I0(GND_net), .I1(n8371[1]), .I2(n271_adj_3978), 
            .I3(n29787), .O(n8363[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3766_4 (.CI(n29787), .I0(n8371[1]), .I1(n271_adj_3978), 
            .CO(n29788));
    SB_LUT4 add_3766_3_lut (.I0(GND_net), .I1(n8371[0]), .I2(n198_adj_3979), 
            .I3(n29786), .O(n8363[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3766_3 (.CI(n29786), .I0(n8371[0]), .I1(n198_adj_3979), 
            .CO(n29787));
    SB_LUT4 add_3766_2_lut (.I0(GND_net), .I1(n56_adj_3980), .I2(n125_adj_3981), 
            .I3(GND_net), .O(n8363[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3766_2 (.CI(GND_net), .I0(n56_adj_3980), .I1(n125_adj_3981), 
            .CO(n29786));
    SB_LUT4 add_3765_8_lut (.I0(GND_net), .I1(n8363[5]), .I2(n560_adj_3982), 
            .I3(n29785), .O(n8354[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3765_7_lut (.I0(GND_net), .I1(n8363[4]), .I2(n487_adj_3983), 
            .I3(n29784), .O(n8354[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_7 (.CI(n29784), .I0(n8363[4]), .I1(n487_adj_3983), 
            .CO(n29785));
    SB_LUT4 add_3765_6_lut (.I0(GND_net), .I1(n8363[3]), .I2(n414_adj_3984), 
            .I3(n29783), .O(n8354[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_6 (.CI(n29783), .I0(n8363[3]), .I1(n414_adj_3984), 
            .CO(n29784));
    SB_LUT4 add_3765_5_lut (.I0(GND_net), .I1(n8363[2]), .I2(n341_adj_3985), 
            .I3(n29782), .O(n8354[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_5 (.CI(n29782), .I0(n8363[2]), .I1(n341_adj_3985), 
            .CO(n29783));
    SB_LUT4 add_3765_4_lut (.I0(GND_net), .I1(n8363[1]), .I2(n268_adj_3986), 
            .I3(n29781), .O(n8354[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_4 (.CI(n29781), .I0(n8363[1]), .I1(n268_adj_3986), 
            .CO(n29782));
    SB_LUT4 add_3765_3_lut (.I0(GND_net), .I1(n8363[0]), .I2(n195_adj_3987), 
            .I3(n29780), .O(n8354[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_3 (.CI(n29780), .I0(n8363[0]), .I1(n195_adj_3987), 
            .CO(n29781));
    SB_LUT4 add_3765_2_lut (.I0(GND_net), .I1(n53_adj_3988), .I2(n122_adj_3989), 
            .I3(GND_net), .O(n8354[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3765_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3765_2 (.CI(GND_net), .I0(n53_adj_3988), .I1(n122_adj_3989), 
            .CO(n29780));
    SB_LUT4 add_3764_9_lut (.I0(GND_net), .I1(n8354[6]), .I2(n630_adj_3990), 
            .I3(n29779), .O(n8344[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3764_8_lut (.I0(GND_net), .I1(n8354[5]), .I2(n557_adj_3991), 
            .I3(n29778), .O(n8344[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3764_8 (.CI(n29778), .I0(n8354[5]), .I1(n557_adj_3991), 
            .CO(n29779));
    SB_LUT4 add_3764_7_lut (.I0(GND_net), .I1(n8354[4]), .I2(n484_adj_3992), 
            .I3(n29777), .O(n8344[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3764_7 (.CI(n29777), .I0(n8354[4]), .I1(n484_adj_3992), 
            .CO(n29778));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n23909), .I1(n7802[10]), .I2(n877), 
            .I3(n29336), .O(n3050[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n29336), .I0(n7802[10]), .I1(n877), 
            .CO(n29337));
    SB_LUT4 add_3764_6_lut (.I0(GND_net), .I1(n8354[3]), .I2(n411_adj_3993), 
            .I3(n29776), .O(n8344[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3974), .I1(n11_adj_3973), .I2(n8_adj_3972), 
            .I3(n12_adj_3971), .O(n18_adj_3994));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3764_6 (.CI(n29776), .I0(n8354[3]), .I1(n411_adj_3993), 
            .CO(n29777));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n23909), .I1(n7802[9]), .I2(n804), 
            .I3(n29335), .O(n3050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3764_5_lut (.I0(GND_net), .I1(n8354[2]), .I2(n338_adj_3995), 
            .I3(n29775), .O(n8344[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3764_5 (.CI(n29775), .I0(n8354[2]), .I1(n338_adj_3995), 
            .CO(n29776));
    SB_CARRY mult_10_add_1225_12 (.CI(n29335), .I0(n7802[9]), .I1(n804), 
            .CO(n29336));
    SB_LUT4 add_3764_4_lut (.I0(GND_net), .I1(n8354[1]), .I2(n265_adj_3996), 
            .I3(n29774), .O(n8344[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3764_4 (.CI(n29774), .I0(n8354[1]), .I1(n265_adj_3996), 
            .CO(n29775));
    SB_LUT4 add_3764_3_lut (.I0(GND_net), .I1(n8354[0]), .I2(n192_adj_3997), 
            .I3(n29773), .O(n8344[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3764_3 (.CI(n29773), .I0(n8354[0]), .I1(n192_adj_3997), 
            .CO(n29774));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n23909), .I1(n7802[8]), .I2(n731), 
            .I3(n29334), .O(n3050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_11 (.CI(n29334), .I0(n7802[8]), .I1(n731), 
            .CO(n29335));
    SB_LUT4 add_3764_2_lut (.I0(GND_net), .I1(n50_adj_3998), .I2(n119_adj_3999), 
            .I3(GND_net), .O(n8344[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3764_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n23909), .I1(n7802[7]), .I2(n658), 
            .I3(n29333), .O(n3050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_10 (.CI(n29333), .I0(n7802[7]), .I1(n658), 
            .CO(n29334));
    SB_CARRY add_3764_2 (.CI(GND_net), .I0(n50_adj_3998), .I1(n119_adj_3999), 
            .CO(n29773));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n23909), .I1(n7802[6]), .I2(n585), 
            .I3(n29332), .O(n3050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3763_10_lut (.I0(GND_net), .I1(n8344[7]), .I2(n700_adj_4000), 
            .I3(n29772), .O(n8333[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3763_9_lut (.I0(GND_net), .I1(n8344[6]), .I2(n627_adj_4001), 
            .I3(n29771), .O(n8333[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_9 (.CI(n29771), .I0(n8344[6]), .I1(n627_adj_4001), 
            .CO(n29772));
    SB_LUT4 add_3763_8_lut (.I0(GND_net), .I1(n8344[5]), .I2(n554_adj_4002), 
            .I3(n29770), .O(n8333[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_8 (.CI(n29770), .I0(n8344[5]), .I1(n554_adj_4002), 
            .CO(n29771));
    SB_LUT4 add_3763_7_lut (.I0(GND_net), .I1(n8344[4]), .I2(n481_adj_4003), 
            .I3(n29769), .O(n8333[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_7 (.CI(n29769), .I0(n8344[4]), .I1(n481_adj_4003), 
            .CO(n29770));
    SB_LUT4 add_3763_6_lut (.I0(GND_net), .I1(n8344[3]), .I2(n408_adj_4004), 
            .I3(n29768), .O(n8333[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_6 (.CI(n29768), .I0(n8344[3]), .I1(n408_adj_4004), 
            .CO(n29769));
    SB_LUT4 add_3763_5_lut (.I0(GND_net), .I1(n8344[2]), .I2(n335_adj_4005), 
            .I3(n29767), .O(n8333[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_5 (.CI(n29767), .I0(n8344[2]), .I1(n335_adj_4005), 
            .CO(n29768));
    SB_LUT4 add_3763_4_lut (.I0(GND_net), .I1(n8344[1]), .I2(n262_adj_4006), 
            .I3(n29766), .O(n8333[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_4 (.CI(n29766), .I0(n8344[1]), .I1(n262_adj_4006), 
            .CO(n29767));
    SB_LUT4 add_3763_3_lut (.I0(GND_net), .I1(n8344[0]), .I2(n189_adj_4007), 
            .I3(n29765), .O(n8333[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_3 (.CI(n29765), .I0(n8344[0]), .I1(n189_adj_4007), 
            .CO(n29766));
    SB_LUT4 add_3763_2_lut (.I0(GND_net), .I1(n47_adj_4008), .I2(n116_adj_4009), 
            .I3(GND_net), .O(n8333[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3763_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3763_2 (.CI(GND_net), .I0(n47_adj_4008), .I1(n116_adj_4009), 
            .CO(n29765));
    SB_LUT4 add_3762_11_lut (.I0(GND_net), .I1(n8333[8]), .I2(n770_adj_4010), 
            .I3(n29764), .O(n8321[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3762_10_lut (.I0(GND_net), .I1(n8333[7]), .I2(n697_adj_4011), 
            .I3(n29763), .O(n8321[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_10 (.CI(n29763), .I0(n8333[7]), .I1(n697_adj_4011), 
            .CO(n29764));
    SB_LUT4 add_3762_9_lut (.I0(GND_net), .I1(n8333[6]), .I2(n624_adj_4012), 
            .I3(n29762), .O(n8321[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_9 (.CI(n29762), .I0(n8333[6]), .I1(n624_adj_4012), 
            .CO(n29763));
    SB_LUT4 add_3762_8_lut (.I0(GND_net), .I1(n8333[5]), .I2(n551_adj_4013), 
            .I3(n29761), .O(n8321[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_8 (.CI(n29761), .I0(n8333[5]), .I1(n551_adj_4013), 
            .CO(n29762));
    SB_LUT4 add_3762_7_lut (.I0(GND_net), .I1(n8333[4]), .I2(n478_adj_4014), 
            .I3(n29760), .O(n8321[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_7 (.CI(n29760), .I0(n8333[4]), .I1(n478_adj_4014), 
            .CO(n29761));
    SB_LUT4 add_3762_6_lut (.I0(GND_net), .I1(n8333[3]), .I2(n405_adj_4015), 
            .I3(n29759), .O(n8321[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_6 (.CI(n29759), .I0(n8333[3]), .I1(n405_adj_4015), 
            .CO(n29760));
    SB_CARRY mult_10_add_1225_9 (.CI(n29332), .I0(n7802[6]), .I1(n585), 
            .CO(n29333));
    SB_LUT4 add_3762_5_lut (.I0(GND_net), .I1(n8333[2]), .I2(n332_adj_4016), 
            .I3(n29758), .O(n8321[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n23909), .I1(n7802[5]), .I2(n512), 
            .I3(n29331), .O(n3050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3762_5 (.CI(n29758), .I0(n8333[2]), .I1(n332_adj_4016), 
            .CO(n29759));
    SB_LUT4 add_3762_4_lut (.I0(GND_net), .I1(n8333[1]), .I2(n259_adj_4017), 
            .I3(n29757), .O(n8321[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_4 (.CI(n29757), .I0(n8333[1]), .I1(n259_adj_4017), 
            .CO(n29758));
    SB_LUT4 add_3762_3_lut (.I0(GND_net), .I1(n8333[0]), .I2(n186_adj_4018), 
            .I3(n29756), .O(n8321[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_3 (.CI(n29756), .I0(n8333[0]), .I1(n186_adj_4018), 
            .CO(n29757));
    SB_LUT4 add_3762_2_lut (.I0(GND_net), .I1(n44_adj_4019), .I2(n113_adj_4020), 
            .I3(GND_net), .O(n8321[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3762_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3762_2 (.CI(GND_net), .I0(n44_adj_4019), .I1(n113_adj_4020), 
            .CO(n29756));
    SB_LUT4 add_3761_12_lut (.I0(GND_net), .I1(n8321[9]), .I2(n840_adj_4021), 
            .I3(n29755), .O(n8308[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3761_11_lut (.I0(GND_net), .I1(n8321[8]), .I2(n767_adj_4022), 
            .I3(n29754), .O(n8308[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_11 (.CI(n29754), .I0(n8321[8]), .I1(n767_adj_4022), 
            .CO(n29755));
    SB_LUT4 add_3761_10_lut (.I0(GND_net), .I1(n8321[7]), .I2(n694_adj_4023), 
            .I3(n29753), .O(n8308[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_10 (.CI(n29753), .I0(n8321[7]), .I1(n694_adj_4023), 
            .CO(n29754));
    SB_LUT4 add_3761_9_lut (.I0(GND_net), .I1(n8321[6]), .I2(n621_adj_4024), 
            .I3(n29752), .O(n8308[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_9 (.CI(n29752), .I0(n8321[6]), .I1(n621_adj_4024), 
            .CO(n29753));
    SB_LUT4 add_3761_8_lut (.I0(GND_net), .I1(n8321[5]), .I2(n548_adj_4025), 
            .I3(n29751), .O(n8308[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_8 (.CI(n29751), .I0(n8321[5]), .I1(n548_adj_4025), 
            .CO(n29752));
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13_adj_4026));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_3761_7_lut (.I0(GND_net), .I1(n8321[4]), .I2(n475_adj_4027), 
            .I3(n29750), .O(n8308[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n29331), .I0(n7802[5]), .I1(n512), 
            .CO(n29332));
    SB_CARRY add_3761_7 (.CI(n29750), .I0(n8321[4]), .I1(n475_adj_4027), 
            .CO(n29751));
    SB_LUT4 add_3761_6_lut (.I0(GND_net), .I1(n8321[3]), .I2(n402_adj_4028), 
            .I3(n29749), .O(n8308[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_6 (.CI(n29749), .I0(n8321[3]), .I1(n402_adj_4028), 
            .CO(n29750));
    SB_LUT4 add_3761_5_lut (.I0(GND_net), .I1(n8321[2]), .I2(n329_adj_4029), 
            .I3(n29748), .O(n8308[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_5 (.CI(n29748), .I0(n8321[2]), .I1(n329_adj_4029), 
            .CO(n29749));
    SB_LUT4 add_3761_4_lut (.I0(GND_net), .I1(n8321[1]), .I2(n256_adj_4030), 
            .I3(n29747), .O(n8308[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_4 (.CI(n29747), .I0(n8321[1]), .I1(n256_adj_4030), 
            .CO(n29748));
    SB_LUT4 add_3761_3_lut (.I0(GND_net), .I1(n8321[0]), .I2(n183_adj_4031), 
            .I3(n29746), .O(n8308[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3761_3 (.CI(n29746), .I0(n8321[0]), .I1(n183_adj_4031), 
            .CO(n29747));
    SB_LUT4 add_3761_2_lut (.I0(GND_net), .I1(n41_adj_4032), .I2(n110_adj_4033), 
            .I3(GND_net), .O(n8308[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3761_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4026), .I1(n18_adj_3994), .I2(n27550), 
            .I3(n4_adj_4034), .O(n36490));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3761_2 (.CI(GND_net), .I0(n41_adj_4032), .I1(n110_adj_4033), 
            .CO(n29746));
    SB_LUT4 add_3760_13_lut (.I0(GND_net), .I1(n8308[10]), .I2(n910_adj_4035), 
            .I3(n29745), .O(n8294[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3760_12_lut (.I0(GND_net), .I1(n8308[9]), .I2(n837_adj_4036), 
            .I3(n29744), .O(n8294[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_12 (.CI(n29744), .I0(n8308[9]), .I1(n837_adj_4036), 
            .CO(n29745));
    SB_LUT4 add_3760_11_lut (.I0(GND_net), .I1(n8308[8]), .I2(n764_adj_4037), 
            .I3(n29743), .O(n8294[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_11 (.CI(n29743), .I0(n8308[8]), .I1(n764_adj_4037), 
            .CO(n29744));
    SB_LUT4 add_3760_10_lut (.I0(GND_net), .I1(n8308[7]), .I2(n691_adj_4038), 
            .I3(n29742), .O(n8294[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_10 (.CI(n29742), .I0(n8308[7]), .I1(n691_adj_4038), 
            .CO(n29743));
    SB_LUT4 add_3760_9_lut (.I0(GND_net), .I1(n8308[6]), .I2(n618_adj_4039), 
            .I3(n29741), .O(n8294[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_9 (.CI(n29741), .I0(n8308[6]), .I1(n618_adj_4039), 
            .CO(n29742));
    SB_LUT4 add_3760_8_lut (.I0(GND_net), .I1(n8308[5]), .I2(n545_adj_4040), 
            .I3(n29740), .O(n8294[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_8 (.CI(n29740), .I0(n8308[5]), .I1(n545_adj_4040), 
            .CO(n29741));
    SB_LUT4 add_3760_7_lut (.I0(GND_net), .I1(n8308[4]), .I2(n472_adj_4041), 
            .I3(n29739), .O(n8294[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_7 (.CI(n29739), .I0(n8308[4]), .I1(n472_adj_4041), 
            .CO(n29740));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n23909), .I1(n7802[4]), .I2(n439), 
            .I3(n29330), .O(n3050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3760_6_lut (.I0(GND_net), .I1(n8308[3]), .I2(n399_adj_4042), 
            .I3(n29738), .O(n8294[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_6 (.CI(n29738), .I0(n8308[3]), .I1(n399_adj_4042), 
            .CO(n29739));
    SB_LUT4 add_3760_5_lut (.I0(GND_net), .I1(n8308[2]), .I2(n326_adj_4043), 
            .I3(n29737), .O(n8294[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_5 (.CI(n29737), .I0(n8308[2]), .I1(n326_adj_4043), 
            .CO(n29738));
    SB_LUT4 add_3760_4_lut (.I0(GND_net), .I1(n8308[1]), .I2(n253_adj_4044), 
            .I3(n29736), .O(n8294[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_4 (.CI(n29736), .I0(n8308[1]), .I1(n253_adj_4044), 
            .CO(n29737));
    SB_LUT4 add_3760_3_lut (.I0(GND_net), .I1(n8308[0]), .I2(n180_adj_4045), 
            .I3(n29735), .O(n8294[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3760_3 (.CI(n29735), .I0(n8308[0]), .I1(n180_adj_4045), 
            .CO(n29736));
    SB_LUT4 add_3760_2_lut (.I0(GND_net), .I1(n38_adj_4046), .I2(n107_adj_4047), 
            .I3(GND_net), .O(n8294[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3760_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n29330), .I0(n7802[4]), .I1(n439), 
            .CO(n29331));
    SB_CARRY add_3760_2 (.CI(GND_net), .I0(n38_adj_4046), .I1(n107_adj_4047), 
            .CO(n29735));
    SB_LUT4 add_3759_14_lut (.I0(GND_net), .I1(n8294[11]), .I2(n980_adj_4048), 
            .I3(n29734), .O(n8279[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4049));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4050));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3759_13_lut (.I0(GND_net), .I1(n8294[10]), .I2(n907_adj_4051), 
            .I3(n29733), .O(n8279[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_13 (.CI(n29733), .I0(n8294[10]), .I1(n907_adj_4051), 
            .CO(n29734));
    SB_LUT4 add_3759_12_lut (.I0(GND_net), .I1(n8294[9]), .I2(n834_adj_4052), 
            .I3(n29732), .O(n8279[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_12 (.CI(n29732), .I0(n8294[9]), .I1(n834_adj_4052), 
            .CO(n29733));
    SB_LUT4 add_3759_11_lut (.I0(GND_net), .I1(n8294[8]), .I2(n761_adj_4053), 
            .I3(n29731), .O(n8279[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_11 (.CI(n29731), .I0(n8294[8]), .I1(n761_adj_4053), 
            .CO(n29732));
    SB_LUT4 add_3759_10_lut (.I0(GND_net), .I1(n8294[7]), .I2(n688_adj_4054), 
            .I3(n29730), .O(n8279[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_10 (.CI(n29730), .I0(n8294[7]), .I1(n688_adj_4054), 
            .CO(n29731));
    SB_LUT4 add_3759_9_lut (.I0(GND_net), .I1(n8294[6]), .I2(n615_adj_4055), 
            .I3(n29729), .O(n8279[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_9 (.CI(n29729), .I0(n8294[6]), .I1(n615_adj_4055), 
            .CO(n29730));
    SB_LUT4 add_3759_8_lut (.I0(GND_net), .I1(n8294[5]), .I2(n542_adj_4056), 
            .I3(n29728), .O(n8279[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_8 (.CI(n29728), .I0(n8294[5]), .I1(n542_adj_4056), 
            .CO(n29729));
    SB_LUT4 add_3759_7_lut (.I0(GND_net), .I1(n8294[4]), .I2(n469_adj_4057), 
            .I3(n29727), .O(n8279[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_7 (.CI(n29727), .I0(n8294[4]), .I1(n469_adj_4057), 
            .CO(n29728));
    SB_LUT4 add_3759_6_lut (.I0(GND_net), .I1(n8294[3]), .I2(n396_adj_4058), 
            .I3(n29726), .O(n8279[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_6 (.CI(n29726), .I0(n8294[3]), .I1(n396_adj_4058), 
            .CO(n29727));
    SB_LUT4 add_3759_5_lut (.I0(GND_net), .I1(n8294[2]), .I2(n323_adj_4059), 
            .I3(n29725), .O(n8279[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_5 (.CI(n29725), .I0(n8294[2]), .I1(n323_adj_4059), 
            .CO(n29726));
    SB_LUT4 add_3759_4_lut (.I0(GND_net), .I1(n8294[1]), .I2(n250_adj_4060), 
            .I3(n29724), .O(n8279[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_4 (.CI(n29724), .I0(n8294[1]), .I1(n250_adj_4060), 
            .CO(n29725));
    SB_LUT4 add_3759_3_lut (.I0(GND_net), .I1(n8294[0]), .I2(n177_adj_4061), 
            .I3(n29723), .O(n8279[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_3 (.CI(n29723), .I0(n8294[0]), .I1(n177_adj_4061), 
            .CO(n29724));
    SB_LUT4 add_3759_2_lut (.I0(GND_net), .I1(n35_adj_4062), .I2(n104_adj_4063), 
            .I3(GND_net), .O(n8279[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3759_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3759_2 (.CI(GND_net), .I0(n35_adj_4062), .I1(n104_adj_4063), 
            .CO(n29723));
    SB_LUT4 add_3758_15_lut (.I0(GND_net), .I1(n8279[12]), .I2(n1050_adj_4064), 
            .I3(n29722), .O(n8263[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3758_14_lut (.I0(GND_net), .I1(n8279[11]), .I2(n977_adj_4065), 
            .I3(n29721), .O(n8263[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n23909), .I1(n7802[3]), .I2(n366), 
            .I3(n29329), .O(n3050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_6 (.CI(n29329), .I0(n7802[3]), .I1(n366), 
            .CO(n29330));
    SB_CARRY add_3758_14 (.CI(n29721), .I0(n8279[11]), .I1(n977_adj_4065), 
            .CO(n29722));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n23909), .I1(n7802[2]), .I2(n293), 
            .I3(n29328), .O(n3050[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3758_13_lut (.I0(GND_net), .I1(n8279[10]), .I2(n904_adj_4066), 
            .I3(n29720), .O(n8263[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3758_13 (.CI(n29720), .I0(n8279[10]), .I1(n904_adj_4066), 
            .CO(n29721));
    SB_LUT4 add_3758_12_lut (.I0(GND_net), .I1(n8279[9]), .I2(n831_adj_4068), 
            .I3(n29719), .O(n8263[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_12 (.CI(n29719), .I0(n8279[9]), .I1(n831_adj_4068), 
            .CO(n29720));
    SB_LUT4 add_3758_11_lut (.I0(GND_net), .I1(n8279[8]), .I2(n758_adj_4069), 
            .I3(n29718), .O(n8263[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n29328), .I0(n7802[2]), .I1(n293), 
            .CO(n29329));
    SB_CARRY add_3758_11 (.CI(n29718), .I0(n8279[8]), .I1(n758_adj_4069), 
            .CO(n29719));
    SB_LUT4 add_3758_10_lut (.I0(GND_net), .I1(n8279[7]), .I2(n685_adj_4070), 
            .I3(n29717), .O(n8263[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_10 (.CI(n29717), .I0(n8279[7]), .I1(n685_adj_4070), 
            .CO(n29718));
    SB_LUT4 add_3758_9_lut (.I0(GND_net), .I1(n8279[6]), .I2(n612_adj_4071), 
            .I3(n29716), .O(n8263[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_9 (.CI(n29716), .I0(n8279[6]), .I1(n612_adj_4071), 
            .CO(n29717));
    SB_LUT4 add_3758_8_lut (.I0(GND_net), .I1(n8279[5]), .I2(n539_adj_4072), 
            .I3(n29715), .O(n8263[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_8 (.CI(n29715), .I0(n8279[5]), .I1(n539_adj_4072), 
            .CO(n29716));
    SB_LUT4 add_3758_7_lut (.I0(GND_net), .I1(n8279[4]), .I2(n466_adj_4073), 
            .I3(n29714), .O(n8263[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_7 (.CI(n29714), .I0(n8279[4]), .I1(n466_adj_4073), 
            .CO(n29715));
    SB_LUT4 add_3758_6_lut (.I0(GND_net), .I1(n8279[3]), .I2(n393_adj_4074), 
            .I3(n29713), .O(n8263[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_6 (.CI(n29713), .I0(n8279[3]), .I1(n393_adj_4074), 
            .CO(n29714));
    SB_LUT4 add_3758_5_lut (.I0(GND_net), .I1(n8279[2]), .I2(n320_adj_4075), 
            .I3(n29712), .O(n8263[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_5 (.CI(n29712), .I0(n8279[2]), .I1(n320_adj_4075), 
            .CO(n29713));
    SB_LUT4 add_3758_4_lut (.I0(GND_net), .I1(n8279[1]), .I2(n247_adj_4076), 
            .I3(n29711), .O(n8263[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n23909), .I1(n7802[1]), .I2(n220), 
            .I3(n29327), .O(n3050[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_4 (.CI(n29327), .I0(n7802[1]), .I1(n220), 
            .CO(n29328));
    SB_CARRY add_3758_4 (.CI(n29711), .I0(n8279[1]), .I1(n247_adj_4076), 
            .CO(n29712));
    SB_LUT4 add_3758_3_lut (.I0(GND_net), .I1(n8279[0]), .I2(n174_adj_4077), 
            .I3(n29710), .O(n8263[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_3 (.CI(n29710), .I0(n8279[0]), .I1(n174_adj_4077), 
            .CO(n29711));
    SB_LUT4 add_3758_2_lut (.I0(GND_net), .I1(n32_adj_4078), .I2(n101_adj_4079), 
            .I3(GND_net), .O(n8263[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3758_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3758_2 (.CI(GND_net), .I0(n32_adj_4078), .I1(n101_adj_4079), 
            .CO(n29710));
    SB_LUT4 add_3757_16_lut (.I0(GND_net), .I1(n8263[13]), .I2(n1120_adj_4080), 
            .I3(n29709), .O(n8246[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3757_15_lut (.I0(GND_net), .I1(n8263[12]), .I2(n1047_adj_4081), 
            .I3(n29708), .O(n8246[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_15 (.CI(n29708), .I0(n8263[12]), .I1(n1047_adj_4081), 
            .CO(n29709));
    SB_LUT4 add_3757_14_lut (.I0(GND_net), .I1(n8263[11]), .I2(n974_adj_4082), 
            .I3(n29707), .O(n8246[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_14 (.CI(n29707), .I0(n8263[11]), .I1(n974_adj_4082), 
            .CO(n29708));
    SB_LUT4 add_3757_13_lut (.I0(GND_net), .I1(n8263[10]), .I2(n901_adj_4083), 
            .I3(n29706), .O(n8246[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_13 (.CI(n29706), .I0(n8263[10]), .I1(n901_adj_4083), 
            .CO(n29707));
    SB_LUT4 add_3757_12_lut (.I0(GND_net), .I1(n8263[9]), .I2(n828_adj_4084), 
            .I3(n29705), .O(n8246[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_12 (.CI(n29705), .I0(n8263[9]), .I1(n828_adj_4084), 
            .CO(n29706));
    SB_LUT4 add_3757_11_lut (.I0(GND_net), .I1(n8263[8]), .I2(n755_adj_4085), 
            .I3(n29704), .O(n8246[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_11 (.CI(n29704), .I0(n8263[8]), .I1(n755_adj_4085), 
            .CO(n29705));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n23909), .I1(n7802[0]), .I2(n147), 
            .I3(n29326), .O(n3050[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3757_10_lut (.I0(GND_net), .I1(n8263[7]), .I2(n682_adj_4086), 
            .I3(n29703), .O(n8246[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_10 (.CI(n29703), .I0(n8263[7]), .I1(n682_adj_4086), 
            .CO(n29704));
    SB_LUT4 add_3757_9_lut (.I0(GND_net), .I1(n8263[6]), .I2(n609_adj_4087), 
            .I3(n29702), .O(n8246[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_9 (.CI(n29702), .I0(n8263[6]), .I1(n609_adj_4087), 
            .CO(n29703));
    SB_LUT4 add_3757_8_lut (.I0(GND_net), .I1(n8263[5]), .I2(n536_adj_4088), 
            .I3(n29701), .O(n8246[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_8 (.CI(n29701), .I0(n8263[5]), .I1(n536_adj_4088), 
            .CO(n29702));
    SB_LUT4 add_3757_7_lut (.I0(GND_net), .I1(n8263[4]), .I2(n463_adj_4089), 
            .I3(n29700), .O(n8246[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n29326), .I0(n7802[0]), .I1(n147), 
            .CO(n29327));
    SB_CARRY add_3757_7 (.CI(n29700), .I0(n8263[4]), .I1(n463_adj_4089), 
            .CO(n29701));
    SB_LUT4 add_3757_6_lut (.I0(GND_net), .I1(n8263[3]), .I2(n390_adj_4090), 
            .I3(n29699), .O(n8246[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_6 (.CI(n29699), .I0(n8263[3]), .I1(n390_adj_4090), 
            .CO(n29700));
    SB_LUT4 add_3757_5_lut (.I0(GND_net), .I1(n8263[2]), .I2(n317_adj_4091), 
            .I3(n29698), .O(n8246[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_5 (.CI(n29698), .I0(n8263[2]), .I1(n317_adj_4091), 
            .CO(n29699));
    SB_LUT4 add_3757_4_lut (.I0(GND_net), .I1(n8263[1]), .I2(n244_adj_4092), 
            .I3(n29697), .O(n8246[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3757_4 (.CI(n29697), .I0(n8263[1]), .I1(n244_adj_4092), 
            .CO(n29698));
    SB_LUT4 add_3757_3_lut (.I0(GND_net), .I1(n8263[0]), .I2(n171_adj_4093), 
            .I3(n29696), .O(n8246[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n23909), .I1(n5_adj_4094), .I2(n74), 
            .I3(GND_net), .O(n3050[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3757_3 (.CI(n29696), .I0(n8263[0]), .I1(n171_adj_4093), 
            .CO(n29697));
    SB_LUT4 add_3757_2_lut (.I0(GND_net), .I1(n29_adj_4095), .I2(n98_adj_4096), 
            .I3(GND_net), .O(n8246[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3757_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4094), .I1(n74), 
            .CO(n29326));
    SB_CARRY add_3757_2 (.CI(GND_net), .I0(n29_adj_4095), .I1(n98_adj_4096), 
            .CO(n29696));
    SB_LUT4 add_3756_17_lut (.I0(GND_net), .I1(n8246[14]), .I2(GND_net), 
            .I3(n29695), .O(n8228[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3756_16_lut (.I0(GND_net), .I1(n8246[13]), .I2(n1117_adj_4097), 
            .I3(n29694), .O(n8228[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_16 (.CI(n29694), .I0(n8246[13]), .I1(n1117_adj_4097), 
            .CO(n29695));
    SB_LUT4 add_3728_23_lut (.I0(GND_net), .I1(n7826[20]), .I2(GND_net), 
            .I3(n29325), .O(n7802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3756_15_lut (.I0(GND_net), .I1(n8246[12]), .I2(n1044_adj_4098), 
            .I3(n29693), .O(n8228[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_15 (.CI(n29693), .I0(n8246[12]), .I1(n1044_adj_4098), 
            .CO(n29694));
    SB_LUT4 add_3756_14_lut (.I0(GND_net), .I1(n8246[11]), .I2(n971_adj_4099), 
            .I3(n29692), .O(n8228[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_14 (.CI(n29692), .I0(n8246[11]), .I1(n971_adj_4099), 
            .CO(n29693));
    SB_LUT4 add_3756_13_lut (.I0(GND_net), .I1(n8246[10]), .I2(n898_adj_4100), 
            .I3(n29691), .O(n8228[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_13 (.CI(n29691), .I0(n8246[10]), .I1(n898_adj_4100), 
            .CO(n29692));
    SB_LUT4 add_3756_12_lut (.I0(GND_net), .I1(n8246[9]), .I2(n825_adj_4101), 
            .I3(n29690), .O(n8228[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_12 (.CI(n29690), .I0(n8246[9]), .I1(n825_adj_4101), 
            .CO(n29691));
    SB_LUT4 add_3756_11_lut (.I0(GND_net), .I1(n8246[8]), .I2(n752_adj_4102), 
            .I3(n29689), .O(n8228[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_11 (.CI(n29689), .I0(n8246[8]), .I1(n752_adj_4102), 
            .CO(n29690));
    SB_LUT4 add_3756_10_lut (.I0(GND_net), .I1(n8246[7]), .I2(n679_adj_4103), 
            .I3(n29688), .O(n8228[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_10 (.CI(n29688), .I0(n8246[7]), .I1(n679_adj_4103), 
            .CO(n29689));
    SB_LUT4 add_3756_9_lut (.I0(GND_net), .I1(n8246[6]), .I2(n606_adj_4104), 
            .I3(n29687), .O(n8228[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_9 (.CI(n29687), .I0(n8246[6]), .I1(n606_adj_4104), 
            .CO(n29688));
    SB_LUT4 add_3756_8_lut (.I0(GND_net), .I1(n8246[5]), .I2(n533_adj_4105), 
            .I3(n29686), .O(n8228[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_8 (.CI(n29686), .I0(n8246[5]), .I1(n533_adj_4105), 
            .CO(n29687));
    SB_LUT4 add_3756_7_lut (.I0(GND_net), .I1(n8246[4]), .I2(n460_adj_4106), 
            .I3(n29685), .O(n8228[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_7 (.CI(n29685), .I0(n8246[4]), .I1(n460_adj_4106), 
            .CO(n29686));
    SB_LUT4 add_3756_6_lut (.I0(GND_net), .I1(n8246[3]), .I2(n387_adj_4107), 
            .I3(n29684), .O(n8228[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_6 (.CI(n29684), .I0(n8246[3]), .I1(n387_adj_4107), 
            .CO(n29685));
    SB_LUT4 add_3728_22_lut (.I0(GND_net), .I1(n7826[19]), .I2(GND_net), 
            .I3(n29324), .O(n7802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3756_5_lut (.I0(GND_net), .I1(n8246[2]), .I2(n314_adj_4108), 
            .I3(n29683), .O(n8228[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_5 (.CI(n29683), .I0(n8246[2]), .I1(n314_adj_4108), 
            .CO(n29684));
    SB_LUT4 add_3756_4_lut (.I0(GND_net), .I1(n8246[1]), .I2(n241_adj_4109), 
            .I3(n29682), .O(n8228[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_4 (.CI(n29682), .I0(n8246[1]), .I1(n241_adj_4109), 
            .CO(n29683));
    SB_LUT4 add_3756_3_lut (.I0(GND_net), .I1(n8246[0]), .I2(n168_adj_4110), 
            .I3(n29681), .O(n8228[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_3 (.CI(n29681), .I0(n8246[0]), .I1(n168_adj_4110), 
            .CO(n29682));
    SB_LUT4 add_3756_2_lut (.I0(GND_net), .I1(n26_adj_4111), .I2(n95_adj_4112), 
            .I3(GND_net), .O(n8228[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3756_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3756_2 (.CI(GND_net), .I0(n26_adj_4111), .I1(n95_adj_4112), 
            .CO(n29681));
    SB_LUT4 add_3755_18_lut (.I0(GND_net), .I1(n8228[15]), .I2(GND_net), 
            .I3(n29680), .O(n8209[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_22 (.CI(n29324), .I0(n7826[19]), .I1(GND_net), .CO(n29325));
    SB_LUT4 add_3755_17_lut (.I0(GND_net), .I1(n8228[14]), .I2(GND_net), 
            .I3(n29679), .O(n8209[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_17 (.CI(n29679), .I0(n8228[14]), .I1(GND_net), .CO(n29680));
    SB_LUT4 add_3755_16_lut (.I0(GND_net), .I1(n8228[13]), .I2(n1114_adj_4113), 
            .I3(n29678), .O(n8209[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_16 (.CI(n29678), .I0(n8228[13]), .I1(n1114_adj_4113), 
            .CO(n29679));
    SB_LUT4 add_3755_15_lut (.I0(GND_net), .I1(n8228[12]), .I2(n1041_adj_4114), 
            .I3(n29677), .O(n8209[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_15 (.CI(n29677), .I0(n8228[12]), .I1(n1041_adj_4114), 
            .CO(n29678));
    SB_LUT4 add_3755_14_lut (.I0(GND_net), .I1(n8228[11]), .I2(n968_adj_4115), 
            .I3(n29676), .O(n8209[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_14 (.CI(n29676), .I0(n8228[11]), .I1(n968_adj_4115), 
            .CO(n29677));
    SB_LUT4 add_3755_13_lut (.I0(GND_net), .I1(n8228[10]), .I2(n895_adj_4116), 
            .I3(n29675), .O(n8209[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_13 (.CI(n29675), .I0(n8228[10]), .I1(n895_adj_4116), 
            .CO(n29676));
    SB_LUT4 add_3755_12_lut (.I0(GND_net), .I1(n8228[9]), .I2(n822_adj_4117), 
            .I3(n29674), .O(n8209[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_12 (.CI(n29674), .I0(n8228[9]), .I1(n822_adj_4117), 
            .CO(n29675));
    SB_LUT4 add_3755_11_lut (.I0(GND_net), .I1(n8228[8]), .I2(n749_adj_4118), 
            .I3(n29673), .O(n8209[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_11 (.CI(n29673), .I0(n8228[8]), .I1(n749_adj_4118), 
            .CO(n29674));
    SB_LUT4 add_3755_10_lut (.I0(GND_net), .I1(n8228[7]), .I2(n676_adj_4119), 
            .I3(n29672), .O(n8209[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_10 (.CI(n29672), .I0(n8228[7]), .I1(n676_adj_4119), 
            .CO(n29673));
    SB_LUT4 add_3755_9_lut (.I0(GND_net), .I1(n8228[6]), .I2(n603_adj_4120), 
            .I3(n29671), .O(n8209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_9 (.CI(n29671), .I0(n8228[6]), .I1(n603_adj_4120), 
            .CO(n29672));
    SB_LUT4 add_3728_21_lut (.I0(GND_net), .I1(n7826[18]), .I2(GND_net), 
            .I3(n29323), .O(n7802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3755_8_lut (.I0(GND_net), .I1(n8228[5]), .I2(n530_adj_4121), 
            .I3(n29670), .O(n8209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_8 (.CI(n29670), .I0(n8228[5]), .I1(n530_adj_4121), 
            .CO(n29671));
    SB_LUT4 add_3755_7_lut (.I0(GND_net), .I1(n8228[4]), .I2(n457_adj_4122), 
            .I3(n29669), .O(n8209[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_7 (.CI(n29669), .I0(n8228[4]), .I1(n457_adj_4122), 
            .CO(n29670));
    SB_LUT4 add_3755_6_lut (.I0(GND_net), .I1(n8228[3]), .I2(n384_adj_4123), 
            .I3(n29668), .O(n8209[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_6 (.CI(n29668), .I0(n8228[3]), .I1(n384_adj_4123), 
            .CO(n29669));
    SB_LUT4 add_3755_5_lut (.I0(GND_net), .I1(n8228[2]), .I2(n311_adj_4124), 
            .I3(n29667), .O(n8209[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_5 (.CI(n29667), .I0(n8228[2]), .I1(n311_adj_4124), 
            .CO(n29668));
    SB_LUT4 add_3755_4_lut (.I0(GND_net), .I1(n8228[1]), .I2(n238_adj_4125), 
            .I3(n29666), .O(n8209[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_4 (.CI(n29666), .I0(n8228[1]), .I1(n238_adj_4125), 
            .CO(n29667));
    SB_LUT4 add_3755_3_lut (.I0(GND_net), .I1(n8228[0]), .I2(n165_adj_4126), 
            .I3(n29665), .O(n8209[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_3 (.CI(n29665), .I0(n8228[0]), .I1(n165_adj_4126), 
            .CO(n29666));
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4127));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3755_2_lut (.I0(GND_net), .I1(n23_adj_4128), .I2(n92_adj_4129), 
            .I3(GND_net), .O(n8209[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3755_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3755_2 (.CI(GND_net), .I0(n23_adj_4128), .I1(n92_adj_4129), 
            .CO(n29665));
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4130));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4131));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3754_19_lut (.I0(GND_net), .I1(n8209[16]), .I2(GND_net), 
            .I3(n29664), .O(n8189[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3754_18_lut (.I0(GND_net), .I1(n8209[15]), .I2(GND_net), 
            .I3(n29663), .O(n8189[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_18 (.CI(n29663), .I0(n8209[15]), .I1(GND_net), .CO(n29664));
    SB_LUT4 add_3754_17_lut (.I0(GND_net), .I1(n8209[14]), .I2(GND_net), 
            .I3(n29662), .O(n8189[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_17 (.CI(n29662), .I0(n8209[14]), .I1(GND_net), .CO(n29663));
    SB_LUT4 add_3754_16_lut (.I0(GND_net), .I1(n8209[13]), .I2(n1111_adj_4132), 
            .I3(n29661), .O(n8189[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_16 (.CI(n29661), .I0(n8209[13]), .I1(n1111_adj_4132), 
            .CO(n29662));
    SB_LUT4 add_3754_15_lut (.I0(GND_net), .I1(n8209[12]), .I2(n1038_adj_4133), 
            .I3(n29660), .O(n8189[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_15 (.CI(n29660), .I0(n8209[12]), .I1(n1038_adj_4133), 
            .CO(n29661));
    SB_LUT4 add_3754_14_lut (.I0(GND_net), .I1(n8209[11]), .I2(n965_adj_4134), 
            .I3(n29659), .O(n8189[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_14 (.CI(n29659), .I0(n8209[11]), .I1(n965_adj_4134), 
            .CO(n29660));
    SB_LUT4 add_3754_13_lut (.I0(GND_net), .I1(n8209[10]), .I2(n892_adj_4135), 
            .I3(n29658), .O(n8189[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_13 (.CI(n29658), .I0(n8209[10]), .I1(n892_adj_4135), 
            .CO(n29659));
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4136));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3754_12_lut (.I0(GND_net), .I1(n8209[9]), .I2(n819_adj_4137), 
            .I3(n29657), .O(n8189[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_12 (.CI(n29657), .I0(n8209[9]), .I1(n819_adj_4137), 
            .CO(n29658));
    SB_LUT4 add_3754_11_lut (.I0(GND_net), .I1(n8209[8]), .I2(n746_adj_4138), 
            .I3(n29656), .O(n8189[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_11 (.CI(n29656), .I0(n8209[8]), .I1(n746_adj_4138), 
            .CO(n29657));
    SB_LUT4 add_3754_10_lut (.I0(GND_net), .I1(n8209[7]), .I2(n673_adj_4139), 
            .I3(n29655), .O(n8189[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_10 (.CI(n29655), .I0(n8209[7]), .I1(n673_adj_4139), 
            .CO(n29656));
    SB_LUT4 add_3754_9_lut (.I0(GND_net), .I1(n8209[6]), .I2(n600_adj_4140), 
            .I3(n29654), .O(n8189[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_9 (.CI(n29654), .I0(n8209[6]), .I1(n600_adj_4140), 
            .CO(n29655));
    SB_LUT4 add_3754_8_lut (.I0(GND_net), .I1(n8209[5]), .I2(n527_adj_4141), 
            .I3(n29653), .O(n8189[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_8 (.CI(n29653), .I0(n8209[5]), .I1(n527_adj_4141), 
            .CO(n29654));
    SB_LUT4 add_3754_7_lut (.I0(GND_net), .I1(n8209[4]), .I2(n454_adj_4142), 
            .I3(n29652), .O(n8189[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4143));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3754_7 (.CI(n29652), .I0(n8209[4]), .I1(n454_adj_4142), 
            .CO(n29653));
    SB_LUT4 add_3754_6_lut (.I0(GND_net), .I1(n8209[3]), .I2(n381_adj_4144), 
            .I3(n29651), .O(n8189[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_6 (.CI(n29651), .I0(n8209[3]), .I1(n381_adj_4144), 
            .CO(n29652));
    SB_LUT4 add_3754_5_lut (.I0(GND_net), .I1(n8209[2]), .I2(n308_adj_4145), 
            .I3(n29650), .O(n8189[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_5 (.CI(n29650), .I0(n8209[2]), .I1(n308_adj_4145), 
            .CO(n29651));
    SB_LUT4 add_3754_4_lut (.I0(GND_net), .I1(n8209[1]), .I2(n235_adj_4146), 
            .I3(n29649), .O(n8189[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_4 (.CI(n29649), .I0(n8209[1]), .I1(n235_adj_4146), 
            .CO(n29650));
    SB_LUT4 add_3754_3_lut (.I0(GND_net), .I1(n8209[0]), .I2(n162_adj_4147), 
            .I3(n29648), .O(n8189[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_3 (.CI(n29648), .I0(n8209[0]), .I1(n162_adj_4147), 
            .CO(n29649));
    SB_LUT4 add_3754_2_lut (.I0(GND_net), .I1(n20_adj_4148), .I2(n89_adj_4149), 
            .I3(GND_net), .O(n8189[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3754_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3754_2 (.CI(GND_net), .I0(n20_adj_4148), .I1(n89_adj_4149), 
            .CO(n29648));
    SB_LUT4 add_3753_20_lut (.I0(GND_net), .I1(n8189[17]), .I2(GND_net), 
            .I3(n29647), .O(n8168[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22838_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n27491), .I3(n8087[0]), .O(n4_adj_3970));   // verilog/motorControl.v(42[17:23])
    defparam i22838_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_3753_19_lut (.I0(GND_net), .I1(n8189[16]), .I2(GND_net), 
            .I3(n29646), .O(n8168[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_21 (.CI(n29323), .I0(n7826[18]), .I1(GND_net), .CO(n29324));
    SB_CARRY add_3753_19 (.CI(n29646), .I0(n8189[16]), .I1(GND_net), .CO(n29647));
    SB_LUT4 add_3753_18_lut (.I0(GND_net), .I1(n8189[15]), .I2(GND_net), 
            .I3(n29645), .O(n8168[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_978 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n8087[0]), .I3(n27491), .O(n8081[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_978.LUT_INIT = 16'h8778;
    SB_CARRY add_3753_18 (.CI(n29645), .I0(n8189[15]), .I1(GND_net), .CO(n29646));
    SB_LUT4 add_3753_17_lut (.I0(GND_net), .I1(n8189[14]), .I2(GND_net), 
            .I3(n29644), .O(n8168[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22869_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n27525), .I3(n8092[0]), .O(n4_adj_4034));   // verilog/motorControl.v(42[17:23])
    defparam i22869_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_3753_17 (.CI(n29644), .I0(n8189[14]), .I1(GND_net), .CO(n29645));
    SB_LUT4 add_3753_16_lut (.I0(GND_net), .I1(n8189[13]), .I2(n1108_adj_4150), 
            .I3(n29643), .O(n8168[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_16 (.CI(n29643), .I0(n8189[13]), .I1(n1108_adj_4150), 
            .CO(n29644));
    SB_LUT4 add_3753_15_lut (.I0(GND_net), .I1(n8189[12]), .I2(n1035_adj_4151), 
            .I3(n29642), .O(n8168[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_15 (.CI(n29642), .I0(n8189[12]), .I1(n1035_adj_4151), 
            .CO(n29643));
    SB_LUT4 add_3753_14_lut (.I0(GND_net), .I1(n8189[11]), .I2(n962_adj_4152), 
            .I3(n29641), .O(n8168[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_14 (.CI(n29641), .I0(n8189[11]), .I1(n962_adj_4152), 
            .CO(n29642));
    SB_LUT4 add_3753_13_lut (.I0(GND_net), .I1(n8189[10]), .I2(n889_adj_4153), 
            .I3(n29640), .O(n8168[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_13 (.CI(n29640), .I0(n8189[10]), .I1(n889_adj_4153), 
            .CO(n29641));
    SB_LUT4 add_3753_12_lut (.I0(GND_net), .I1(n8189[9]), .I2(n816_adj_4154), 
            .I3(n29639), .O(n8168[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_12 (.CI(n29639), .I0(n8189[9]), .I1(n816_adj_4154), 
            .CO(n29640));
    SB_LUT4 add_3753_11_lut (.I0(GND_net), .I1(n8189[8]), .I2(n743_adj_4155), 
            .I3(n29638), .O(n8168[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_20_lut (.I0(GND_net), .I1(n7826[17]), .I2(GND_net), 
            .I3(n29322), .O(n7802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_11 (.CI(n29638), .I0(n8189[8]), .I1(n743_adj_4155), 
            .CO(n29639));
    SB_LUT4 add_3753_10_lut (.I0(GND_net), .I1(n8189[7]), .I2(n670_adj_4156), 
            .I3(n29637), .O(n8168[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_10 (.CI(n29637), .I0(n8189[7]), .I1(n670_adj_4156), 
            .CO(n29638));
    SB_LUT4 add_3753_9_lut (.I0(GND_net), .I1(n8189[6]), .I2(n597_adj_4157), 
            .I3(n29636), .O(n8168[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_9 (.CI(n29636), .I0(n8189[6]), .I1(n597_adj_4157), 
            .CO(n29637));
    SB_LUT4 add_3753_8_lut (.I0(GND_net), .I1(n8189[5]), .I2(n524_adj_4158), 
            .I3(n29635), .O(n8168[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_8 (.CI(n29635), .I0(n8189[5]), .I1(n524_adj_4158), 
            .CO(n29636));
    SB_LUT4 add_3753_7_lut (.I0(GND_net), .I1(n8189[4]), .I2(n451_adj_4159), 
            .I3(n29634), .O(n8168[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_7 (.CI(n29634), .I0(n8189[4]), .I1(n451_adj_4159), 
            .CO(n29635));
    SB_LUT4 add_3753_6_lut (.I0(GND_net), .I1(n8189[3]), .I2(n378_adj_4160), 
            .I3(n29633), .O(n8168[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_6 (.CI(n29633), .I0(n8189[3]), .I1(n378_adj_4160), 
            .CO(n29634));
    SB_LUT4 add_3753_5_lut (.I0(GND_net), .I1(n8189[2]), .I2(n305_adj_4161), 
            .I3(n29632), .O(n8168[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_5 (.CI(n29632), .I0(n8189[2]), .I1(n305_adj_4161), 
            .CO(n29633));
    SB_LUT4 add_3753_4_lut (.I0(GND_net), .I1(n8189[1]), .I2(n232_adj_4162), 
            .I3(n29631), .O(n8168[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_4 (.CI(n29631), .I0(n8189[1]), .I1(n232_adj_4162), 
            .CO(n29632));
    SB_LUT4 add_3753_3_lut (.I0(GND_net), .I1(n8189[0]), .I2(n159_adj_4163), 
            .I3(n29630), .O(n8168[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_20 (.CI(n29322), .I0(n7826[17]), .I1(GND_net), .CO(n29323));
    SB_CARRY add_3753_3 (.CI(n29630), .I0(n8189[0]), .I1(n159_adj_4163), 
            .CO(n29631));
    SB_LUT4 add_3753_2_lut (.I0(GND_net), .I1(n17_adj_4164), .I2(n86_adj_4165), 
            .I3(GND_net), .O(n8168[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3753_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3753_2 (.CI(GND_net), .I0(n17_adj_4164), .I1(n86_adj_4165), 
            .CO(n29630));
    SB_LUT4 add_3752_21_lut (.I0(GND_net), .I1(n8168[18]), .I2(GND_net), 
            .I3(n29629), .O(n8146[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_20_lut (.I0(GND_net), .I1(n8168[17]), .I2(GND_net), 
            .I3(n29628), .O(n8146[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_20 (.CI(n29628), .I0(n8168[17]), .I1(GND_net), .CO(n29629));
    SB_LUT4 add_3752_19_lut (.I0(GND_net), .I1(n8168[16]), .I2(GND_net), 
            .I3(n29627), .O(n8146[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_19 (.CI(n29627), .I0(n8168[16]), .I1(GND_net), .CO(n29628));
    SB_LUT4 add_3752_18_lut (.I0(GND_net), .I1(n8168[15]), .I2(GND_net), 
            .I3(n29626), .O(n8146[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_18 (.CI(n29626), .I0(n8168[15]), .I1(GND_net), .CO(n29627));
    SB_LUT4 add_3752_17_lut (.I0(GND_net), .I1(n8168[14]), .I2(GND_net), 
            .I3(n29625), .O(n8146[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_17 (.CI(n29625), .I0(n8168[14]), .I1(GND_net), .CO(n29626));
    SB_LUT4 add_3752_16_lut (.I0(GND_net), .I1(n8168[13]), .I2(n1105_adj_4166), 
            .I3(n29624), .O(n8146[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_16 (.CI(n29624), .I0(n8168[13]), .I1(n1105_adj_4166), 
            .CO(n29625));
    SB_LUT4 add_3752_15_lut (.I0(GND_net), .I1(n8168[12]), .I2(n1032_adj_4167), 
            .I3(n29623), .O(n8146[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_15 (.CI(n29623), .I0(n8168[12]), .I1(n1032_adj_4167), 
            .CO(n29624));
    SB_LUT4 add_3752_14_lut (.I0(GND_net), .I1(n8168[11]), .I2(n959_adj_4168), 
            .I3(n29622), .O(n8146[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_14 (.CI(n29622), .I0(n8168[11]), .I1(n959_adj_4168), 
            .CO(n29623));
    SB_LUT4 add_3728_19_lut (.I0(GND_net), .I1(n7826[16]), .I2(GND_net), 
            .I3(n29321), .O(n7802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_13_lut (.I0(GND_net), .I1(n8168[10]), .I2(n886_adj_4169), 
            .I3(n29621), .O(n8146[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_13 (.CI(n29621), .I0(n8168[10]), .I1(n886_adj_4169), 
            .CO(n29622));
    SB_LUT4 add_3752_12_lut (.I0(GND_net), .I1(n8168[9]), .I2(n813_adj_4170), 
            .I3(n29620), .O(n8146[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_12 (.CI(n29620), .I0(n8168[9]), .I1(n813_adj_4170), 
            .CO(n29621));
    SB_LUT4 i2_3_lut_4_lut_adj_979 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8092[0]), .I3(n27525), .O(n8087[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_979.LUT_INIT = 16'h8778;
    SB_LUT4 add_3752_11_lut (.I0(GND_net), .I1(n8168[8]), .I2(n740_adj_4171), 
            .I3(n29619), .O(n8146[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_11 (.CI(n29619), .I0(n8168[8]), .I1(n740_adj_4171), 
            .CO(n29620));
    SB_CARRY add_3728_19 (.CI(n29321), .I0(n7826[16]), .I1(GND_net), .CO(n29322));
    SB_LUT4 add_3752_10_lut (.I0(GND_net), .I1(n8168[7]), .I2(n667_adj_4172), 
            .I3(n29618), .O(n8146[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_10 (.CI(n29618), .I0(n8168[7]), .I1(n667_adj_4172), 
            .CO(n29619));
    SB_LUT4 add_3752_9_lut (.I0(GND_net), .I1(n8168[6]), .I2(n594_adj_4173), 
            .I3(n29617), .O(n8146[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_9 (.CI(n29617), .I0(n8168[6]), .I1(n594_adj_4173), 
            .CO(n29618));
    SB_LUT4 add_3752_8_lut (.I0(GND_net), .I1(n8168[5]), .I2(n521_adj_4174), 
            .I3(n29616), .O(n8146[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_8 (.CI(n29616), .I0(n8168[5]), .I1(n521_adj_4174), 
            .CO(n29617));
    SB_LUT4 add_3728_18_lut (.I0(GND_net), .I1(n7826[15]), .I2(GND_net), 
            .I3(n29320), .O(n7802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3752_7_lut (.I0(GND_net), .I1(n8168[4]), .I2(n448_adj_4175), 
            .I3(n29615), .O(n8146[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_7 (.CI(n29615), .I0(n8168[4]), .I1(n448_adj_4175), 
            .CO(n29616));
    SB_LUT4 add_3752_6_lut (.I0(GND_net), .I1(n8168[3]), .I2(n375_adj_4176), 
            .I3(n29614), .O(n8146[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_6 (.CI(n29614), .I0(n8168[3]), .I1(n375_adj_4176), 
            .CO(n29615));
    SB_LUT4 add_3752_5_lut (.I0(GND_net), .I1(n8168[2]), .I2(n302_adj_4177), 
            .I3(n29613), .O(n8146[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_5 (.CI(n29613), .I0(n8168[2]), .I1(n302_adj_4177), 
            .CO(n29614));
    SB_LUT4 add_3752_4_lut (.I0(GND_net), .I1(n8168[1]), .I2(n229_adj_4178), 
            .I3(n29612), .O(n8146[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_4 (.CI(n29612), .I0(n8168[1]), .I1(n229_adj_4178), 
            .CO(n29613));
    SB_LUT4 add_3752_3_lut (.I0(GND_net), .I1(n8168[0]), .I2(n156_adj_4179), 
            .I3(n29611), .O(n8146[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_3 (.CI(n29611), .I0(n8168[0]), .I1(n156_adj_4179), 
            .CO(n29612));
    SB_LUT4 add_3752_2_lut (.I0(GND_net), .I1(n14_adj_4180), .I2(n83_adj_4181), 
            .I3(GND_net), .O(n8146[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3752_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3752_2 (.CI(GND_net), .I0(n14_adj_4180), .I1(n83_adj_4181), 
            .CO(n29611));
    SB_LUT4 add_3751_22_lut (.I0(GND_net), .I1(n8146[19]), .I2(GND_net), 
            .I3(n29610), .O(n8123[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_21_lut (.I0(GND_net), .I1(n8146[18]), .I2(GND_net), 
            .I3(n29609), .O(n8123[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22858_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n27525));   // verilog/motorControl.v(42[17:23])
    defparam i22858_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_3751_21 (.CI(n29609), .I0(n8146[18]), .I1(GND_net), .CO(n29610));
    SB_LUT4 add_3751_20_lut (.I0(GND_net), .I1(n8146[17]), .I2(GND_net), 
            .I3(n29608), .O(n8123[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_20 (.CI(n29608), .I0(n8146[17]), .I1(GND_net), .CO(n29609));
    SB_LUT4 add_3751_19_lut (.I0(GND_net), .I1(n8146[16]), .I2(GND_net), 
            .I3(n29607), .O(n8123[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_19 (.CI(n29607), .I0(n8146[16]), .I1(GND_net), .CO(n29608));
    SB_LUT4 add_3751_18_lut (.I0(GND_net), .I1(n8146[15]), .I2(GND_net), 
            .I3(n29606), .O(n8123[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_18 (.CI(n29320), .I0(n7826[15]), .I1(GND_net), .CO(n29321));
    SB_LUT4 i22856_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8087[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22856_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_3751_18 (.CI(n29606), .I0(n8146[15]), .I1(GND_net), .CO(n29607));
    SB_LUT4 add_3751_17_lut (.I0(GND_net), .I1(n8146[14]), .I2(GND_net), 
            .I3(n29605), .O(n8123[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_17 (.CI(n29605), .I0(n8146[14]), .I1(GND_net), .CO(n29606));
    SB_LUT4 add_3751_16_lut (.I0(GND_net), .I1(n8146[13]), .I2(n1102_adj_4182), 
            .I3(n29604), .O(n8123[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_16 (.CI(n29604), .I0(n8146[13]), .I1(n1102_adj_4182), 
            .CO(n29605));
    SB_LUT4 add_3751_15_lut (.I0(GND_net), .I1(n8146[12]), .I2(n1029_adj_4183), 
            .I3(n29603), .O(n8123[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_15 (.CI(n29603), .I0(n8146[12]), .I1(n1029_adj_4183), 
            .CO(n29604));
    SB_LUT4 add_3751_14_lut (.I0(GND_net), .I1(n8146[11]), .I2(n956_adj_4184), 
            .I3(n29602), .O(n8123[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_14 (.CI(n29602), .I0(n8146[11]), .I1(n956_adj_4184), 
            .CO(n29603));
    SB_LUT4 add_3751_13_lut (.I0(GND_net), .I1(n8146[10]), .I2(n883_adj_4185), 
            .I3(n29601), .O(n8123[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_13 (.CI(n29601), .I0(n8146[10]), .I1(n883_adj_4185), 
            .CO(n29602));
    SB_LUT4 add_3751_12_lut (.I0(GND_net), .I1(n8146[9]), .I2(n810_adj_4186), 
            .I3(n29600), .O(n8123[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_12 (.CI(n29600), .I0(n8146[9]), .I1(n810_adj_4186), 
            .CO(n29601));
    SB_LUT4 add_3751_11_lut (.I0(GND_net), .I1(n8146[8]), .I2(n737_adj_4187), 
            .I3(n29599), .O(n8123[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_11 (.CI(n29599), .I0(n8146[8]), .I1(n737_adj_4187), 
            .CO(n29600));
    SB_LUT4 add_3751_10_lut (.I0(GND_net), .I1(n8146[7]), .I2(n664_adj_4188), 
            .I3(n29598), .O(n8123[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_10 (.CI(n29598), .I0(n8146[7]), .I1(n664_adj_4188), 
            .CO(n29599));
    SB_LUT4 add_3751_9_lut (.I0(GND_net), .I1(n8146[6]), .I2(n591_adj_4189), 
            .I3(n29597), .O(n8123[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_9 (.CI(n29597), .I0(n8146[6]), .I1(n591_adj_4189), 
            .CO(n29598));
    SB_LUT4 add_3728_17_lut (.I0(GND_net), .I1(n7826[14]), .I2(GND_net), 
            .I3(n29319), .O(n7802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3751_8_lut (.I0(GND_net), .I1(n8146[5]), .I2(n518_adj_4190), 
            .I3(n29596), .O(n8123[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_17 (.CI(n29319), .I0(n7826[14]), .I1(GND_net), .CO(n29320));
    SB_CARRY add_3751_8 (.CI(n29596), .I0(n8146[5]), .I1(n518_adj_4190), 
            .CO(n29597));
    SB_LUT4 add_3751_7_lut (.I0(GND_net), .I1(n8146[4]), .I2(n445_adj_4191), 
            .I3(n29595), .O(n8123[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_7 (.CI(n29595), .I0(n8146[4]), .I1(n445_adj_4191), 
            .CO(n29596));
    SB_LUT4 add_3751_6_lut (.I0(GND_net), .I1(n8146[3]), .I2(n372_adj_4192), 
            .I3(n29594), .O(n8123[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_6 (.CI(n29594), .I0(n8146[3]), .I1(n372_adj_4192), 
            .CO(n29595));
    SB_LUT4 add_3751_5_lut (.I0(GND_net), .I1(n8146[2]), .I2(n299_adj_4193), 
            .I3(n29593), .O(n8123[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_5 (.CI(n29593), .I0(n8146[2]), .I1(n299_adj_4193), 
            .CO(n29594));
    SB_LUT4 add_3751_4_lut (.I0(GND_net), .I1(n8146[1]), .I2(n226_adj_4194), 
            .I3(n29592), .O(n8123[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_4 (.CI(n29592), .I0(n8146[1]), .I1(n226_adj_4194), 
            .CO(n29593));
    SB_LUT4 add_3751_3_lut (.I0(GND_net), .I1(n8146[0]), .I2(n153_adj_4195), 
            .I3(n29591), .O(n8123[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_3 (.CI(n29591), .I0(n8146[0]), .I1(n153_adj_4195), 
            .CO(n29592));
    SB_LUT4 add_3751_2_lut (.I0(GND_net), .I1(n11_adj_4196), .I2(n80_adj_4197), 
            .I3(GND_net), .O(n8123[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3751_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3751_2 (.CI(GND_net), .I0(n11_adj_4196), .I1(n80_adj_4197), 
            .CO(n29591));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n8099[21]), 
            .I2(GND_net), .I3(n29590), .O(n40206)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8099[20]), .I2(GND_net), 
            .I3(n29589), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n29589), .I0(n8099[20]), .I1(GND_net), 
            .CO(n29590));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8099[19]), .I2(GND_net), 
            .I3(n29588), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n29588), .I0(n8099[19]), .I1(GND_net), 
            .CO(n29589));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8099[18]), .I2(GND_net), 
            .I3(n29587), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29587), .I0(n8099[18]), .I1(GND_net), 
            .CO(n29588));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8099[17]), .I2(GND_net), 
            .I3(n29586), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n29586), .I0(n8099[17]), .I1(GND_net), 
            .CO(n29587));
    SB_LUT4 add_3728_16_lut (.I0(GND_net), .I1(n7826[13]), .I2(n1099), 
            .I3(n29318), .O(n7802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8099[16]), .I2(GND_net), 
            .I3(n29585), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n29585), .I0(n8099[16]), .I1(GND_net), 
            .CO(n29586));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8099[15]), .I2(GND_net), 
            .I3(n29584), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n29584), .I0(n8099[15]), .I1(GND_net), 
            .CO(n29585));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8099[14]), .I2(GND_net), 
            .I3(n29583), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n29583), .I0(n8099[14]), .I1(GND_net), 
            .CO(n29584));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8099[13]), .I2(n1096_adj_4198), 
            .I3(n29582), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29582), .I0(n8099[13]), .I1(n1096_adj_4198), 
            .CO(n29583));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_4253[23]), .I3(n28083), .O(\PID_CONTROLLER.err_23__N_3638 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8099[12]), .I2(n1023_adj_4201), 
            .I3(n29581), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n29581), .I0(n8099[12]), .I1(n1023_adj_4201), 
            .CO(n29582));
    SB_CARRY add_3728_16 (.CI(n29318), .I0(n7826[13]), .I1(n1099), .CO(n29319));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8099[11]), .I2(n950_adj_4202), 
            .I3(n29580), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29580), .I0(n8099[11]), .I1(n950_adj_4202), 
            .CO(n29581));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_4253[22]), .I3(n28082), .O(\PID_CONTROLLER.err_23__N_3638 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8099[10]), .I2(n877_adj_4204), 
            .I3(n29579), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n29579), .I0(n8099[10]), .I1(n877_adj_4204), 
            .CO(n29580));
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3728_15_lut (.I0(GND_net), .I1(n7826[12]), .I2(n1026), 
            .I3(n29317), .O(n7802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8099[9]), .I2(n804_adj_4207), 
            .I3(n29578), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_15 (.CI(n29317), .I0(n7826[12]), .I1(n1026), .CO(n29318));
    SB_CARRY state_23__I_0_add_2_24 (.CI(n28082), .I0(motor_state[22]), 
            .I1(n1_adj_4253[22]), .CO(n28083));
    SB_CARRY mult_11_add_1225_12 (.CI(n29578), .I0(n8099[9]), .I1(n804_adj_4207), 
            .CO(n29579));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8099[8]), .I2(n731_adj_4208), 
            .I3(n29577), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_4253[21]), .I3(n28081), .O(\PID_CONTROLLER.err_23__N_3638 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n28081), .I0(motor_state[21]), 
            .I1(n1_adj_4253[21]), .CO(n28082));
    SB_CARRY mult_11_add_1225_11 (.CI(n29577), .I0(n8099[8]), .I1(n731_adj_4208), 
            .CO(n29578));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_4253[20]), .I3(n28080), .O(\PID_CONTROLLER.err_23__N_3638 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8099[7]), .I2(n658_adj_4211), 
            .I3(n29576), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n29576), .I0(n8099[7]), .I1(n658_adj_4211), 
            .CO(n29577));
    SB_CARRY state_23__I_0_add_2_22 (.CI(n28080), .I0(motor_state[20]), 
            .I1(n1_adj_4253[20]), .CO(n28081));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8099[6]), .I2(n585_adj_4213), 
            .I3(n29575), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_4253[19]), .I3(n28079), .O(\PID_CONTROLLER.err_23__N_3638 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n29575), .I0(n8099[6]), .I1(n585_adj_4213), 
            .CO(n29576));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8099[5]), .I2(n512_adj_4215), 
            .I3(n29574), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n29574), .I0(n8099[5]), .I1(n512_adj_4215), 
            .CO(n29575));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8099[4]), .I2(n439_adj_4216), 
            .I3(n29573), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n29573), .I0(n8099[4]), .I1(n439_adj_4216), 
            .CO(n29574));
    SB_LUT4 i22807_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4217), .I3(n8081[1]), .O(n6_adj_3967));   // verilog/motorControl.v(42[17:23])
    defparam i22807_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8099[3]), .I2(n366_adj_4219), 
            .I3(n29572), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n28079), .I0(motor_state[19]), 
            .I1(n1_adj_4253[19]), .CO(n28080));
    SB_CARRY mult_11_add_1225_6 (.CI(n29572), .I0(n8099[3]), .I1(n366_adj_4219), 
            .CO(n29573));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_4253[18]), .I3(n28078), .O(\PID_CONTROLLER.err_23__N_3638 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8099[2]), .I2(n293_adj_4221), 
            .I3(n29571), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n28078), .I0(motor_state[18]), 
            .I1(n1_adj_4253[18]), .CO(n28079));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_4253[17]), .I3(n28077), .O(\PID_CONTROLLER.err_23__N_3638 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n28077), .I0(motor_state[17]), 
            .I1(n1_adj_4253[17]), .CO(n28078));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_4253[16]), .I3(n28076), .O(\PID_CONTROLLER.err_23__N_3638 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n28076), .I0(motor_state[16]), 
            .I1(n1_adj_4253[16]), .CO(n28077));
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_4253[15]), .I3(n28075), .O(\PID_CONTROLLER.err_23__N_3638 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n28075), .I0(motor_state[15]), 
            .I1(n1_adj_4253[15]), .CO(n28076));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_4253[14]), .I3(n28074), .O(\PID_CONTROLLER.err_23__N_3638 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n29571), .I0(n8099[2]), .I1(n293_adj_4221), 
            .CO(n29572));
    SB_CARRY state_23__I_0_add_2_16 (.CI(n28074), .I0(motor_state[14]), 
            .I1(n1_adj_4253[14]), .CO(n28075));
    SB_LUT4 add_3728_14_lut (.I0(GND_net), .I1(n7826[11]), .I2(n953), 
            .I3(n29316), .O(n7802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_4253[13]), .I3(n28073), .O(\PID_CONTROLLER.err_23__N_3638 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n28073), .I0(motor_state[13]), 
            .I1(n1_adj_4253[13]), .CO(n28074));
    SB_CARRY add_3728_14 (.CI(n29316), .I0(n7826[11]), .I1(n953), .CO(n29317));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8099[1]), .I2(n220_adj_4227), 
            .I3(n29570), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n29570), .I0(n8099[1]), .I1(n220_adj_4227), 
            .CO(n29571));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8099[0]), .I2(n147_adj_4228), 
            .I3(n29569), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_4253[12]), .I3(n28072), .O(\PID_CONTROLLER.err_23__N_3638 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29569), .I0(n8099[0]), .I1(n147_adj_4228), 
            .CO(n29570));
    SB_CARRY state_23__I_0_add_2_14 (.CI(n28072), .I0(motor_state[12]), 
            .I1(n1_adj_4253[12]), .CO(n28073));
    SB_LUT4 add_3728_13_lut (.I0(GND_net), .I1(n7826[10]), .I2(n880), 
            .I3(n29315), .O(n7802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_980 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8081[1]), .I3(n4_adj_4217), .O(n8074[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_980.LUT_INIT = 16'h8778;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_4253[11]), .I3(n28071), .O(\PID_CONTROLLER.err_23__N_3638 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_13 (.CI(n29315), .I0(n7826[10]), .I1(n880), .CO(n29316));
    SB_CARRY state_23__I_0_add_2_13 (.CI(n28071), .I0(motor_state[11]), 
            .I1(n1_adj_4253[11]), .CO(n28072));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4231), .I2(n74_adj_4232), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4231), .I1(n74_adj_4232), 
            .CO(n29569));
    SB_LUT4 add_3750_23_lut (.I0(GND_net), .I1(n8123[20]), .I2(GND_net), 
            .I3(n29568), .O(n8099[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_4253[10]), .I3(n28070), .O(\PID_CONTROLLER.err_23__N_3638 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3750_22_lut (.I0(GND_net), .I1(n8123[19]), .I2(GND_net), 
            .I3(n29567), .O(n8099[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_22 (.CI(n29567), .I0(n8123[19]), .I1(GND_net), .CO(n29568));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n28070), .I0(motor_state[10]), 
            .I1(n1_adj_4253[10]), .CO(n28071));
    SB_LUT4 add_3750_21_lut (.I0(GND_net), .I1(n8123[18]), .I2(GND_net), 
            .I3(n29566), .O(n8099[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_21 (.CI(n29566), .I0(n8123[18]), .I1(GND_net), .CO(n29567));
    SB_LUT4 add_3750_20_lut (.I0(GND_net), .I1(n8123[17]), .I2(GND_net), 
            .I3(n29565), .O(n8099[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_12_lut (.I0(GND_net), .I1(n7826[9]), .I2(n807), .I3(n29314), 
            .O(n7802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_12 (.CI(n29314), .I0(n7826[9]), .I1(n807), .CO(n29315));
    SB_CARRY add_3750_20 (.CI(n29565), .I0(n8123[17]), .I1(GND_net), .CO(n29566));
    SB_LUT4 add_3728_11_lut (.I0(GND_net), .I1(n7826[8]), .I2(n734), .I3(n29313), 
            .O(n7802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_11 (.CI(n29313), .I0(n7826[8]), .I1(n734), .CO(n29314));
    SB_LUT4 add_3750_19_lut (.I0(GND_net), .I1(n8123[16]), .I2(GND_net), 
            .I3(n29564), .O(n8099[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_19 (.CI(n29564), .I0(n8123[16]), .I1(GND_net), .CO(n29565));
    SB_LUT4 add_3750_18_lut (.I0(GND_net), .I1(n8123[15]), .I2(GND_net), 
            .I3(n29563), .O(n8099[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_18 (.CI(n29563), .I0(n8123[15]), .I1(GND_net), .CO(n29564));
    SB_LUT4 add_3750_17_lut (.I0(GND_net), .I1(n8123[14]), .I2(GND_net), 
            .I3(n29562), .O(n8099[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_17 (.CI(n29562), .I0(n8123[14]), .I1(GND_net), .CO(n29563));
    SB_LUT4 add_3750_16_lut (.I0(GND_net), .I1(n8123[13]), .I2(n1099_adj_4234), 
            .I3(n29561), .O(n8099[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_16 (.CI(n29561), .I0(n8123[13]), .I1(n1099_adj_4234), 
            .CO(n29562));
    SB_LUT4 add_3750_15_lut (.I0(GND_net), .I1(n8123[12]), .I2(n1026_adj_4235), 
            .I3(n29560), .O(n8099[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_15 (.CI(n29560), .I0(n8123[12]), .I1(n1026_adj_4235), 
            .CO(n29561));
    SB_LUT4 add_3750_14_lut (.I0(GND_net), .I1(n8123[11]), .I2(n953_adj_4236), 
            .I3(n29559), .O(n8099[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_14 (.CI(n29559), .I0(n8123[11]), .I1(n953_adj_4236), 
            .CO(n29560));
    SB_LUT4 add_3750_13_lut (.I0(GND_net), .I1(n8123[10]), .I2(n880_adj_4237), 
            .I3(n29558), .O(n8099[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_13 (.CI(n29558), .I0(n8123[10]), .I1(n880_adj_4237), 
            .CO(n29559));
    SB_LUT4 add_3750_12_lut (.I0(GND_net), .I1(n8123[9]), .I2(n807_adj_4238), 
            .I3(n29557), .O(n8099[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_12 (.CI(n29557), .I0(n8123[9]), .I1(n807_adj_4238), 
            .CO(n29558));
    SB_LUT4 add_3750_11_lut (.I0(GND_net), .I1(n8123[8]), .I2(n734_adj_4239), 
            .I3(n29556), .O(n8099[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_11 (.CI(n29556), .I0(n8123[8]), .I1(n734_adj_4239), 
            .CO(n29557));
    SB_LUT4 add_3750_10_lut (.I0(GND_net), .I1(n8123[7]), .I2(n661), .I3(n29555), 
            .O(n8099[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_10 (.CI(n29555), .I0(n8123[7]), .I1(n661), .CO(n29556));
    SB_LUT4 add_3750_9_lut (.I0(GND_net), .I1(n8123[6]), .I2(n588_adj_4240), 
            .I3(n29554), .O(n8099[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_9 (.CI(n29554), .I0(n8123[6]), .I1(n588_adj_4240), 
            .CO(n29555));
    SB_LUT4 add_3728_10_lut (.I0(GND_net), .I1(n7826[7]), .I2(n661_adj_4241), 
            .I3(n29312), .O(n7802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_4253[9]), .I3(n28069), .O(\PID_CONTROLLER.err_23__N_3638 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n28069), .I0(motor_state[9]), .I1(n1_adj_4253[9]), 
            .CO(n28070));
    SB_LUT4 i2_3_lut_4_lut_adj_981 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8081[0]), .I3(n27448), .O(n8074[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_981.LUT_INIT = 16'h8778;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_4253[8]), .I3(n28068), .O(\PID_CONTROLLER.err_23__N_3638 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n28068), .I0(motor_state[8]), .I1(n1_adj_4253[8]), 
            .CO(n28069));
    SB_LUT4 add_3750_8_lut (.I0(GND_net), .I1(n8123[5]), .I2(n515_adj_4244), 
            .I3(n29553), .O(n8099[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_4253[7]), .I3(n28067), .O(\PID_CONTROLLER.err_23__N_3638 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_10 (.CI(n29312), .I0(n7826[7]), .I1(n661_adj_4241), 
            .CO(n29313));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n28067), .I0(motor_state[7]), .I1(n1_adj_4253[7]), 
            .CO(n28068));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_4253[6]), .I3(n28066), .O(\PID_CONTROLLER.err_23__N_3638 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_8 (.CI(n29553), .I0(n8123[5]), .I1(n515_adj_4244), 
            .CO(n29554));
    SB_LUT4 add_3750_7_lut (.I0(GND_net), .I1(n8123[4]), .I2(n442_adj_4143), 
            .I3(n29552), .O(n8099[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_7 (.CI(n29552), .I0(n8123[4]), .I1(n442_adj_4143), 
            .CO(n29553));
    SB_LUT4 add_3750_6_lut (.I0(GND_net), .I1(n8123[3]), .I2(n369_adj_4136), 
            .I3(n29551), .O(n8099[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_6 (.CI(n29551), .I0(n8123[3]), .I1(n369_adj_4136), 
            .CO(n29552));
    SB_LUT4 add_3750_5_lut (.I0(GND_net), .I1(n8123[2]), .I2(n296_adj_4131), 
            .I3(n29550), .O(n8099[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_5 (.CI(n29550), .I0(n8123[2]), .I1(n296_adj_4131), 
            .CO(n29551));
    SB_CARRY state_23__I_0_add_2_8 (.CI(n28066), .I0(motor_state[6]), .I1(n1_adj_4253[6]), 
            .CO(n28067));
    SB_LUT4 add_3750_4_lut (.I0(GND_net), .I1(n8123[1]), .I2(n223_adj_4130), 
            .I3(n29549), .O(n8099[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_4 (.CI(n29549), .I0(n8123[1]), .I1(n223_adj_4130), 
            .CO(n29550));
    SB_LUT4 add_3750_3_lut (.I0(GND_net), .I1(n8123[0]), .I2(n150_adj_4127), 
            .I3(n29548), .O(n8099[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_4253[5]), .I3(n28065), .O(\PID_CONTROLLER.err_23__N_3638 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_3 (.CI(n29548), .I0(n8123[0]), .I1(n150_adj_4127), 
            .CO(n29549));
    SB_LUT4 add_3750_2_lut (.I0(GND_net), .I1(n8_adj_4050), .I2(n77_adj_4049), 
            .I3(GND_net), .O(n8099[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3750_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3750_2 (.CI(GND_net), .I0(n8_adj_4050), .I1(n77_adj_4049), 
            .CO(n29548));
    SB_CARRY state_23__I_0_add_2_7 (.CI(n28065), .I0(motor_state[5]), .I1(n1_adj_4253[5]), 
            .CO(n28066));
    SB_LUT4 add_3744_7_lut (.I0(GND_net), .I1(n36490), .I2(n490), .I3(n29547), 
            .O(n8066[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_4253[4]), .I3(n28064), .O(\PID_CONTROLLER.err_23__N_3638 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n28064), .I0(motor_state[4]), .I1(n1_adj_4253[4]), 
            .CO(n28065));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_4253[3]), .I3(n28063), .O(\PID_CONTROLLER.err_23__N_3638 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n28063), .I0(motor_state[3]), .I1(n1_adj_4253[3]), 
            .CO(n28064));
    SB_LUT4 add_3744_6_lut (.I0(GND_net), .I1(n8074[3]), .I2(n417), .I3(n29546), 
            .O(n8066[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_6 (.CI(n29546), .I0(n8074[3]), .I1(n417), .CO(n29547));
    SB_LUT4 add_3744_5_lut (.I0(GND_net), .I1(n8074[2]), .I2(n344), .I3(n29545), 
            .O(n8066[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_9_lut (.I0(GND_net), .I1(n7826[6]), .I2(n588), .I3(n29311), 
            .O(n7802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_5 (.CI(n29545), .I0(n8074[2]), .I1(n344), .CO(n29546));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_4253[2]), .I3(n28062), .O(\PID_CONTROLLER.err_23__N_3638 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3744_4_lut (.I0(GND_net), .I1(n8074[1]), .I2(n271_adj_3965), 
            .I3(n29544), .O(n8066[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_4 (.CI(n29544), .I0(n8074[1]), .I1(n271_adj_3965), 
            .CO(n29545));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n28062), .I0(motor_state[2]), .I1(n1_adj_4253[2]), 
            .CO(n28063));
    SB_LUT4 add_3744_3_lut (.I0(GND_net), .I1(n8074[0]), .I2(n198), .I3(n29543), 
            .O(n8066[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_3 (.CI(n29543), .I0(n8074[0]), .I1(n198), .CO(n29544));
    SB_LUT4 add_3744_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_3964), 
            .I3(GND_net), .O(n8066[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3744_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_4253[1]), .I3(n28061), .O(\PID_CONTROLLER.err_23__N_3638 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3744_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_3964), .CO(n29543));
    SB_CARRY add_3728_9 (.CI(n29311), .I0(n7826[6]), .I1(n588), .CO(n29312));
    SB_LUT4 add_3743_8_lut (.I0(GND_net), .I1(n8066[5]), .I2(n560), .I3(n29542), 
            .O(n8057[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22799_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n27448), .I3(n8081[0]), .O(n4_adj_4217));   // verilog/motorControl.v(42[17:23])
    defparam i22799_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_3743_7_lut (.I0(GND_net), .I1(n8066[4]), .I2(n487), .I3(n29541), 
            .O(n8057[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_7 (.CI(n29541), .I0(n8066[4]), .I1(n487), .CO(n29542));
    SB_LUT4 add_3743_6_lut (.I0(GND_net), .I1(n8066[3]), .I2(n414), .I3(n29540), 
            .O(n8057[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_6 (.CI(n29540), .I0(n8066[3]), .I1(n414), .CO(n29541));
    SB_LUT4 add_3743_5_lut (.I0(GND_net), .I1(n8066[2]), .I2(n341), .I3(n29539), 
            .O(n8057[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n28061), .I0(motor_state[1]), .I1(n1_adj_4253[1]), 
            .CO(n28062));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_4253[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3638 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_4253[0]), 
            .CO(n28061));
    SB_LUT4 add_3728_8_lut (.I0(GND_net), .I1(n7826[5]), .I2(n515), .I3(n29310), 
            .O(n7802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3743_5 (.CI(n29539), .I0(n8066[2]), .I1(n341), .CO(n29540));
    SB_CARRY add_3728_8 (.CI(n29310), .I0(n7826[5]), .I1(n515), .CO(n29311));
    SB_LUT4 add_3728_7_lut (.I0(GND_net), .I1(n7826[4]), .I2(n442), .I3(n29309), 
            .O(n7802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_7 (.CI(n29309), .I0(n7826[4]), .I1(n442), .CO(n29310));
    SB_LUT4 add_3728_6_lut (.I0(GND_net), .I1(n7826[3]), .I2(n369), .I3(n29308), 
            .O(n7802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_6 (.CI(n29308), .I0(n7826[3]), .I1(n369), .CO(n29309));
    SB_LUT4 add_3743_4_lut (.I0(GND_net), .I1(n8066[1]), .I2(n268_adj_3961), 
            .I3(n29538), .O(n8057[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_5_lut (.I0(GND_net), .I1(n7826[2]), .I2(n296), .I3(n29307), 
            .O(n7802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_5 (.CI(n29307), .I0(n7826[2]), .I1(n296), .CO(n29308));
    SB_LUT4 add_3728_4_lut (.I0(GND_net), .I1(n7826[1]), .I2(n223), .I3(n29306), 
            .O(n7802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_4 (.CI(n29306), .I0(n7826[1]), .I1(n223), .CO(n29307));
    SB_LUT4 i22786_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8074[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22786_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3728_3_lut (.I0(GND_net), .I1(n7826[0]), .I2(n150), .I3(n29305), 
            .O(n7802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_4 (.CI(n29538), .I0(n8066[1]), .I1(n268_adj_3961), 
            .CO(n29539));
    SB_CARRY add_3728_3 (.CI(n29305), .I0(n7826[0]), .I1(n150), .CO(n29306));
    SB_LUT4 add_3728_2_lut (.I0(GND_net), .I1(n8_adj_3960), .I2(n77), 
            .I3(GND_net), .O(n7802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_2 (.CI(GND_net), .I0(n8_adj_3960), .I1(n77), .CO(n29305));
    SB_LUT4 add_3743_3_lut (.I0(GND_net), .I1(n8066[0]), .I2(n195), .I3(n29537), 
            .O(n8057[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_3 (.CI(n29537), .I0(n8066[0]), .I1(n195), .CO(n29538));
    SB_LUT4 add_3743_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_3959), 
            .I3(GND_net), .O(n8057[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3743_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3743_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_3959), .CO(n29537));
    SB_LUT4 add_3742_9_lut (.I0(GND_net), .I1(n8057[6]), .I2(n630), .I3(n29536), 
            .O(n8047[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3742_8_lut (.I0(GND_net), .I1(n8057[5]), .I2(n557), .I3(n29535), 
            .O(n8047[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_8 (.CI(n29535), .I0(n8057[5]), .I1(n557), .CO(n29536));
    SB_LUT4 add_3742_7_lut (.I0(GND_net), .I1(n8057[4]), .I2(n484), .I3(n29534), 
            .O(n8047[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_7 (.CI(n29534), .I0(n8057[4]), .I1(n484), .CO(n29535));
    SB_LUT4 add_3742_6_lut (.I0(GND_net), .I1(n8057[3]), .I2(n411), .I3(n29533), 
            .O(n8047[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_6 (.CI(n29533), .I0(n8057[3]), .I1(n411), .CO(n29534));
    SB_LUT4 add_3742_5_lut (.I0(GND_net), .I1(n8057[2]), .I2(n338), .I3(n29532), 
            .O(n8047[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_5 (.CI(n29532), .I0(n8057[2]), .I1(n338), .CO(n29533));
    SB_LUT4 add_3742_4_lut (.I0(GND_net), .I1(n8057[1]), .I2(n265_adj_3957), 
            .I3(n29531), .O(n8047[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_4 (.CI(n29531), .I0(n8057[1]), .I1(n265_adj_3957), 
            .CO(n29532));
    SB_LUT4 add_3742_3_lut (.I0(GND_net), .I1(n8057[0]), .I2(n192), .I3(n29530), 
            .O(n8047[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_3 (.CI(n29530), .I0(n8057[0]), .I1(n192), .CO(n29531));
    SB_LUT4 add_3742_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_3956), 
            .I3(GND_net), .O(n8047[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3742_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3742_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_3956), .CO(n29530));
    SB_LUT4 add_3741_10_lut (.I0(GND_net), .I1(n8047[7]), .I2(n700), .I3(n29529), 
            .O(n8036[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3741_9_lut (.I0(GND_net), .I1(n8047[6]), .I2(n627), .I3(n29528), 
            .O(n8036[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_9 (.CI(n29528), .I0(n8047[6]), .I1(n627), .CO(n29529));
    SB_LUT4 add_3741_8_lut (.I0(GND_net), .I1(n8047[5]), .I2(n554), .I3(n29527), 
            .O(n8036[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_8 (.CI(n29527), .I0(n8047[5]), .I1(n554), .CO(n29528));
    SB_LUT4 add_3741_7_lut (.I0(GND_net), .I1(n8047[4]), .I2(n481), .I3(n29526), 
            .O(n8036[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_7 (.CI(n29526), .I0(n8047[4]), .I1(n481), .CO(n29527));
    SB_LUT4 add_3741_6_lut (.I0(GND_net), .I1(n8047[3]), .I2(n408), .I3(n29525), 
            .O(n8036[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_6 (.CI(n29525), .I0(n8047[3]), .I1(n408), .CO(n29526));
    SB_LUT4 add_3741_5_lut (.I0(GND_net), .I1(n8047[2]), .I2(n335), .I3(n29524), 
            .O(n8036[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_5 (.CI(n29524), .I0(n8047[2]), .I1(n335), .CO(n29525));
    SB_LUT4 add_3741_4_lut (.I0(GND_net), .I1(n8047[1]), .I2(n262_adj_3955), 
            .I3(n29523), .O(n8036[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_4 (.CI(n29523), .I0(n8047[1]), .I1(n262_adj_3955), 
            .CO(n29524));
    SB_LUT4 add_3741_3_lut (.I0(GND_net), .I1(n8047[0]), .I2(n189), .I3(n29522), 
            .O(n8036[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_3 (.CI(n29522), .I0(n8047[0]), .I1(n189), .CO(n29523));
    SB_LUT4 add_3741_2_lut (.I0(GND_net), .I1(n47_adj_3954), .I2(n116_adj_3953), 
            .I3(GND_net), .O(n8036[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3741_2 (.CI(GND_net), .I0(n47_adj_3954), .I1(n116_adj_3953), 
            .CO(n29522));
    SB_LUT4 add_3740_11_lut (.I0(GND_net), .I1(n8036[8]), .I2(n770), .I3(n29521), 
            .O(n8024[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3740_10_lut (.I0(GND_net), .I1(n8036[7]), .I2(n697), .I3(n29520), 
            .O(n8024[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_10 (.CI(n29520), .I0(n8036[7]), .I1(n697), .CO(n29521));
    SB_LUT4 i22788_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n27448));   // verilog/motorControl.v(42[17:23])
    defparam i22788_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3740_9_lut (.I0(GND_net), .I1(n8036[6]), .I2(n624), .I3(n29519), 
            .O(n8024[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4244));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3740_9 (.CI(n29519), .I0(n8036[6]), .I1(n624), .CO(n29520));
    SB_LUT4 add_3740_8_lut (.I0(GND_net), .I1(n8036[5]), .I2(n551), .I3(n29518), 
            .O(n8024[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_8 (.CI(n29518), .I0(n8036[5]), .I1(n551), .CO(n29519));
    SB_LUT4 add_3740_7_lut (.I0(GND_net), .I1(n8036[4]), .I2(n478), .I3(n29517), 
            .O(n8024[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_7 (.CI(n29517), .I0(n8036[4]), .I1(n478), .CO(n29518));
    SB_LUT4 add_3740_6_lut (.I0(GND_net), .I1(n8036[3]), .I2(n405), .I3(n29516), 
            .O(n8024[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_6 (.CI(n29516), .I0(n8036[3]), .I1(n405), .CO(n29517));
    SB_LUT4 add_3740_5_lut (.I0(GND_net), .I1(n8036[2]), .I2(n332), .I3(n29515), 
            .O(n8024[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_5 (.CI(n29515), .I0(n8036[2]), .I1(n332), .CO(n29516));
    SB_LUT4 add_3740_4_lut (.I0(GND_net), .I1(n8036[1]), .I2(n259_adj_3950), 
            .I3(n29514), .O(n8024[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_4 (.CI(n29514), .I0(n8036[1]), .I1(n259_adj_3950), 
            .CO(n29515));
    SB_LUT4 add_3740_3_lut (.I0(GND_net), .I1(n8036[0]), .I2(n186_adj_3948), 
            .I3(n29513), .O(n8024[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_3 (.CI(n29513), .I0(n8036[0]), .I1(n186_adj_3948), 
            .CO(n29514));
    SB_LUT4 add_3740_2_lut (.I0(GND_net), .I1(n44), .I2(n113_adj_3946), 
            .I3(GND_net), .O(n8024[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3740_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3740_2 (.CI(GND_net), .I0(n44), .I1(n113_adj_3946), .CO(n29513));
    SB_LUT4 add_3739_12_lut (.I0(GND_net), .I1(n8024[9]), .I2(n840), .I3(n29512), 
            .O(n8011[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3739_11_lut (.I0(GND_net), .I1(n8024[8]), .I2(n767), .I3(n29511), 
            .O(n8011[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_11 (.CI(n29511), .I0(n8024[8]), .I1(n767), .CO(n29512));
    SB_LUT4 add_3739_10_lut (.I0(GND_net), .I1(n8024[7]), .I2(n694), .I3(n29510), 
            .O(n8011[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_10 (.CI(n29510), .I0(n8024[7]), .I1(n694), .CO(n29511));
    SB_LUT4 add_3739_9_lut (.I0(GND_net), .I1(n8024[6]), .I2(n621), .I3(n29509), 
            .O(n8011[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_9 (.CI(n29509), .I0(n8024[6]), .I1(n621), .CO(n29510));
    SB_LUT4 add_3739_8_lut (.I0(GND_net), .I1(n8024[5]), .I2(n548), .I3(n29508), 
            .O(n8011[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_8 (.CI(n29508), .I0(n8024[5]), .I1(n548), .CO(n29509));
    SB_LUT4 add_3739_7_lut (.I0(GND_net), .I1(n8024[4]), .I2(n475), .I3(n29507), 
            .O(n8011[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_7 (.CI(n29507), .I0(n8024[4]), .I1(n475), .CO(n29508));
    SB_LUT4 add_3739_6_lut (.I0(GND_net), .I1(n8024[3]), .I2(n402), .I3(n29506), 
            .O(n8011[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_6 (.CI(n29506), .I0(n8024[3]), .I1(n402), .CO(n29507));
    SB_LUT4 add_3739_5_lut (.I0(GND_net), .I1(n8024[2]), .I2(n329), .I3(n29505), 
            .O(n8011[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_5 (.CI(n29505), .I0(n8024[2]), .I1(n329), .CO(n29506));
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3739_4_lut (.I0(GND_net), .I1(n8024[1]), .I2(n256_adj_3941), 
            .I3(n29504), .O(n8011[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_4 (.CI(n29504), .I0(n8024[1]), .I1(n256_adj_3941), 
            .CO(n29505));
    SB_LUT4 add_3739_3_lut (.I0(GND_net), .I1(n8024[0]), .I2(n183_adj_3939), 
            .I3(n29503), .O(n8011[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_3 (.CI(n29503), .I0(n8024[0]), .I1(n183_adj_3939), 
            .CO(n29504));
    SB_LUT4 add_3739_2_lut (.I0(GND_net), .I1(n41_adj_3938), .I2(n110_adj_3937), 
            .I3(GND_net), .O(n8011[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3739_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3739_2 (.CI(GND_net), .I0(n41_adj_3938), .I1(n110_adj_3937), 
            .CO(n29503));
    SB_LUT4 add_3738_13_lut (.I0(GND_net), .I1(n8011[10]), .I2(n910), 
            .I3(n29502), .O(n7997[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3738_12_lut (.I0(GND_net), .I1(n8011[9]), .I2(n837), .I3(n29501), 
            .O(n7997[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_12 (.CI(n29501), .I0(n8011[9]), .I1(n837), .CO(n29502));
    SB_LUT4 add_3738_11_lut (.I0(GND_net), .I1(n8011[8]), .I2(n764), .I3(n29500), 
            .O(n7997[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_11 (.CI(n29500), .I0(n8011[8]), .I1(n764), .CO(n29501));
    SB_LUT4 add_3738_10_lut (.I0(GND_net), .I1(n8011[7]), .I2(n691), .I3(n29499), 
            .O(n7997[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_10 (.CI(n29499), .I0(n8011[7]), .I1(n691), .CO(n29500));
    SB_LUT4 add_3738_9_lut (.I0(GND_net), .I1(n8011[6]), .I2(n618), .I3(n29498), 
            .O(n7997[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_9 (.CI(n29498), .I0(n8011[6]), .I1(n618), .CO(n29499));
    SB_LUT4 i22825_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n8081[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22825_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3738_8_lut (.I0(GND_net), .I1(n8011[5]), .I2(n545), .I3(n29497), 
            .O(n7997[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_8 (.CI(n29497), .I0(n8011[5]), .I1(n545), .CO(n29498));
    SB_LUT4 add_3738_7_lut (.I0(GND_net), .I1(n8011[4]), .I2(n472), .I3(n29496), 
            .O(n7997[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_7 (.CI(n29496), .I0(n8011[4]), .I1(n472), .CO(n29497));
    SB_LUT4 add_3738_6_lut (.I0(GND_net), .I1(n8011[3]), .I2(n399), .I3(n29495), 
            .O(n7997[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_6 (.CI(n29495), .I0(n8011[3]), .I1(n399), .CO(n29496));
    SB_LUT4 add_3738_5_lut (.I0(GND_net), .I1(n8011[2]), .I2(n326), .I3(n29494), 
            .O(n7997[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_5 (.CI(n29494), .I0(n8011[2]), .I1(n326), .CO(n29495));
    SB_LUT4 add_3738_4_lut (.I0(GND_net), .I1(n8011[1]), .I2(n253), .I3(n29493), 
            .O(n7997[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_4 (.CI(n29493), .I0(n8011[1]), .I1(n253), .CO(n29494));
    SB_LUT4 i22827_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n27491));   // verilog/motorControl.v(42[17:23])
    defparam i22827_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3738_3_lut (.I0(GND_net), .I1(n8011[0]), .I2(n180), .I3(n29492), 
            .O(n7997[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_3 (.CI(n29492), .I0(n8011[0]), .I1(n180), .CO(n29493));
    SB_LUT4 add_3738_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_3935), 
            .I3(GND_net), .O(n7997[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3738_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3738_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_3935), .CO(n29492));
    SB_LUT4 add_3737_14_lut (.I0(GND_net), .I1(n7997[11]), .I2(n980), 
            .I3(n29491), .O(n7982[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3737_13_lut (.I0(GND_net), .I1(n7997[10]), .I2(n907), 
            .I3(n29490), .O(n7982[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_13 (.CI(n29490), .I0(n7997[10]), .I1(n907), .CO(n29491));
    SB_LUT4 add_3737_12_lut (.I0(GND_net), .I1(n7997[9]), .I2(n834), .I3(n29489), 
            .O(n7982[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_12 (.CI(n29489), .I0(n7997[9]), .I1(n834), .CO(n29490));
    SB_LUT4 add_3737_11_lut (.I0(GND_net), .I1(n7997[8]), .I2(n761), .I3(n29488), 
            .O(n7982[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_11 (.CI(n29488), .I0(n7997[8]), .I1(n761), .CO(n29489));
    SB_LUT4 add_3737_10_lut (.I0(GND_net), .I1(n7997[7]), .I2(n688), .I3(n29487), 
            .O(n7982[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_10 (.CI(n29487), .I0(n7997[7]), .I1(n688), .CO(n29488));
    SB_LUT4 add_3737_9_lut (.I0(GND_net), .I1(n7997[6]), .I2(n615), .I3(n29486), 
            .O(n7982[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_9 (.CI(n29486), .I0(n7997[6]), .I1(n615), .CO(n29487));
    SB_LUT4 add_3737_8_lut (.I0(GND_net), .I1(n7997[5]), .I2(n542), .I3(n29485), 
            .O(n7982[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_8 (.CI(n29485), .I0(n7997[5]), .I1(n542), .CO(n29486));
    SB_LUT4 add_3737_7_lut (.I0(GND_net), .I1(n7997[4]), .I2(n469), .I3(n29484), 
            .O(n7982[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_7 (.CI(n29484), .I0(n7997[4]), .I1(n469), .CO(n29485));
    SB_LUT4 add_3737_6_lut (.I0(GND_net), .I1(n7997[3]), .I2(n396), .I3(n29483), 
            .O(n7982[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_6 (.CI(n29483), .I0(n7997[3]), .I1(n396), .CO(n29484));
    SB_LUT4 add_3737_5_lut (.I0(GND_net), .I1(n7997[2]), .I2(n323), .I3(n29482), 
            .O(n7982[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_5 (.CI(n29482), .I0(n7997[2]), .I1(n323), .CO(n29483));
    SB_LUT4 add_3737_4_lut (.I0(GND_net), .I1(n7997[1]), .I2(n250), .I3(n29481), 
            .O(n7982[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_4 (.CI(n29481), .I0(n7997[1]), .I1(n250), .CO(n29482));
    SB_LUT4 add_3737_3_lut (.I0(GND_net), .I1(n7997[0]), .I2(n177), .I3(n29480), 
            .O(n7982[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_3 (.CI(n29480), .I0(n7997[0]), .I1(n177), .CO(n29481));
    SB_LUT4 add_3737_2_lut (.I0(GND_net), .I1(n35_adj_3930), .I2(n104_adj_3929), 
            .I3(GND_net), .O(n7982[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3737_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3737_2 (.CI(GND_net), .I0(n35_adj_3930), .I1(n104_adj_3929), 
            .CO(n29480));
    SB_LUT4 add_3736_15_lut (.I0(GND_net), .I1(n7982[12]), .I2(n1050), 
            .I3(n29479), .O(n7966[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3736_14_lut (.I0(GND_net), .I1(n7982[11]), .I2(n977), 
            .I3(n29478), .O(n7966[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_14 (.CI(n29478), .I0(n7982[11]), .I1(n977), .CO(n29479));
    SB_LUT4 add_3736_13_lut (.I0(GND_net), .I1(n7982[10]), .I2(n904), 
            .I3(n29477), .O(n7966[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_13 (.CI(n29477), .I0(n7982[10]), .I1(n904), .CO(n29478));
    SB_LUT4 add_3736_12_lut (.I0(GND_net), .I1(n7982[9]), .I2(n831), .I3(n29476), 
            .O(n7966[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_12 (.CI(n29476), .I0(n7982[9]), .I1(n831), .CO(n29477));
    SB_LUT4 add_3736_11_lut (.I0(GND_net), .I1(n7982[8]), .I2(n758), .I3(n29475), 
            .O(n7966[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_11 (.CI(n29475), .I0(n7982[8]), .I1(n758), .CO(n29476));
    SB_LUT4 add_3736_10_lut (.I0(GND_net), .I1(n7982[7]), .I2(n685), .I3(n29474), 
            .O(n7966[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_10 (.CI(n29474), .I0(n7982[7]), .I1(n685), .CO(n29475));
    SB_LUT4 add_3736_9_lut (.I0(GND_net), .I1(n7982[6]), .I2(n612), .I3(n29473), 
            .O(n7966[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_9 (.CI(n29473), .I0(n7982[6]), .I1(n612), .CO(n29474));
    SB_LUT4 add_3736_8_lut (.I0(GND_net), .I1(n7982[5]), .I2(n539), .I3(n29472), 
            .O(n7966[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_8 (.CI(n29472), .I0(n7982[5]), .I1(n539), .CO(n29473));
    SB_LUT4 add_3736_7_lut (.I0(GND_net), .I1(n7982[4]), .I2(n466), .I3(n29471), 
            .O(n7966[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_7 (.CI(n29471), .I0(n7982[4]), .I1(n466), .CO(n29472));
    SB_LUT4 add_3736_6_lut (.I0(GND_net), .I1(n7982[3]), .I2(n393), .I3(n29470), 
            .O(n7966[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_6 (.CI(n29470), .I0(n7982[3]), .I1(n393), .CO(n29471));
    SB_LUT4 add_3736_5_lut (.I0(GND_net), .I1(n7982[2]), .I2(n320), .I3(n29469), 
            .O(n7966[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_5 (.CI(n29469), .I0(n7982[2]), .I1(n320), .CO(n29470));
    SB_LUT4 add_3736_4_lut (.I0(GND_net), .I1(n7982[1]), .I2(n247), .I3(n29468), 
            .O(n7966[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_4 (.CI(n29468), .I0(n7982[1]), .I1(n247), .CO(n29469));
    SB_LUT4 add_3736_3_lut (.I0(GND_net), .I1(n7982[0]), .I2(n174), .I3(n29467), 
            .O(n7966[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_3 (.CI(n29467), .I0(n7982[0]), .I1(n174), .CO(n29468));
    SB_LUT4 add_3736_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n7966[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3736_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3736_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29467));
    SB_LUT4 add_3735_16_lut (.I0(GND_net), .I1(n7966[13]), .I2(n1120), 
            .I3(n29466), .O(n7949[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3735_15_lut (.I0(GND_net), .I1(n7966[12]), .I2(n1047), 
            .I3(n29465), .O(n7949[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_15 (.CI(n29465), .I0(n7966[12]), .I1(n1047), .CO(n29466));
    SB_LUT4 add_3735_14_lut (.I0(GND_net), .I1(n7966[11]), .I2(n974), 
            .I3(n29464), .O(n7949[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_14 (.CI(n29464), .I0(n7966[11]), .I1(n974), .CO(n29465));
    SB_LUT4 add_3735_13_lut (.I0(GND_net), .I1(n7966[10]), .I2(n901), 
            .I3(n29463), .O(n7949[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_13 (.CI(n29463), .I0(n7966[10]), .I1(n901), .CO(n29464));
    SB_LUT4 add_3735_12_lut (.I0(GND_net), .I1(n7966[9]), .I2(n828), .I3(n29462), 
            .O(n7949[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_12 (.CI(n29462), .I0(n7966[9]), .I1(n828), .CO(n29463));
    SB_LUT4 add_3735_11_lut (.I0(GND_net), .I1(n7966[8]), .I2(n755), .I3(n29461), 
            .O(n7949[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_11 (.CI(n29461), .I0(n7966[8]), .I1(n755), .CO(n29462));
    SB_LUT4 add_3735_10_lut (.I0(GND_net), .I1(n7966[7]), .I2(n682), .I3(n29460), 
            .O(n7949[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_10 (.CI(n29460), .I0(n7966[7]), .I1(n682), .CO(n29461));
    SB_LUT4 add_3735_9_lut (.I0(GND_net), .I1(n7966[6]), .I2(n609), .I3(n29459), 
            .O(n7949[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_9 (.CI(n29459), .I0(n7966[6]), .I1(n609), .CO(n29460));
    SB_LUT4 add_3735_8_lut (.I0(GND_net), .I1(n7966[5]), .I2(n536), .I3(n29458), 
            .O(n7949[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3735_8 (.CI(n29458), .I0(n7966[5]), .I1(n536), .CO(n29459));
    SB_LUT4 add_3735_7_lut (.I0(GND_net), .I1(n7966[4]), .I2(n463), .I3(n29457), 
            .O(n7949[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3735_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4241));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4240));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4239));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4238));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4237));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4236));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4235));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4234));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4232));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4231));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4228));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4227));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3879));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4221));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4219));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4216));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4215));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4213));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4211));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4208));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4207));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4204));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4202));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4201));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4198));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4197));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4196));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4195));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4194));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4193));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4192));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4191));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4190));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4189));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4188));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4187));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4186));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4185));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4184));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4183));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4182));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4181));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4180));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4179));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4178));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4177));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4176));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3868));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4175));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4174));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4173));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33775_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n40606));   // verilog/motorControl.v(46[19:35])
    defparam i33775_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4172));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_3916));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4170));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4169));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4168));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4167));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4166));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4164));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4163));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4161));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4160));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4159));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4158));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4157));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4156));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4155));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4154));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4153));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4152));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4151));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4150));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4149));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4148));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4147));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4146));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4145));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4144));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4142));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4141));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4140));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4139));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4138));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4137));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4135));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4134));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4133));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4132));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4129));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4128));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4126));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4125));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4124));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4123));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4122));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4121));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4120));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4119));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4118));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4117));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4116));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3851));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4115));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4114));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4113));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4112));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4111));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4110));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4109));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4108));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4107));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4106));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4105));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4104));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4103));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4102));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4101));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4100));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4099));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4098));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4097));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4096));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4095));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4094));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4093));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4092));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4091));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4090));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4089));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4088));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4087));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4086));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4085));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4084));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4083));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4082));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4081));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4080));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4079));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4078));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4077));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4076));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4075));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4074));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4073));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4252[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4072));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4071));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4070));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18905_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n3050[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i18905_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4069));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4068));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4066));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i2_3_lut (.I0(n155[1]), .I1(n1[1]), .I2(n256), .I3(GND_net), 
            .O(n3075[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4065));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4064));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4063));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4062));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4061));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4060));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4059));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4058));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256), 
            .I3(GND_net), .O(n3075[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4057));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4056));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4055));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4054));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4053));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4052));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4051));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4048));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4047));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4046));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4045));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4044));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4043));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256), 
            .I3(GND_net), .O(n3075[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_640_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256), 
            .I3(GND_net), .O(n3075[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4042));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4041));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4040));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4039));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256), 
            .I3(GND_net), .O(n3075[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4038));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4037));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256), 
            .I3(GND_net), .O(n3075[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3835));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256), 
            .I3(GND_net), .O(n3075[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4036));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4035));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4033));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4032));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4031));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256), 
            .I3(GND_net), .O(n3075[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4030));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4029));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4028));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4027));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4025));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4024));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256), 
            .I3(GND_net), .O(n3075[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4023));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4022));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4021));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4020));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4019));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4018));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4017));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4016));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4015));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4014));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4013));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4012));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4011));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4010));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4009));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4008));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256), 
            .I3(GND_net), .O(n3075[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256), 
            .I3(GND_net), .O(n3075[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_640_i13_3_lut (.I0(n155[12]), .I1(n1[12]), .I2(n256), 
            .I3(GND_net), .O(n3075[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4007));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4006));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4005));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4004));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4003));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4002));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4001));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4000));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3999));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3998));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3997));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3996));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_3995));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_3993));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_3992));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_3991));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_3990));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3989));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3988));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3987));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_640_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256), 
            .I3(GND_net), .O(n3075[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3986));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_3985));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_3984));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_3983));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_3982));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3981));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3980));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3979));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_640_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256), 
            .I3(GND_net), .O(n3075[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3978));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_3977));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_3976));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_982 (.I0(n6_adj_3922), .I1(\Ki[4] ), .I2(n8378[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8371[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_982.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23039_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n8389[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23039_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_983 (.I0(n4_adj_3940), .I1(\Ki[3] ), .I2(n8384[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8378[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_983.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_3975));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_984 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4246));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_984.LUT_INIT = 16'h9c50;
    SB_LUT4 i22975_4_lut (.I0(n8378[2]), .I1(\Ki[4] ), .I2(n6_adj_3922), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4247));   // verilog/motorControl.v(42[26:37])
    defparam i22975_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_985 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4248));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_985.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23006_4_lut (.I0(n8384[1]), .I1(\Ki[3] ), .I2(n4_adj_3940), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4249));   // verilog/motorControl.v(42[26:37])
    defparam i23006_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23041_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n27720));   // verilog/motorControl.v(42[26:37])
    defparam i23041_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_986 (.I0(n6_adj_4249), .I1(n11_adj_4248), .I2(n8_adj_4247), 
            .I3(n12_adj_4246), .O(n18_adj_4250));   // verilog/motorControl.v(42[26:37])
    defparam i8_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_987 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4251));   // verilog/motorControl.v(42[26:37])
    defparam i3_4_lut_adj_987.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_988 (.I0(n13_adj_4251), .I1(n18_adj_4250), .I2(n27720), 
            .I3(n4_adj_3934), .O(n35988));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33948_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n40780));   // verilog/motorControl.v(44[10:25])
    defparam i33948_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i19188_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n23909));   // verilog/motorControl.v(46[19:35])
    defparam i19188_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3920));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3737[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3737[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3737[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3737[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3737[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3737[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3737[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3737[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3737[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3737[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3737[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3737[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3737[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3737[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3737[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3737[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3737[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3737[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3737[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3737[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3737[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3737[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3737[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3761), .I3(GND_net), .O(duty_23__N_3614[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22985_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n8378[0]));   // verilog/motorControl.v(42[26:37])
    defparam i22985_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_640_i1_4_lut_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n3075[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_640_i1_4_lut_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3944));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33595_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n40425));
    defparam i33595_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i33649_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n40479));
    defparam i33649_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33842_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n40674));
    defparam i33842_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33779_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n40610));
    defparam i33779_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (pwm_setpoint, GND_net, \half_duty_new[0] , 
            CLK_c, PIN_19_c_0, n18061, \half_duty[0][1] , n18062, 
            \half_duty[0][2] , n18063, \half_duty[0][3] , n18064, \half_duty[0][4] , 
            n18066, \half_duty[0][6] , n18067, \half_duty[0][7] , n1172, 
            VCC_net, \half_duty_new[1] , \half_duty[0][0] , \half_duty_new[2] , 
            \half_duty_new[3] , \half_duty_new[4] , \half_duty_new[6] , 
            \half_duty_new[7] , n17424) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input [22:0]pwm_setpoint;
    input GND_net;
    output \half_duty_new[0] ;
    input CLK_c;
    output PIN_19_c_0;
    input n18061;
    output \half_duty[0][1] ;
    input n18062;
    output \half_duty[0][2] ;
    input n18063;
    output \half_duty[0][3] ;
    input n18064;
    output \half_duty[0][4] ;
    input n18066;
    output \half_duty[0][6] ;
    input n18067;
    output \half_duty[0][7] ;
    output n1172;
    input VCC_net;
    output \half_duty_new[1] ;
    output \half_duty[0][0] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n17424;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [22:0]n5595;
    
    wire n27834;
    wire [9:0]half_duty_new_9__N_664;
    
    wire pwm_out_0__N_582, n17004, n27835, n27833, n22157;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    wire [10:0]n49;
    
    wire pause_counter_0__N_612;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n27832, n27831, n35412, pause_counter_0, n27830, n27829, 
        n27828, n27827, n28575, n28574, n28573, n28572, n28571, 
        n28570, n28569, n28568, n28567, n27826, n28566, n27825, 
        n27824, n27823, n27822, n18, n20, n38006, n4, n42408, 
        n42404, pwm_out_0__N_586, n20_adj_3820, n5, n13, n8, n42406, 
        n22, n2, n10, n3, n1, n38116, n13_adj_3821, n12, n18_adj_3822, 
        n3_adj_3823, n16, n20_adj_3824;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n15, n27789, n27788, n27787, n27786;
    wire [10:0]pwm_out_0__N_587;
    
    wire n27785, n27784, n27783, n27782, n27781, n28184, n28183, 
        n28182, n28181, n28180, n28179, n28178, n28177, n28176, 
        n28175, n28174, n28173, n28172, n28171, n28170, n28169, 
        n28168, n27780, n28167, n28166, n28165, n28164, n28163, 
        n27779, n27842, n27841, n27840, n27839, n27838, n27837, 
        n27836;
    
    SB_LUT4 add_2054_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n27834), .O(n5595[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_664[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n17004), .D(pwm_out_0__N_582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2054_15 (.CI(n27834), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n27835));
    SB_LUT4 add_2054_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n27833), .O(n5595[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n18061));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n18062));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n18063));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n18064));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0] [5]), .C(CLK_c), .D(n22157));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n18066));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n18067));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1187__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[10]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[9]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[8]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[7]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[6]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[5]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[4]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[3]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[2]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1187__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[1]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY add_2054_14 (.CI(n27833), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n27834));
    SB_LUT4 add_2054_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n27832), .O(n5595[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_13 (.CI(n27832), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n27833));
    SB_LUT4 add_2054_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n27831), .O(n5595[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_12 (.CI(n27831), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n27832));
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n35412));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_2054_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n27830), .O(n5595[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_11 (.CI(n27830), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n27831));
    SB_LUT4 add_2054_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n27829), .O(n5595[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_10 (.CI(n27829), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n27830));
    SB_LUT4 add_2054_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n27828), .O(n5595[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_9 (.CI(n27828), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n27829));
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_612));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2054_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n27827), .O(n5595[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1187_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n28575), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1187_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n28574), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_11 (.CI(n28574), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n28575));
    SB_LUT4 count_0__1187_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n28573), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_10 (.CI(n28573), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n28574));
    SB_LUT4 count_0__1187_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n28572), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_9 (.CI(n28572), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n28573));
    SB_LUT4 count_0__1187_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n28571), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_8 (.CI(n28571), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n28572));
    SB_LUT4 count_0__1187_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n28570), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_7 (.CI(n28570), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n28571));
    SB_LUT4 count_0__1187_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n28569), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_6 (.CI(n28569), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n28570));
    SB_LUT4 count_0__1187_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n28568), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_5 (.CI(n28568), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n28569));
    SB_LUT4 count_0__1187_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n28567), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_4 (.CI(n28567), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n28568));
    SB_CARRY add_2054_8 (.CI(n27827), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n27828));
    SB_LUT4 add_2054_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n27826), .O(n5595[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_7 (.CI(n27826), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n27827));
    SB_DFFESR count_0__1187__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[0]), .R(n1172));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 count_0__1187_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n28566), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2054_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n27825), .O(n5595[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_6 (.CI(n27825), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n27826));
    SB_LUT4 add_2054_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n27824), .O(n5595[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_5 (.CI(n27824), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n27825));
    SB_LUT4 add_2054_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n27823), .O(n5595[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_4 (.CI(n27823), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n27824));
    SB_CARRY count_0__1187_add_4_3 (.CI(n28566), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n28567));
    SB_LUT4 count_0__1187_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1187_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1187_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n28566));
    SB_LUT4 add_2054_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n27822), .O(n5595[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_3 (.CI(n27822), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n27823));
    SB_LUT4 add_2054_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5595[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n27822));
    SB_LUT4 i9_4_lut (.I0(\count[0] [5]), .I1(n18), .I2(\count[0] [9]), 
            .I3(\count[0] [7]), .O(n20));
    defparam i9_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i7_4_lut (.I0(\count[0] [10]), .I1(\count[0] [4]), .I2(\count[0] [2]), 
            .I3(n38006), .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'h0080;
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_664[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i8_4_lut (.I0(n4), .I1(n42408), .I2(n42404), .I3(pwm_out_0__N_586), 
            .O(n20_adj_3820));
    defparam i8_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut (.I0(\count[0] [10]), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n13));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10_4_lut (.I0(n13), .I1(n20_adj_3820), .I2(n8), .I3(n42406), 
            .O(n22));
    defparam i10_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i31350_4_lut (.I0(n2), .I1(n10), .I2(n3), .I3(n1), .O(n38116));
    defparam i31350_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n38116), .I1(pause_counter_0), .I2(pwm_out_0__N_582), 
            .I3(n22), .O(n17004));
    defparam i1_4_lut.LUT_INIT = 16'h1303;
    SB_LUT4 i2_4_lut (.I0(\count[0] [6]), .I1(\count[0] [5]), .I2(\half_duty[0][6] ), 
            .I3(\half_duty[0] [5]), .O(n13_adj_3821));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut (.I0(\half_duty[0][3] ), .I1(\count[0] [10]), .I2(\count[0] [3]), 
            .I3(GND_net), .O(n12));   // vhdl/pwm.vhd(80[8:31])
    defparam i1_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i7_4_lut_adj_969 (.I0(n13_adj_3821), .I1(\half_duty[0][7] ), 
            .I2(\count[0] [9]), .I3(\count[0] [7]), .O(n18_adj_3822));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_4_lut_adj_969.LUT_INIT = 16'hfbfe;
    SB_LUT4 half_duty_0__9__I_0_47_i3_2_lut (.I0(\half_duty[0][2] ), .I1(\count[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3823));   // vhdl/pwm.vhd(80[8:31])
    defparam half_duty_0__9__I_0_47_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\half_duty[0][1] ), .I1(\count[0] [0]), .I2(\count[0] [1]), 
            .I3(\half_duty[0][0] ), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9_4_lut_adj_970 (.I0(\half_duty[0][4] ), .I1(n18_adj_3822), 
            .I2(n12), .I3(\count[0] [4]), .O(n20_adj_3824));   // vhdl/pwm.vhd(80[8:31])
    defparam i9_4_lut_adj_970.LUT_INIT = 16'hfdfe;
    SB_LUT4 i10_4_lut_adj_971 (.I0(\count[0] [8]), .I1(n20_adj_3824), .I2(n16), 
            .I3(n3_adj_3823), .O(pwm_out_0__N_582));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_971.LUT_INIT = 16'hfffe;
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_664[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_664[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_664[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(half_duty_new[5]), .C(CLK_c), .D(half_duty_new_9__N_664[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_664[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_664[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n17424));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i4_2_lut (.I0(\count[0] [1]), .I1(\count[0] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n15));
    defparam i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10_4_lut_adj_972 (.I0(n15), .I1(n20), .I2(\count[0] [8]), 
            .I3(\count[0] [3]), .O(n1172));
    defparam i10_4_lut_adj_972.LUT_INIT = 16'h0800;
    SB_CARRY pwm_out_0__I_20_13 (.CI(n27789), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_586));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n27788), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27789));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n27787), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n27787), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27788));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n27786), .O(n42408)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_10 (.CI(n27786), .I0(GND_net), .I1(VCC_net), 
            .CO(n27787));
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_587[7]), 
            .I3(n27785), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n27785), .I0(GND_net), .I1(pwm_out_0__N_587[7]), 
            .CO(n27786));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_587[6]), 
            .I3(n27784), .O(n42404)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n27784), .I0(VCC_net), .I1(pwm_out_0__N_587[6]), 
            .CO(n27785));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_587[5]), 
            .I3(n27783), .O(n42406)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n27783), .I0(GND_net), .I1(pwm_out_0__N_587[5]), 
            .CO(n27784));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_587[4]), 
            .I3(n27782), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n27782), .I0(GND_net), .I1(pwm_out_0__N_587[4]), 
            .CO(n27783));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_587[3]), 
            .I3(n27781), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_2043_24_lut (.I0(GND_net), .I1(n5595[22]), .I2(pwm_setpoint[22]), 
            .I3(n28184), .O(half_duty_new_9__N_664[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2043_23_lut (.I0(GND_net), .I1(n5595[21]), .I2(pwm_setpoint[21]), 
            .I3(n28183), .O(half_duty_new_9__N_664[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_23 (.CI(n28183), .I0(n5595[21]), .I1(pwm_setpoint[21]), 
            .CO(n28184));
    SB_LUT4 add_2043_22_lut (.I0(GND_net), .I1(n5595[20]), .I2(pwm_setpoint[20]), 
            .I3(n28182), .O(half_duty_new_9__N_664[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_22 (.CI(n28182), .I0(n5595[20]), .I1(pwm_setpoint[20]), 
            .CO(n28183));
    SB_LUT4 add_2043_21_lut (.I0(GND_net), .I1(n5595[19]), .I2(pwm_setpoint[19]), 
            .I3(n28181), .O(half_duty_new_9__N_664[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_21 (.CI(n28181), .I0(n5595[19]), .I1(pwm_setpoint[19]), 
            .CO(n28182));
    SB_LUT4 add_2043_20_lut (.I0(GND_net), .I1(n5595[18]), .I2(pwm_setpoint[18]), 
            .I3(n28180), .O(half_duty_new_9__N_664[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n27781), .I0(GND_net), .I1(pwm_out_0__N_587[3]), 
            .CO(n27782));
    SB_CARRY add_2043_20 (.CI(n28180), .I0(n5595[18]), .I1(pwm_setpoint[18]), 
            .CO(n28181));
    SB_LUT4 add_2043_19_lut (.I0(GND_net), .I1(n5595[17]), .I2(pwm_setpoint[17]), 
            .I3(n28179), .O(half_duty_new_9__N_664[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_19 (.CI(n28179), .I0(n5595[17]), .I1(pwm_setpoint[17]), 
            .CO(n28180));
    SB_LUT4 add_2043_18_lut (.I0(GND_net), .I1(n5595[16]), .I2(pwm_setpoint[16]), 
            .I3(n28178), .O(half_duty_new_9__N_664[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_18 (.CI(n28178), .I0(n5595[16]), .I1(pwm_setpoint[16]), 
            .CO(n28179));
    SB_LUT4 add_2043_17_lut (.I0(GND_net), .I1(n5595[15]), .I2(pwm_setpoint[15]), 
            .I3(n28177), .O(half_duty_new_9__N_664[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2043_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2043_17 (.CI(n28177), .I0(n5595[15]), .I1(pwm_setpoint[15]), 
            .CO(n28178));
    SB_CARRY add_2043_16 (.CI(n28176), .I0(n5595[14]), .I1(pwm_setpoint[14]), 
            .CO(n28177));
    SB_CARRY add_2043_15 (.CI(n28175), .I0(n5595[13]), .I1(pwm_setpoint[13]), 
            .CO(n28176));
    SB_CARRY add_2043_14 (.CI(n28174), .I0(n5595[12]), .I1(pwm_setpoint[12]), 
            .CO(n28175));
    SB_CARRY add_2043_13 (.CI(n28173), .I0(n5595[11]), .I1(pwm_setpoint[11]), 
            .CO(n28174));
    SB_CARRY add_2043_12 (.CI(n28172), .I0(n5595[10]), .I1(pwm_setpoint[10]), 
            .CO(n28173));
    SB_CARRY add_2043_11 (.CI(n28171), .I0(n5595[9]), .I1(pwm_setpoint[9]), 
            .CO(n28172));
    SB_CARRY add_2043_10 (.CI(n28170), .I0(n5595[8]), .I1(pwm_setpoint[8]), 
            .CO(n28171));
    SB_CARRY add_2043_9 (.CI(n28169), .I0(n5595[7]), .I1(pwm_setpoint[7]), 
            .CO(n28170));
    SB_CARRY add_2043_8 (.CI(n28168), .I0(n5595[6]), .I1(pwm_setpoint[6]), 
            .CO(n28169));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_587[2]), 
            .I3(n27780), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2043_7 (.CI(n28167), .I0(n5595[5]), .I1(pwm_setpoint[5]), 
            .CO(n28168));
    SB_CARRY add_2043_6 (.CI(n28166), .I0(n5595[4]), .I1(pwm_setpoint[4]), 
            .CO(n28167));
    SB_CARRY add_2043_5 (.CI(n28165), .I0(n5595[3]), .I1(pwm_setpoint[3]), 
            .CO(n28166));
    SB_CARRY add_2043_4 (.CI(n28164), .I0(n5595[2]), .I1(pwm_setpoint[2]), 
            .CO(n28165));
    SB_CARRY add_2043_3 (.CI(n28163), .I0(n5595[1]), .I1(pwm_setpoint[1]), 
            .CO(n28164));
    SB_CARRY add_2043_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n28163));
    SB_CARRY pwm_out_0__I_20_4 (.CI(n27780), .I0(GND_net), .I1(pwm_out_0__N_587[2]), 
            .CO(n27781));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_587[1]), 
            .I3(n27779), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_3 (.CI(n27779), .I0(GND_net), .I1(pwm_out_0__N_587[1]), 
            .CO(n27780));
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_587[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_587[0]), 
            .CO(n27779));
    SB_LUT4 add_2054_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n27842), .O(n5595[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2054_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n27841), .O(n5595[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_22 (.CI(n27841), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n27842));
    SB_LUT4 add_2054_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n27840), .O(n5595[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_21 (.CI(n27840), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n27841));
    SB_LUT4 add_2054_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n27839), .O(n5595[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_20 (.CI(n27839), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n27840));
    SB_LUT4 add_2054_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n27838), .O(n5595[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_19 (.CI(n27838), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n27839));
    SB_LUT4 add_2054_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n27837), .O(n5595[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_18 (.CI(n27837), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n27838));
    SB_LUT4 add_2054_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n27836), .O(n5595[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_17 (.CI(n27836), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n27837));
    SB_LUT4 add_2054_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n27835), .O(n5595[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2054_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2054_16 (.CI(n27835), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n27836));
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36306_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_582), .I2(GND_net), 
            .I3(GND_net), .O(n35412));
    defparam i36306_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0] [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17436_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1172), .I3(GND_net), .O(n22157));
    defparam i17436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17444_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_out_0__N_587[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i17444_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31240_2_lut (.I0(pause_counter_0), .I1(\count[0] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n38006));
    defparam i31240_2_lut.LUT_INIT = 16'heeee;
    
endmodule
