// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Feb  1 10:54:27 2022
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    
    wire n1767;
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    
    wire n41195;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(353[11:24])
    
    wire n59929;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(361[15:20])
    
    wire pwm_setpoint_23__N_207, n11439, n11441, n11443, n11445, n11447, 
        n11449, n11451, n11453, n11455, n11457, n11459, n11461, 
        n11463, n11465, n11467, n11469, n60023, n260, n11477, 
        n11475, n294, n298, n299, n300, n301, n302, n303, n304, 
        n305, n306, n307, n308, n309;
    wire [23:0]pwm_setpoint_23__N_3;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    
    wire n71355, n1769, n1771, n1773;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, n32202, RX_N_2, n1765, n1763, n1761, n1759, 
        n68483, n1757, n1755;
    wire [31:0]motor_state_23__N_91;
    wire [44:0]encoder1_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
        read_N_409, n1331, n21540, n21539, n62, n6, n26, n68937, 
        n1805;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    wire [5:0]color_bit_N_502;
    
    wire n70437, n25, n24, n23, n22, n21, n20, n19, n32199, 
        n19_adj_5734, n17, n16, n15, n13, n11, n9, n18, n17_adj_5735, 
        n2834, n16_adj_5736, n15_adj_5737, n14, n13_adj_5738, n52728, 
        n2, n14_adj_5739, n15_adj_5740, n16_adj_5741, n17_adj_5742, 
        n18_adj_5743, n19_adj_5744, n20_adj_5745, n21_adj_5746, n22_adj_5747, 
        n23_adj_5748, n24_adj_5749, n25_adj_5750, n24_adj_5751, n15015, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n4943, n4942, n4941, n4921, 
        n4920, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
        n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, 
        n4937, n4938, n4939, n4940, n59928, n3489, n2887, n65, 
        n12, n40902, n40859, n70408, n40795, n62546, n1, n52711, 
        n52727, n52710, n52726, n52709, n59932, n70680, n35072, 
        n52725, n52724, n52723, n71337, n8, n20277, Kp_23__N_869, 
        n69780, Kp_23__N_715, n70104, n15_adj_5752, n13533, n8_adj_5753, 
        n68877, n69736, n69750, n32171, \FRAME_MATCHER.i_31__N_2509 , 
        \FRAME_MATCHER.i_31__N_2513 , n54060, n39619, n54059, n54058, 
        n32168, n32165, n61815, n32162, n32158, n32155, n32152, 
        n32149, n32146, n32143, n32140, n32137, n32134, n32130, 
        n32127, n32124, n32109, n32068, n32065, n32062, n32059, 
        n32056, n32053, n32050, n32047, n32044, n32041, n59777, 
        n32038, n32028, n32018, n32015, n32012, n32009, n32005, 
        n54057, n54056, n11890, n53495, n54055, n54054, n54053, 
        n54052, n31925, n31922, n31919, n31916, n31915, n31914, 
        n31913, n31912, n31911, n31910, n31909, n31908, n31907, 
        n31906, n31874, n31873, n31872, n31871, n31870, n31869, 
        n31868, n31867, n31866, n31865, n31864, n31863, n31862, 
        n31861, n31860, n31859, n31858, n31857, n31856, n31853, 
        n31821, n31820, n31819, n31818, n31817, n31811, n31806, 
        n54051, n31802, n54050, n31796, n31793, n31787, n31784, 
        n54049, n54048, n54047, n53494, n54046, n53493, n54045, 
        n54044, n31772, n54043, n53492, n31766, n54042, n7, n6_adj_5754, 
        n5, n4, n24_adj_5755, n21_adj_5756, n19_adj_5757, n17_adj_5758, 
        n15_adj_5759, n53491, n54041, n54040, n53490, n54039, n53489, 
        n54038, n54037, n54036, n54035, n54034, n54033, n54032, 
        n54031, n54030, n14_adj_5760, n12_adj_5761, n10, n54029, 
        n4_adj_5762, n54028, n40, n70436, n70422, n30, n23_adj_5763, 
        n22_adj_5764, n21_adj_5765, n19_adj_5766, n17_adj_5767, n16_adj_5768, 
        n15_adj_5769, n13_adj_5770, n11_adj_5771, n10_adj_5772, n9_adj_5773, 
        n8_adj_5774, n7_adj_5775, n6_adj_5776, n4_adj_5777, n54027, 
        n54026, n54025, n54024, n54023, n54022, n54021, n54020, 
        n54019, n54018, n54017, n59927, n59926, n59925, n59924, 
        n59923, n60028, n59934, n60029, n59922, n54016, n54015, 
        n54014, n54013, n54012, n15_adj_5778, n54011, n54010, n54009, 
        n54008, n54007, n54006, n54005, n59921, n60031, n59920, 
        n59919, n59918, n59917, n54004, n4_adj_5779, n54003, n4_adj_5780, 
        n54002, n4_adj_5781, n54001, n54000, n53999, n27754, n53998, 
        n10_adj_5782, n53997, n70124, n53996, n53995, n53994, n53993, 
        n53992, n53991, n53990, n53989, n53988, control_update, 
        n53987, n53986;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n53985, n53984, n59916, n53983, n32704, n55760, n53982, 
        n53981, n11437, n53980, n59915, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344, n345, n346, n347, n348, 
        n349, n350, n351, n352, n353, n354, n355, n356, n357, 
        n358, n359, n53979, n53978, n53977, n53976, n5233, n5230, 
        n53975, n53974, n31757, n3178, n31754, n59914, n5_adj_5783, 
        n32677, n32676, n32675, n32674, n32673, n32672, n32671, 
        n32670, n32669, n11_adj_5784, n32668, n32667, n32666, n32665, 
        n32663;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, position_31__N_3836, n53967, 
        n53966, n70112, n70672, n70119, n32651, n32650, n32649, 
        n25253, n53965, n52722, n15_adj_5785, n32645, n32644, n53964, 
        n32640, n53963;
    wire [1:0]a_new_adj_5905;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5906;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5788, b_prev_adj_5789, debounce_cnt_N_3833_adj_5790, 
        n32632, position_31__N_3836_adj_5791, n70311, n53962, n20276, 
        n53961, n20274, n64704, n53960, n59265, n12_adj_5792, n11_adj_5793, 
        n10_adj_5794, n4_adj_5795, n3, n2_adj_5796, n53959;
    wire [7:0]data_adj_5919;   // verilog/eeprom.v(23[12:16])
    
    wire n30278;
    wire [7:0]state_7__N_3918;
    
    wire n53958, n52962, n52961, n53957, n31751, n53956, n53955, 
        n53954, n53953, n53952, n53951, n53950, n53949, n52960, 
        n52959, n31748, n5_adj_5797, n31745, n14_adj_5798, n53948, 
        n60030, n52958, n53947, n13_adj_5799, n52957, n6916, n53946, 
        n32606, n32605, n52956, n32604, n32603, n70111, n32600, 
        n32599, n32598, n53945, n32594, n32593, n27752, n52955, 
        n53944, n52954, n53943, n52953, n52952, n32592, n53942, 
        n52951, n32591, n53941, n32590, n32589, n32588, n32587, 
        n53940, n27938, n32586, n52950;
    wire [15:0]data_adj_5926;   // verilog/tli4970.v(27[14:18])
    
    wire n53939, n53938, n32585, n53937, n53936, n32584, n32583, 
        n32582, n32581, n32580, n32579, n32578, n53935, n32577, 
        n32576, n32575, n32574, n32573, n32570, n53934, n53933, 
        n53932, n53931, n15_adj_5808, n52721, n53930, n52720, n5_adj_5809, 
        n53929, n31742, n40832, n11471, n31739, n11473, n53928, 
        state_7__N_4319, n61776, n70115, n9_adj_5810, n8_adj_5811, 
        n7_adj_5812, n6_adj_5813, n5_adj_5814, n53927, n27749, n53926, 
        r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n8_adj_5815, n53925, n53924, n31736, n53923;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n71313, n71307, n53922;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n53921, n17531, n52708, n69776, n32489, n32488, n32487, 
        n32484, n32483, n32482, n32481, n32480, n53920;
    wire [2:0]r_SM_Main_adj_5942;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5943;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5944;   // verilog/uart_tx.v(34[16:27])
    
    wire n53919, n32479, n32478, n32477, n32475, n32474;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n32472, n32471, n32470, n32469, n32468, n32467, n32462, 
        n32461, n32460, n32459, n32458, n32457, n32455, n32454, 
        n32452, n32451, n32450;
    wire [7:0]state_adj_5952;   // verilog/i2c_controller.v(33[12:17])
    
    wire n32449, n32448, n32447, n32446, n32445, n32444, n21523, 
        n6720;
    wire [7:0]state_7__N_4126;
    
    wire n32409, n32406, n32403, n32396, n32393, n32390, n32387, 
        n20278, n59913, n60038, n60044, n60043, n59912, n53891, 
        n30237, n59911, n60042, n59910, n60041, n59909, n60046, 
        n60045, n59908, n53890, n60025, n60047, n53889, n59907, 
        n30217, n59906, n53888, n53887, n59931, n53886, n60039, 
        n59905, n59904, n59903, n59902, n59901, n60024, n53885, 
        n43, n53884, n53883, n31492, n59900, n31490, n53882, n53881, 
        n59939, n59899, n59898, n53880, n53879, n53878, n53877, 
        n53876, n60026, n59897, n60035, n59896, n59895, n59930, 
        n31484, n53875, n53874, n53873, n67418, n53872, n53871, 
        n21531, n20279, n60609, n17525, n21537, n17532, n15009, 
        n13527, n11884, n59938, n15016, n13534, n11891, n10009, 
        n21532, n17526, n59894, n59935, n17533, n11885, n13528, 
        n15010, n21533, n59893, n32363, n20280, n59892, n59891, 
        n15017, n13535, n11892, n59890, n64710, n17527, n21534, 
        n64707, n59772, n11886, n4_adj_5829, n15011, n13529, n17534, 
        n15018, n59889, n71301, n20281, n13536, n11893, n53792, 
        n52719, n52707, n53791, n53790, n53789, n53788, n17528, 
        n21535, n11887, n53787, n53786, n13530, n53785, n53784, 
        n15012, n53783, n53782, n53781, n53780, n53779, n64705, 
        n17535, n53778, n53777, n52718, n53776, n53775, n15019, 
        n13537, n11894, n53774, n52880, n17529, n20282, n53773, 
        n52879, n52878, n11888, n13531, n52877, n52876, n15013, 
        n71295, n52875, n52874, n28460, n52873, n52872, n59888, 
        n60051, n52871, n52870, n52869, n52868, n15020, n37892, 
        n13538, n11895, n59798, n52867, n59887, n17530, n52866, 
        n52706, n30137, n37917, n52865, n52864, n69468, n21520, 
        n20275, n27881, n20283, n31475, n60049, n31474, n30093, 
        n30087, n4_adj_5830, n6_adj_5831, n8_adj_5832, n9_adj_5833, 
        n11_adj_5834, n13_adj_5835, n14_adj_5836, n15_adj_5837, n30084, 
        n4_adj_5838, n6_adj_5839, n8_adj_5840, n9_adj_5841, n59886, 
        n30080, n52863, n55567, n60050, n30062, n60048, n52862, 
        n17515, n38, n39, n40_adj_5842, n41, n42, n43_adj_5843, 
        n44, n45, n55, n11897, n30039, n59885, n21521, n31471, 
        n55737, n30015, n69830, n31470, n59884, n59883, n31467, 
        n60040, n59882, n59881, n59880, n59879, n60021, n59874, 
        n60037, n60022, n31461, n60036, n29991, n52861, n52860, 
        n52859, n52858, n55781, n55748, n55746, n31653, n31460, 
        n60020, n59878, n60019, n59877, n60018, n59876, n60017, 
        n60016, n31455, n60015, n60082, n60014, n60081, n60013, 
        n60077, n60012, n31451, n60011, n60078, n60010, n60076, 
        n60009, n60073, n60008, n31447, n60007, n60074, n60006, 
        n60079, n60005, n60080, n60004, n31443, n60003, n60072, 
        n60002, n60075, n60001, n60000, n59999, n59998, n59997, 
        n59996, n59995, n59994, n59993, n59992, n59991, n59990, 
        n59989, n59988, n59987, n59986, n59985, n59984, n59983, 
        n59982, n59981, n59980, n59979, n59978, n59977, n59976, 
        n59975, n59974, n59973, n59972, n59936, n59971, n59970, 
        n59969, n59968, n59967, n59966, n59965, n59964, n59963, 
        n59962, n59961, n59960, n59959, n59958, n59957, n59956, 
        n59955, n59954, n59953, n59952, n62587, n59951, n59950, 
        n59949, n59948, n59947, n59875, n59946, n31358, n59945, 
        n59944, n59943, n59942, n59941, n59940, n30709, n30708, 
        n30702, n30700, n30698, n59789, n59773, n59779, n60134, 
        n30673, n30671, n30669, n40695, n31122, n30629, n30627, 
        n30623, n30621, n30619, n60027, n20284, n21538, n21522, 
        n60033, n20285, n9946, n9944, n13517, n11874, n14999, 
        n20286, n17517, n13518, n4_adj_5844, n15000, n11875, n17516, 
        n71265, n71253, n59313, n11876, n13519, n15001, n25082, 
        n11877, n13520, n15002, n17518, n15003, n17519, n32306, 
        n11879, n13522, n15004, n17520, n71703, n11878, n13521, 
        n71229, n71223, n71220, n71217, n59937, n6_adj_5845, n32300, 
        n32299, n15005, n17521, n32290, n32286, n11880, n13523, 
        n31708, n31707, n27930, n32278, n55802, n32272, n17522, 
        n11881, n15006, n13524, n31706, n31705, n31699, n11882, 
        n13525, n15007, n21524, n17523, n59315, n32250, n52826, 
        n21536, n17524, n31695, n31693, n11883, n13526, n15008, 
        n52825, n59203, n59933, n20287, n52824, n71697, n21525, 
        n11896, n13539, n52823, n20288, n27925, n21526, n20289, 
        n21527, n20290, n21528, n20291, n21529, n20292, n21530, 
        n15014, n27891, n10_adj_5846, n52717, n11435, n7_adj_5847, 
        n64584, n55267, n13511, n11868, n6_adj_5848, n60150, n27360, 
        n14994, n13512, n11869, n64411, n13532, n14995, n13513, 
        n11870, n17512, n14996, n25151, n13514, n71658, n55993, 
        n11871, n71655, n17513, n14997, n13515, n11872, n54840, 
        n11889, n17514, n71628, n14998, n13516, n11873, n60538, 
        n24010, n24006, n52822, n68976, n60034, n60032, n20293, 
        n20294, n20295, n52716, n52821, n6_adj_5849, n52820, n52819, 
        n52715, n52818, n52817, n52816, n52815, n52814, n27916, 
        n68947, n27889, n52813, n68944, n52812, n52811, n52714, 
        n52810, n52809, n52734, n64581, n64815, n52808, n52807, 
        n52733, n52705, n15_adj_5850, n14_adj_5851, n64809, n39602, 
        n39603, n52806, n52805, n52804, n89, n52732, n52731, n39634, 
        n30323, n41236, n40683, n76, n52704, n31682, n52713, n52712, 
        n52730, n52729, n71737, n68869, n68851, n62287, n71580, 
        n61124, n71397, n70310, n71391, n63671, n71577, n14_adj_5852, 
        n64493, n71574, n64491, n10_adj_5853, n63653, n70420, n71385, 
        n63647, n63641, n63635, n63629, n17_adj_5854, n25_adj_5855, 
        n58271, n24_adj_5856, n63623, n63621, n63617, n71379, n63611, 
        n60952, n58351, n63605, n68541, n63599, n63593, n63587, 
        n62692, n63581, n63575, n8_adj_5857, n7_adj_5858, n68520, 
        n63569, n63563, n68512, n22_adj_5859, n60927, n71373, n60925, 
        n63557, n70409, n29, n27, n63551, n67794, n63549, n67793, 
        n23_adj_5860, n63545, n63539, n67782, n63533, n63527, n70740, 
        n6_adj_5861, n63521, n60071, n60414, n63515, n62946, n15_adj_5862, 
        n14_adj_5863, n67745, n61810, n59873, n67713, n67710, n67702, 
        n67701, n67698, n64415, n67697, n64585, n64582, n70888, 
        n4_adj_5864, n70887, n70860, n70859, n59083, n59095, n64465, 
        n59173, n59177, n59181, n59185, n59189, n59193, n59197, 
        n59201, n63279, n70861, n64882, n60086, n64881, n60523, 
        n59255, n59263, n63273, n63269, n71349, n63263, n67938, 
        n59309, n63257, n63255, n6_adj_5865, n8_adj_5866, n60514, 
        n70733, n68883, n71523, n70739, n64817, n67874, n64816, 
        n67604, n64811, n64810, n70639, n71784, n71367, n67858, 
        n59473, n64579, n64578, n70756, n64802, n71361, n67843, 
        n4_adj_5867, n67567, n70096, n64407, n62632, n63077, n63069, 
        n7_adj_5868, n7_adj_5869, n67541;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n29991), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i13824_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n59773), 
            .I3(GND_net), .O(n32015));   // verilog/coms.v(130[12] 305[6])
    defparam i13824_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n9946_bdd_4_lut (.I0(n9946), .I1(current[1]), .I2(duty[4]), 
            .I3(n9944), .O(n71703));
    defparam n9946_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n52860), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13827_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n59773), 
            .I3(GND_net), .O(n32018));   // verilog/coms.v(130[12] 305[6])
    defparam i13827_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .n67418(n67418), 
            .GND_net(GND_net), .bit_ctr({Open_0, bit_ctr[3], Open_1, 
            bit_ctr[1:0]}), .n40859(n40859), .n54840(n54840), .\color_bit_N_502[1] (color_bit_N_502[1]), 
            .n30217(n30217), .state({state}), .n27360(n27360), .\neopxl_color[9] (neopxl_color[9]), 
            .\neopxl_color[8] (neopxl_color[8]), .\neopxl_color[5] (neopxl_color[5]), 
            .\neopxl_color[4] (neopxl_color[4]), .timer({timer}), .LED_c(LED_c), 
            .VCC_net(VCC_net), .n32028(n32028), .n59083(n59083), .\bit_ctr[4] (bit_ctr[4]), 
            .n31915(n31915), .t0({t0}), .n31914(n31914), .n31913(n31913), 
            .n31912(n31912), .n31911(n31911), .n31910(n31910), .n31909(n31909), 
            .n31908(n31908), .n31907(n31907), .n31906(n31906), .NEOPXL_c(NEOPXL_c), 
            .n31708(n31708), .\neopxl_color[14] (neopxl_color[14]), .\neopxl_color[15] (neopxl_color[15]), 
            .\neopxl_color[12] (neopxl_color[12]), .\neopxl_color[13] (neopxl_color[13]), 
            .n71658(n71658), .\neopxl_color[20] (neopxl_color[20]), .\neopxl_color[22] (neopxl_color[22]), 
            .\neopxl_color[21] (neopxl_color[21]), .\neopxl_color[23] (neopxl_color[23]), 
            .\neopxl_color[17] (neopxl_color[17]), .\neopxl_color[19] (neopxl_color[19]), 
            .\neopxl_color[16] (neopxl_color[16]), .\neopxl_color[18] (neopxl_color[18]), 
            .n3178(n3178), .\neopxl_color[6] (neopxl_color[6]), .\neopxl_color[7] (neopxl_color[7]), 
            .\neopxl_color[10] (neopxl_color[10]), .\neopxl_color[11] (neopxl_color[11])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 n71703_bdd_4_lut (.I0(n71703), .I1(duty[1]), .I2(n4942), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n71703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n52706), .O(n1248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n52860), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n52861));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n52859), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_14 (.CI(n52715), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n52716));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n52859), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n52860));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n52858), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19749_3_lut (.I0(n37892), .I1(current[4]), .I2(current_limit[4]), 
            .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i19749_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i50815_3_lut (.I0(n10), .I1(current_limit[8]), .I2(n17_adj_5758), 
            .I3(GND_net), .O(n70310));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n27754));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1795 (.I0(ID[3]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5798));   // verilog/TinyFPGA_B.v(379[12:17])
    defparam i6_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1796 (.I0(ID[0]), .I1(ID[1]), .I2(ID[7]), .I3(ID[2]), 
            .O(n13_adj_5799));   // verilog/TinyFPGA_B.v(379[12:17])
    defparam i5_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 n9946_bdd_4_lut_52117 (.I0(n9946), .I1(current[0]), .I2(duty[3]), 
            .I3(n9944), .O(n71697));
    defparam n9946_bdd_4_lut_52117.LUT_INIT = 16'he4aa;
    SB_LUT4 i22603_4_lut (.I0(n13_adj_5799), .I1(baudrate[0]), .I2(n14_adj_5798), 
            .I3(n27889), .O(n40695));
    defparam i22603_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i1_2_lut (.I0(delay_counter[12]), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5829));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5829), .I2(delay_counter[10]), 
            .I3(n27752), .O(n62287));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1797 (.I0(n62287), .I1(n27749), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n62587));
    defparam i2_4_lut_adj_1797.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5857));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1798 (.I0(delay_counter[22]), .I1(n62587), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5858));
    defparam i2_4_lut_adj_1798.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22632_4_lut (.I0(n7_adj_5858), .I1(delay_counter[31]), .I2(n27754), 
            .I3(n8_adj_5857), .O(n1331));   // verilog/TinyFPGA_B.v(381[14:38])
    defparam i22632_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n27749));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[6]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5863));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n71697_bdd_4_lut (.I0(n71697), .I1(duty[0]), .I2(n4943), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n71697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1799 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[0]), .I3(delay_counter[3]), .O(n15_adj_5862));
    defparam i6_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5862), .I1(delay_counter[1]), .I2(n14_adj_5863), 
            .I3(delay_counter[2]), .O(n27752));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4290_4_lut (.I0(n27752), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5751));
    defparam i4290_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1800 (.I0(n24_adj_5751), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n62632));
    defparam i2_4_lut_adj_1800.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1801 (.I0(n62632), .I1(delay_counter[18]), .I2(n27749), 
            .I3(GND_net), .O(n62546));
    defparam i2_3_lut_adj_1801.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1802 (.I0(delay_counter[23]), .I1(n62546), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5868));
    defparam i2_4_lut_adj_1802.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5868), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n27754), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22702_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(367[12:35])
    defparam i22702_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6165_3_lut (.I0(n4920), .I1(current[15]), .I2(n9944), .I3(GND_net), 
            .O(n24010));
    defparam i6165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6166_3_lut (.I0(n24010), .I1(duty[23]), .I2(n9946), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i6166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i589_2_lut (.I0(n1331), .I1(n40695), .I2(GND_net), .I3(GND_net), 
            .O(n2834));   // verilog/TinyFPGA_B.v(385[18] 387[12])
    defparam i589_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i44979_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64465));
    defparam i44979_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51676_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6916), .I2(n64465), 
            .I3(n25_adj_5855), .O(n17_adj_5854));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i51676_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i50816_3_lut (.I0(n70310), .I1(current_limit[9]), .I2(n19_adj_5757), 
            .I3(GND_net), .O(n70311));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48967_4_lut (.I0(bit_ctr[0]), .I1(n67418), .I2(n54840), .I3(color_bit_N_502[1]), 
            .O(n67745));   // verilog/neopixel.v(34[12] 113[6])
    defparam i48967_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i26_4_lut (.I0(n27360), .I1(n67745), .I2(state[1]), .I3(n4_adj_5844), 
            .O(n59083));   // verilog/neopixel.v(34[12] 113[6])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i13734_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n60134), 
            .I3(GND_net), .O(n31925));   // verilog/coms.v(130[12] 305[6])
    defparam i13734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13731_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n60134), 
            .I3(GND_net), .O(n31922));   // verilog/coms.v(130[12] 305[6])
    defparam i13731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13728_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n60134), 
            .I3(GND_net), .O(n31919));   // verilog/coms.v(130[12] 305[6])
    defparam i13728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13725_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n60134), 
            .I3(GND_net), .O(n31916));   // verilog/coms.v(130[12] 305[6])
    defparam i13725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13662_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n60134), 
            .I3(GND_net), .O(n31853));   // verilog/coms.v(130[12] 305[6])
    defparam i13662_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n52858), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n52859));
    SB_LUT4 i13620_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n60134), 
            .I3(GND_net), .O(n31811));   // verilog/coms.v(130[12] 305[6])
    defparam i13620_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25), .CO(n52858));
    SB_LUT4 i13615_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n60134), 
            .I3(GND_net), .O(n31806));   // verilog/coms.v(130[12] 305[6])
    defparam i13615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13847_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n59773), 
            .I3(GND_net), .O(n32038));   // verilog/coms.v(130[12] 305[6])
    defparam i13847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13850_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n59773), 
            .I3(GND_net), .O(n32041));   // verilog/coms.v(130[12] 305[6])
    defparam i13850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13955_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n59777), .I3(GND_net), .O(n32146));   // verilog/coms.v(130[12] 305[6])
    defparam i13955_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13853_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n59773), 
            .I3(GND_net), .O(n32044));   // verilog/coms.v(130[12] 305[6])
    defparam i13853_3_lut.LUT_INIT = 16'hacac;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n71655_bdd_4_lut (.I0(n71655), .I1(neopxl_color[2]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[0]), .O(n71658));
    defparam n71655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13856_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n59772), .I3(GND_net), .O(n32047));   // verilog/coms.v(130[12] 305[6])
    defparam i13856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13859_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n59772), .I3(GND_net), .O(n32050));   // verilog/coms.v(130[12] 305[6])
    defparam i13859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49973_4_lut (.I0(n19_adj_5757), .I1(n17_adj_5758), .I2(n15_adj_5759), 
            .I3(n68483), .O(n69468));
    defparam i49973_4_lut.LUT_INIT = 16'heeef;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13862_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n59772), .I3(GND_net), .O(n32053));   // verilog/coms.v(130[12] 305[6])
    defparam i13862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13865_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n59772), .I3(GND_net), .O(n32056));   // verilog/coms.v(130[12] 305[6])
    defparam i13865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i14_3_lut (.I0(n12_adj_5761), .I1(current_limit[7]), 
            .I2(n15_adj_5759), .I3(GND_net), .O(n14_adj_5760));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i13868_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n59772), .I3(GND_net), .O(n32059));   // verilog/coms.v(130[12] 305[6])
    defparam i13868_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i1_3_lut (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), .I2(n5233), 
            .I3(GND_net), .O(n63077));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), .I3(n63077), 
            .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_1181_i15_2_lut (.I0(r_Clock_Count_adj_5943[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5837));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i9_2_lut (.I0(r_Clock_Count_adj_5943[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5833));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i13_2_lut (.I0(r_Clock_Count_adj_5943[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5835));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i11_2_lut (.I0(r_Clock_Count_adj_5943[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5834));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i11_2_lut.LUT_INIT = 16'h6666;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 LessThan_1181_i4_4_lut (.I0(r_Clock_Count_adj_5943[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5943[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5830));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50913_3_lut (.I0(n4_adj_5830), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5834), 
            .I3(GND_net), .O(n70408));   // verilog/uart_tx.v(117[17:57])
    defparam i50913_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i13871_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n59772), .I3(GND_net), .O(n32062));   // verilog/coms.v(130[12] 305[6])
    defparam i13871_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i50914_3_lut (.I0(n70408), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5835), 
            .I3(GND_net), .O(n70409));   // verilog/uart_tx.v(117[17:57])
    defparam i50914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49388_4_lut (.I0(n13_adj_5835), .I1(n11_adj_5834), .I2(n9_adj_5833), 
            .I3(n67874), .O(n68883));
    defparam i49388_4_lut.LUT_INIT = 16'heeef;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 LessThan_1181_i8_3_lut (.I0(n6_adj_5831), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5833), .I3(GND_net), .O(n8_adj_5832));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i50693_3_lut (.I0(n70409), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5837), 
            .I3(GND_net), .O(n14_adj_5836));   // verilog/uart_tx.v(117[17:57])
    defparam i50693_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i50335_4_lut (.I0(n14_adj_5836), .I1(n8_adj_5832), .I2(n15_adj_5837), 
            .I3(n68883), .O(n69830));   // verilog/uart_tx.v(117[17:57])
    defparam i50335_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50336_3_lut (.I0(n69830), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5943[8]), 
            .I3(GND_net), .O(n5233));   // verilog/uart_tx.v(117[17:57])
    defparam i50336_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i1_3_lut_adj_1803 (.I0(o_Rx_DV_N_3488[12]), .I1(n5233), .I2(n59789), 
            .I3(GND_net), .O(n63273));
    defparam i1_3_lut_adj_1803.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63273), .O(n63279));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i13874_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n59772), .I3(GND_net), .O(n32065));   // verilog/coms.v(130[12] 305[6])
    defparam i13874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49452_3_lut (.I0(n70311), .I1(current_limit[10]), .I2(n21_adj_5756), 
            .I3(GND_net), .O(n68947));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i49452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13877_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n59772), .I3(GND_net), .O(n32068));   // verilog/coms.v(130[12] 305[6])
    defparam i13877_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 i4_4_lut_adj_1805 (.I0(n55748), .I1(\data_out_frame[16] [4]), 
            .I2(n60150), .I3(n6_adj_5861), .O(n55746));
    defparam i4_4_lut_adj_1805.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1806 (.I0(\data_out_frame[17] [6]), .I1(n60523), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_1806.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1807 (.I0(\data_out_frame[18] [0]), .I1(n55760), 
            .I2(n28460), .I3(n6), .O(n55737));
    defparam i4_4_lut_adj_1807.LUT_INIT = 16'h9669;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n52714), .O(n1240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9946_bdd_4_lut_52112 (.I0(n9946), .I1(current[15]), .I2(duty[22]), 
            .I3(n9944), .O(n71397));
    defparam n9946_bdd_4_lut_52112.LUT_INIT = 16'he4aa;
    SB_LUT4 n71397_bdd_4_lut (.I0(n71397), .I1(duty[19]), .I2(n4924), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[19]));
    defparam n71397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50620_4_lut (.I0(n68947), .I1(n14_adj_5760), .I2(n21_adj_5756), 
            .I3(n69468), .O(n70115));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50620_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50621_3_lut (.I0(n70115), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5755));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50621_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n9946_bdd_4_lut_51865 (.I0(n9946), .I1(current[15]), .I2(duty[21]), 
            .I3(n9944), .O(n71391));
    defparam n9946_bdd_4_lut_51865.LUT_INIT = 16'he4aa;
    SB_CARRY add_151_13 (.CI(n52714), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n52715));
    SB_CARRY add_151_5 (.CI(n52706), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n52707));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n52734), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n52733), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_32 (.CI(n52733), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n52734));
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n52713), .O(n1241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71391_bdd_4_lut (.I0(n71391), .I1(duty[18]), .I2(n4925), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[18]));
    defparam n71391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder1_position_31__I_0_add_2126_32_lut (.I0(encoder1_position[31]), 
            .I1(n11868), .I2(GND_net), .I3(n54060), .O(encoder1_position_scaled_23__N_43[31])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder1_position_31__I_0_add_2126_31_lut (.I0(GND_net), .I1(n11869), 
            .I2(encoder1_position[30]), .I3(n54059), .O(encoder1_position_scaled_23__N_43[30])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_31 (.CI(n54059), .I0(n11869), 
            .I1(encoder1_position[30]), .CO(n54060));
    SB_LUT4 i1_4_lut_adj_1808 (.I0(current_limit[13]), .I1(n24_adj_5755), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n61810));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder1_position_31__I_0_add_2126_30_lut (.I0(GND_net), .I1(n11870), 
            .I2(encoder1_position[29]), .I3(n54058), .O(encoder1_position_scaled_23__N_43[29])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_30 (.CI(n54058), .I0(n11870), 
            .I1(encoder1_position[29]), .CO(n54059));
    SB_LUT4 encoder1_position_31__I_0_add_2126_29_lut (.I0(GND_net), .I1(n11871), 
            .I2(encoder1_position[28]), .I3(n54057), .O(encoder1_position_scaled_23__N_43[28])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_29 (.CI(n54057), .I0(n11871), 
            .I1(encoder1_position[28]), .CO(n54058));
    SB_LUT4 encoder1_position_31__I_0_add_2126_28_lut (.I0(GND_net), .I1(n11872), 
            .I2(encoder1_position[27]), .I3(n54056), .O(encoder1_position_scaled_23__N_43[27])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_28 (.CI(n54056), .I0(n11872), 
            .I1(encoder1_position[27]), .CO(n54057));
    SB_LUT4 encoder1_position_31__I_0_add_2126_27_lut (.I0(GND_net), .I1(n11873), 
            .I2(encoder1_position[26]), .I3(n54055), .O(encoder1_position_scaled_23__N_43[26])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_27 (.CI(n54055), .I0(n11873), 
            .I1(encoder1_position[26]), .CO(n54056));
    SB_LUT4 encoder1_position_31__I_0_add_2126_26_lut (.I0(GND_net), .I1(n11874), 
            .I2(encoder1_position[25]), .I3(n54054), .O(encoder1_position_scaled_23__N_43[25])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_26 (.CI(n54054), .I0(n11874), 
            .I1(encoder1_position[25]), .CO(n54055));
    SB_LUT4 encoder1_position_31__I_0_add_2126_25_lut (.I0(GND_net), .I1(n11875), 
            .I2(encoder1_position[24]), .I3(n54053), .O(encoder1_position_scaled_23__N_43[24])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_25 (.CI(n54053), .I0(n11875), 
            .I1(encoder1_position[24]), .CO(n54054));
    SB_LUT4 encoder1_position_31__I_0_add_2126_24_lut (.I0(GND_net), .I1(n11876), 
            .I2(encoder1_position[23]), .I3(n54052), .O(encoder1_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_24 (.CI(n54052), .I0(n11876), 
            .I1(encoder1_position[23]), .CO(n54053));
    SB_LUT4 encoder1_position_31__I_0_add_2126_23_lut (.I0(GND_net), .I1(n11877), 
            .I2(encoder1_position[22]), .I3(n54051), .O(encoder1_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_23 (.CI(n54051), .I0(n11877), 
            .I1(encoder1_position[22]), .CO(n54052));
    SB_LUT4 encoder1_position_31__I_0_add_2126_22_lut (.I0(GND_net), .I1(n11878), 
            .I2(encoder1_position[21]), .I3(n54050), .O(encoder1_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_22 (.CI(n54050), .I0(n11878), 
            .I1(encoder1_position[21]), .CO(n54051));
    SB_LUT4 encoder1_position_31__I_0_add_2126_21_lut (.I0(GND_net), .I1(n11879), 
            .I2(encoder1_position[20]), .I3(n54049), .O(encoder1_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_21 (.CI(n54049), .I0(n11879), 
            .I1(encoder1_position[20]), .CO(n54050));
    SB_LUT4 encoder1_position_31__I_0_add_2126_20_lut (.I0(GND_net), .I1(n11880), 
            .I2(encoder1_position[19]), .I3(n54048), .O(encoder1_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_20 (.CI(n54048), .I0(n11880), 
            .I1(encoder1_position[19]), .CO(n54049));
    SB_LUT4 encoder1_position_31__I_0_add_2126_19_lut (.I0(GND_net), .I1(n11881), 
            .I2(encoder1_position[18]), .I3(n54047), .O(encoder1_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_19 (.CI(n54047), .I0(n11881), 
            .I1(encoder1_position[18]), .CO(n54048));
    SB_LUT4 encoder1_position_31__I_0_add_2126_18_lut (.I0(GND_net), .I1(n11882), 
            .I2(encoder1_position[17]), .I3(n54046), .O(encoder1_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_18 (.CI(n54046), .I0(n11882), 
            .I1(encoder1_position[17]), .CO(n54047));
    SB_LUT4 encoder1_position_31__I_0_add_2126_17_lut (.I0(GND_net), .I1(n11883), 
            .I2(encoder1_position[16]), .I3(n54045), .O(encoder1_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(current_limit[13]), .I1(n24_adj_5755), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n61815));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'h8000;
    SB_CARRY encoder1_position_31__I_0_add_2126_17 (.CI(n54045), .I0(n11883), 
            .I1(encoder1_position[16]), .CO(n54046));
    SB_LUT4 encoder1_position_31__I_0_add_2126_16_lut (.I0(GND_net), .I1(n11884), 
            .I2(encoder1_position[15]), .I3(n54044), .O(encoder1_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6927_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n24006));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i6927_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY encoder1_position_31__I_0_add_2126_16 (.CI(n54044), .I0(n11884), 
            .I1(encoder1_position[15]), .CO(n54045));
    SB_LUT4 encoder1_position_31__I_0_add_2126_15_lut (.I0(GND_net), .I1(n11885), 
            .I2(encoder1_position[14]), .I3(n54043), .O(encoder1_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6186_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i6186_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY encoder1_position_31__I_0_add_2126_15 (.CI(n54043), .I0(n11885), 
            .I1(encoder1_position[14]), .CO(n54044));
    SB_LUT4 i13918_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n24006), .I3(n4_adj_5867), .O(n32109));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i13918_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 encoder1_position_31__I_0_add_2126_14_lut (.I0(GND_net), .I1(n11886), 
            .I2(encoder1_position[13]), .I3(n54042), .O(encoder1_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5230), .I3(o_Rx_DV_N_3488[8]), .O(n63069));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63069), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_1178_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5841));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1178_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5838));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1178_i8_3_lut (.I0(n6_adj_5839), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5841), .I3(GND_net), .O(n8_adj_5840));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51244_4_lut (.I0(n8_adj_5840), .I1(n4_adj_5838), .I2(n9_adj_5841), 
            .I3(n67858), .O(n70739));   // verilog/uart_rx.v(119[17:57])
    defparam i51244_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51245_3_lut (.I0(n70739), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n70740));   // verilog/uart_rx.v(119[17:57])
    defparam i51245_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51144_3_lut (.I0(n70740), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n70639));   // verilog/uart_rx.v(119[17:57])
    defparam i51144_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51000_3_lut (.I0(n70639), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5230));   // verilog/uart_rx.v(119[17:57])
    defparam i51000_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n59798), .O(n63263));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1813 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63263), .O(n63269));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 n9946_bdd_4_lut_51860 (.I0(n9946), .I1(current[6]), .I2(duty[9]), 
            .I3(n9944), .O(n71385));
    defparam n9946_bdd_4_lut_51860.LUT_INIT = 16'he4aa;
    SB_CARRY encoder1_position_31__I_0_add_2126_14 (.CI(n54042), .I0(n11886), 
            .I1(encoder1_position[13]), .CO(n54043));
    SB_LUT4 encoder1_position_31__I_0_add_2126_13_lut (.I0(GND_net), .I1(n11887), 
            .I2(encoder1_position[12]), .I3(n54041), .O(encoder1_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_13 (.CI(n54041), .I0(n11887), 
            .I1(encoder1_position[12]), .CO(n54042));
    SB_LUT4 encoder1_position_31__I_0_add_2126_12_lut (.I0(GND_net), .I1(n11888), 
            .I2(encoder1_position[11]), .I3(n54040), .O(encoder1_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_12 (.CI(n54040), .I0(n11888), 
            .I1(encoder1_position[11]), .CO(n54041));
    SB_LUT4 encoder1_position_31__I_0_add_2126_11_lut (.I0(GND_net), .I1(n11889), 
            .I2(encoder1_position[10]), .I3(n54039), .O(encoder1_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_11 (.CI(n54039), .I0(n11889), 
            .I1(encoder1_position[10]), .CO(n54040));
    SB_LUT4 encoder1_position_31__I_0_add_2126_10_lut (.I0(GND_net), .I1(n11890), 
            .I2(encoder1_position[9]), .I3(n54038), .O(encoder1_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_10 (.CI(n54038), .I0(n11890), 
            .I1(encoder1_position[9]), .CO(n54039));
    SB_LUT4 encoder1_position_31__I_0_add_2126_9_lut (.I0(GND_net), .I1(n11891), 
            .I2(encoder1_position[8]), .I3(n54037), .O(encoder1_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_31__I_0_add_2126_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_31__I_0_add_2126_9 (.CI(n54037), .I0(n11891), 
            .I1(encoder1_position[8]), .CO(n54038));
    SB_CARRY encoder1_position_31__I_0_add_2126_8 (.CI(n54036), .I0(n11892), 
            .I1(encoder1_position[7]), .CO(n54037));
    SB_CARRY encoder1_position_31__I_0_add_2126_7 (.CI(n54035), .I0(n11893), 
            .I1(encoder1_position[6]), .CO(n54036));
    SB_CARRY encoder1_position_31__I_0_add_2126_6 (.CI(n54034), .I0(n11894), 
            .I1(encoder1_position[5]), .CO(n54035));
    SB_CARRY encoder1_position_31__I_0_add_2126_5 (.CI(n54033), .I0(n11895), 
            .I1(encoder1_position[4]), .CO(n54034));
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder1_position_31__I_0_add_2126_4 (.CI(n54032), .I0(n11896), 
            .I1(encoder1_position[3]), .CO(n54033));
    SB_CARRY encoder1_position_31__I_0_add_2126_3 (.CI(n54031), .I0(n11897), 
            .I1(encoder1_position[2]), .CO(n54032));
    SB_CARRY encoder1_position_31__I_0_add_2126_2 (.CI(GND_net), .I0(encoder1_position[0]), 
            .I1(encoder1_position[1]), .CO(n54031));
    SB_LUT4 add_4929_31_lut (.I0(GND_net), .I1(n13511), .I2(encoder1_position[30]), 
            .I3(n54030), .O(n11868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_30_lut (.I0(GND_net), .I1(n13512), .I2(encoder1_position[29]), 
            .I3(n54029), .O(n11869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_30 (.CI(n54029), .I0(n13512), .I1(encoder1_position[29]), 
            .CO(n54030));
    SB_LUT4 add_4929_29_lut (.I0(GND_net), .I1(n13513), .I2(encoder1_position[28]), 
            .I3(n54028), .O(n11870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_29 (.CI(n54028), .I0(n13513), .I1(encoder1_position[28]), 
            .CO(n54029));
    SB_LUT4 add_4929_28_lut (.I0(GND_net), .I1(n13514), .I2(encoder1_position[27]), 
            .I3(n54027), .O(n11871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_28_lut.LUT_INIT = 16'hC33C;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32109));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_4929_28 (.CI(n54027), .I0(n13514), .I1(encoder1_position[27]), 
            .CO(n54028));
    SB_LUT4 i13611_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n30673), 
            .I3(GND_net), .O(n31802));   // verilog/coms.v(130[12] 305[6])
    defparam i13611_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_4929_27_lut (.I0(GND_net), .I1(n13515), .I2(encoder1_position[26]), 
            .I3(n54026), .O(n11872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_27 (.CI(n54026), .I0(n13515), .I1(encoder1_position[26]), 
            .CO(n54027));
    SB_LUT4 add_4929_26_lut (.I0(GND_net), .I1(n13516), .I2(encoder1_position[25]), 
            .I3(n54025), .O(n11873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_26 (.CI(n54025), .I0(n13516), .I1(encoder1_position[25]), 
            .CO(n54026));
    SB_LUT4 add_4929_25_lut (.I0(GND_net), .I1(n13517), .I2(encoder1_position[24]), 
            .I3(n54024), .O(n11874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_25 (.CI(n54024), .I0(n13517), .I1(encoder1_position[24]), 
            .CO(n54025));
    SB_LUT4 add_4929_24_lut (.I0(GND_net), .I1(n13518), .I2(encoder1_position[23]), 
            .I3(n54023), .O(n11875)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_24 (.CI(n54023), .I0(n13518), .I1(encoder1_position[23]), 
            .CO(n54024));
    SB_LUT4 add_4929_23_lut (.I0(GND_net), .I1(n13519), .I2(encoder1_position[22]), 
            .I3(n54022), .O(n11876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_23 (.CI(n54022), .I0(n13519), .I1(encoder1_position[22]), 
            .CO(n54023));
    SB_LUT4 add_4929_22_lut (.I0(GND_net), .I1(n13520), .I2(encoder1_position[21]), 
            .I3(n54021), .O(n11877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_22 (.CI(n54021), .I0(n13520), .I1(encoder1_position[21]), 
            .CO(n54022));
    SB_LUT4 add_4929_21_lut (.I0(GND_net), .I1(n13521), .I2(encoder1_position[20]), 
            .I3(n54020), .O(n11878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_21 (.CI(n54020), .I0(n13521), .I1(encoder1_position[20]), 
            .CO(n54021));
    SB_LUT4 add_4929_20_lut (.I0(GND_net), .I1(n13522), .I2(encoder1_position[19]), 
            .I3(n54019), .O(n11879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_20 (.CI(n54019), .I0(n13522), .I1(encoder1_position[19]), 
            .CO(n54020));
    SB_LUT4 add_4929_19_lut (.I0(GND_net), .I1(n13523), .I2(encoder1_position[18]), 
            .I3(n54018), .O(n11880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_19 (.CI(n54018), .I0(n13523), .I1(encoder1_position[18]), 
            .CO(n54019));
    SB_LUT4 add_4929_18_lut (.I0(GND_net), .I1(n13524), .I2(encoder1_position[17]), 
            .I3(n54017), .O(n11881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n61815), .I3(n61810), .O(n260));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hb3a2;
    SB_CARRY add_4929_18 (.CI(n54017), .I0(n13524), .I1(encoder1_position[17]), 
            .CO(n54018));
    SB_LUT4 add_4929_17_lut (.I0(GND_net), .I1(n13525), .I2(encoder1_position[16]), 
            .I3(n54016), .O(n11882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_17 (.CI(n54016), .I0(n13525), .I1(encoder1_position[16]), 
            .CO(n54017));
    SB_LUT4 add_4929_16_lut (.I0(GND_net), .I1(n13526), .I2(encoder1_position[15]), 
            .I3(n54015), .O(n11883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_16 (.CI(n54015), .I0(n13526), .I1(encoder1_position[15]), 
            .CO(n54016));
    SB_LUT4 add_4929_15_lut (.I0(GND_net), .I1(n13527), .I2(encoder1_position[14]), 
            .I3(n54014), .O(n11884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_15 (.CI(n54014), .I0(n13527), .I1(encoder1_position[14]), 
            .CO(n54015));
    SB_LUT4 add_4929_14_lut (.I0(GND_net), .I1(n13528), .I2(encoder1_position[13]), 
            .I3(n54013), .O(n11885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_14 (.CI(n54013), .I0(n13528), .I1(encoder1_position[13]), 
            .CO(n54014));
    SB_LUT4 add_4929_13_lut (.I0(GND_net), .I1(n13529), .I2(encoder1_position[12]), 
            .I3(n54012), .O(n11886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_13 (.CI(n54012), .I0(n13529), .I1(encoder1_position[12]), 
            .CO(n54013));
    SB_LUT4 add_4929_12_lut (.I0(GND_net), .I1(n13530), .I2(encoder1_position[11]), 
            .I3(n54011), .O(n11887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_12 (.CI(n54011), .I0(n13530), .I1(encoder1_position[11]), 
            .CO(n54012));
    SB_LUT4 add_4929_11_lut (.I0(GND_net), .I1(n13531), .I2(encoder1_position[10]), 
            .I3(n54010), .O(n11888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_11 (.CI(n54010), .I0(n13531), .I1(encoder1_position[10]), 
            .CO(n54011));
    SB_LUT4 add_4929_10_lut (.I0(GND_net), .I1(n13532), .I2(encoder1_position[9]), 
            .I3(n54009), .O(n11889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_10 (.CI(n54009), .I0(n13532), .I1(encoder1_position[9]), 
            .CO(n54010));
    SB_LUT4 add_4929_9_lut (.I0(GND_net), .I1(n13533), .I2(encoder1_position[8]), 
            .I3(n54008), .O(n11890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_9 (.CI(n54008), .I0(n13533), .I1(encoder1_position[8]), 
            .CO(n54009));
    SB_LUT4 add_4929_8_lut (.I0(GND_net), .I1(n13534), .I2(encoder1_position[7]), 
            .I3(n54007), .O(n11891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_8 (.CI(n54007), .I0(n13534), .I1(encoder1_position[7]), 
            .CO(n54008));
    SB_LUT4 add_4929_7_lut (.I0(GND_net), .I1(n13535), .I2(encoder1_position[6]), 
            .I3(n54006), .O(n11892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_7 (.CI(n54006), .I0(n13535), .I1(encoder1_position[6]), 
            .CO(n54007));
    SB_LUT4 add_4929_6_lut (.I0(GND_net), .I1(n13536), .I2(encoder1_position[5]), 
            .I3(n54005), .O(n11893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_6 (.CI(n54005), .I0(n13536), .I1(encoder1_position[5]), 
            .CO(n54006));
    SB_LUT4 add_4929_5_lut (.I0(GND_net), .I1(n13537), .I2(encoder1_position[4]), 
            .I3(n54004), .O(n11894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_5 (.CI(n54004), .I0(n13537), .I1(encoder1_position[4]), 
            .CO(n54005));
    SB_LUT4 add_4929_4_lut (.I0(GND_net), .I1(n13538), .I2(encoder1_position[3]), 
            .I3(n54003), .O(n11895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_4 (.CI(n54003), .I0(n13538), .I1(encoder1_position[3]), 
            .CO(n54004));
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52063 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[0]), .O(n71577));
    defparam byte_transmit_counter_1__bdd_4_lut_52063.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4929_3_lut (.I0(GND_net), .I1(n13539), .I2(encoder1_position[2]), 
            .I3(n54002), .O(n11896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_3 (.CI(n54002), .I0(n13539), .I1(encoder1_position[2]), 
            .CO(n54003));
    SB_LUT4 add_4929_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n11897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n52705), .O(n1249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71577_bdd_4_lut (.I0(n71577), .I1(\data_out_frame[26] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[0]), 
            .O(n71580));
    defparam n71577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4929_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n54002));
    SB_LUT4 add_4996_30_lut (.I0(GND_net), .I1(n14994), .I2(encoder1_position[29]), 
            .I3(n54001), .O(n13511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4996_29_lut (.I0(GND_net), .I1(n14995), .I2(encoder1_position[28]), 
            .I3(n54000), .O(n13512)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_29 (.CI(n54000), .I0(n14995), .I1(encoder1_position[28]), 
            .CO(n54001));
    SB_LUT4 add_4996_28_lut (.I0(GND_net), .I1(n14996), .I2(encoder1_position[27]), 
            .I3(n53999), .O(n13513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_28 (.CI(n53999), .I0(n14996), .I1(encoder1_position[27]), 
            .CO(n54000));
    SB_LUT4 add_4996_27_lut (.I0(GND_net), .I1(n14997), .I2(encoder1_position[26]), 
            .I3(n53998), .O(n13514)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_27 (.CI(n53998), .I0(n14997), .I1(encoder1_position[26]), 
            .CO(n53999));
    SB_LUT4 add_4996_26_lut (.I0(GND_net), .I1(n14998), .I2(encoder1_position[25]), 
            .I3(n53997), .O(n13515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_26 (.CI(n53997), .I0(n14998), .I1(encoder1_position[25]), 
            .CO(n53998));
    SB_LUT4 add_4996_25_lut (.I0(GND_net), .I1(n14999), .I2(encoder1_position[24]), 
            .I3(n53996), .O(n13516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_25 (.CI(n53996), .I0(n14999), .I1(encoder1_position[24]), 
            .CO(n53997));
    SB_LUT4 add_4996_24_lut (.I0(GND_net), .I1(n15000), .I2(encoder1_position[23]), 
            .I3(n53995), .O(n13517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_24 (.CI(n53995), .I0(n15000), .I1(encoder1_position[23]), 
            .CO(n53996));
    SB_LUT4 add_4996_23_lut (.I0(GND_net), .I1(n15001), .I2(encoder1_position[22]), 
            .I3(n53994), .O(n13518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_23 (.CI(n53994), .I0(n15001), .I1(encoder1_position[22]), 
            .CO(n53995));
    SB_LUT4 add_4996_22_lut (.I0(GND_net), .I1(n15002), .I2(encoder1_position[21]), 
            .I3(n53993), .O(n13519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_22 (.CI(n53993), .I0(n15002), .I1(encoder1_position[21]), 
            .CO(n53994));
    SB_LUT4 add_4996_21_lut (.I0(GND_net), .I1(n15003), .I2(encoder1_position[20]), 
            .I3(n53992), .O(n13520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_21 (.CI(n53992), .I0(n15003), .I1(encoder1_position[20]), 
            .CO(n53993));
    SB_CARRY add_151_12 (.CI(n52713), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n52714));
    SB_LUT4 add_4996_20_lut (.I0(GND_net), .I1(n15004), .I2(encoder1_position[19]), 
            .I3(n53991), .O(n13521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_20 (.CI(n53991), .I0(n15004), .I1(encoder1_position[19]), 
            .CO(n53992));
    SB_LUT4 add_4996_19_lut (.I0(GND_net), .I1(n15005), .I2(encoder1_position[18]), 
            .I3(n53990), .O(n13522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_19 (.CI(n53990), .I0(n15005), .I1(encoder1_position[18]), 
            .CO(n53991));
    SB_LUT4 add_4996_18_lut (.I0(GND_net), .I1(n15006), .I2(encoder1_position[17]), 
            .I3(n53989), .O(n13523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_18 (.CI(n53989), .I0(n15006), .I1(encoder1_position[17]), 
            .CO(n53990));
    SB_LUT4 add_4996_17_lut (.I0(GND_net), .I1(n15007), .I2(encoder1_position[16]), 
            .I3(n53988), .O(n13524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_17 (.CI(n53988), .I0(n15007), .I1(encoder1_position[16]), 
            .CO(n53989));
    SB_LUT4 add_4996_16_lut (.I0(GND_net), .I1(n15008), .I2(encoder1_position[15]), 
            .I3(n53987), .O(n13525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_16 (.CI(n53987), .I0(n15008), .I1(encoder1_position[15]), 
            .CO(n53988));
    SB_LUT4 add_4996_15_lut (.I0(GND_net), .I1(n15009), .I2(encoder1_position[14]), 
            .I3(n53986), .O(n13526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_15 (.CI(n53986), .I0(n15009), .I1(encoder1_position[14]), 
            .CO(n53987));
    SB_LUT4 add_4996_14_lut (.I0(GND_net), .I1(n15010), .I2(encoder1_position[13]), 
            .I3(n53985), .O(n13527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_14 (.CI(n53985), .I0(n15010), .I1(encoder1_position[13]), 
            .CO(n53986));
    SB_LUT4 add_4996_13_lut (.I0(GND_net), .I1(n15011), .I2(encoder1_position[12]), 
            .I3(n53984), .O(n13528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_13 (.CI(n53984), .I0(n15011), .I1(encoder1_position[12]), 
            .CO(n53985));
    SB_LUT4 add_4996_12_lut (.I0(GND_net), .I1(n15012), .I2(encoder1_position[11]), 
            .I3(n53983), .O(n13529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_12 (.CI(n53983), .I0(n15012), .I1(encoder1_position[11]), 
            .CO(n53984));
    SB_LUT4 add_4996_11_lut (.I0(GND_net), .I1(n15013), .I2(encoder1_position[10]), 
            .I3(n53982), .O(n13530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_11 (.CI(n53982), .I0(n15013), .I1(encoder1_position[10]), 
            .CO(n53983));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n52732), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4996_10_lut (.I0(GND_net), .I1(n15014), .I2(encoder1_position[9]), 
            .I3(n53981), .O(n13531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_10 (.CI(n53981), .I0(n15014), .I1(encoder1_position[9]), 
            .CO(n53982));
    SB_LUT4 add_4996_9_lut (.I0(GND_net), .I1(n15015), .I2(encoder1_position[8]), 
            .I3(n53980), .O(n13532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_9 (.CI(n53980), .I0(n15015), .I1(encoder1_position[8]), 
            .CO(n53981));
    SB_LUT4 add_4996_8_lut (.I0(GND_net), .I1(n15016), .I2(encoder1_position[7]), 
            .I3(n53979), .O(n13533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_8 (.CI(n53979), .I0(n15016), .I1(encoder1_position[7]), 
            .CO(n53980));
    SB_LUT4 add_4996_7_lut (.I0(GND_net), .I1(n15017), .I2(encoder1_position[6]), 
            .I3(n53978), .O(n13534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5763));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4996_7 (.CI(n53978), .I0(n15017), .I1(encoder1_position[6]), 
            .CO(n53979));
    SB_LUT4 add_4996_6_lut (.I0(GND_net), .I1(n15018), .I2(encoder1_position[5]), 
            .I3(n53977), .O(n13535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_6 (.CI(n53977), .I0(n15018), .I1(encoder1_position[5]), 
            .CO(n53978));
    SB_LUT4 add_4996_5_lut (.I0(GND_net), .I1(n15019), .I2(encoder1_position[4]), 
            .I3(n53976), .O(n13536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_5 (.CI(n53976), .I0(n15019), .I1(encoder1_position[4]), 
            .CO(n53977));
    SB_LUT4 add_4996_4_lut (.I0(GND_net), .I1(n15020), .I2(encoder1_position[3]), 
            .I3(n53975), .O(n13537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_4 (.CI(n53975), .I0(n15020), .I1(encoder1_position[3]), 
            .CO(n53976));
    SB_LUT4 add_4996_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n53974), .O(n13538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_3 (.CI(n53974), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n53975));
    SB_LUT4 add_4996_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n13539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4996_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4996_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n53974));
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5767));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5766));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5765));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5172_28_lut (.I0(GND_net), .I1(n17512), .I2(encoder1_position[28]), 
            .I3(n53967), .O(n14994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5172_27_lut (.I0(GND_net), .I1(n17513), .I2(encoder1_position[27]), 
            .I3(n53966), .O(n14995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_27 (.CI(n53966), .I0(n17513), .I1(encoder1_position[27]), 
            .CO(n53967));
    SB_LUT4 add_5172_26_lut (.I0(GND_net), .I1(n17514), .I2(encoder1_position[26]), 
            .I3(n53965), .O(n14996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_26 (.CI(n53965), .I0(n17514), .I1(encoder1_position[26]), 
            .CO(n53966));
    SB_LUT4 add_5172_25_lut (.I0(GND_net), .I1(n17515), .I2(encoder1_position[25]), 
            .I3(n53964), .O(n14997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_25 (.CI(n53964), .I0(n17515), .I1(encoder1_position[25]), 
            .CO(n53965));
    SB_LUT4 add_5172_24_lut (.I0(GND_net), .I1(n17516), .I2(encoder1_position[24]), 
            .I3(n53963), .O(n14998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_24 (.CI(n53963), .I0(n17516), .I1(encoder1_position[24]), 
            .CO(n53964));
    SB_LUT4 add_5172_23_lut (.I0(GND_net), .I1(n17517), .I2(encoder1_position[23]), 
            .I3(n53962), .O(n14999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_23 (.CI(n53962), .I0(n17517), .I1(encoder1_position[23]), 
            .CO(n53963));
    SB_LUT4 add_5172_22_lut (.I0(GND_net), .I1(n17518), .I2(encoder1_position[22]), 
            .I3(n53961), .O(n15000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_22 (.CI(n53961), .I0(n17518), .I1(encoder1_position[22]), 
            .CO(n53962));
    SB_LUT4 add_5172_21_lut (.I0(GND_net), .I1(n17519), .I2(encoder1_position[21]), 
            .I3(n53960), .O(n15001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_21 (.CI(n53960), .I0(n17519), .I1(encoder1_position[21]), 
            .CO(n53961));
    SB_LUT4 add_5172_20_lut (.I0(GND_net), .I1(n17520), .I2(encoder1_position[20]), 
            .I3(n53959), .O(n15002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_20 (.CI(n53959), .I0(n17520), .I1(encoder1_position[20]), 
            .CO(n53960));
    SB_LUT4 add_5172_19_lut (.I0(GND_net), .I1(n17521), .I2(encoder1_position[19]), 
            .I3(n53958), .O(n15003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_19 (.CI(n53958), .I0(n17521), .I1(encoder1_position[19]), 
            .CO(n53959));
    SB_LUT4 add_5172_18_lut (.I0(GND_net), .I1(n17522), .I2(encoder1_position[18]), 
            .I3(n53957), .O(n15004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_18 (.CI(n53957), .I0(n17522), .I1(encoder1_position[18]), 
            .CO(n53958));
    SB_LUT4 add_5172_17_lut (.I0(GND_net), .I1(n17523), .I2(encoder1_position[17]), 
            .I3(n53956), .O(n15005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_17 (.CI(n53956), .I0(n17523), .I1(encoder1_position[17]), 
            .CO(n53957));
    SB_LUT4 add_5172_16_lut (.I0(GND_net), .I1(n17524), .I2(encoder1_position[16]), 
            .I3(n53955), .O(n15006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_16 (.CI(n53955), .I0(n17524), .I1(encoder1_position[16]), 
            .CO(n53956));
    SB_LUT4 add_5172_15_lut (.I0(GND_net), .I1(n17525), .I2(encoder1_position[15]), 
            .I3(n53954), .O(n15007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_15 (.CI(n53954), .I0(n17525), .I1(encoder1_position[15]), 
            .CO(n53955));
    SB_LUT4 add_5172_14_lut (.I0(GND_net), .I1(n17526), .I2(encoder1_position[14]), 
            .I3(n53953), .O(n15008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5771));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5770));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5172_14 (.CI(n53953), .I0(n17526), .I1(encoder1_position[14]), 
            .CO(n53954));
    SB_LUT4 add_5172_13_lut (.I0(GND_net), .I1(n17527), .I2(encoder1_position[13]), 
            .I3(n53952), .O(n15009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_13 (.CI(n53952), .I0(n17527), .I1(encoder1_position[13]), 
            .CO(n53953));
    SB_LUT4 add_5172_12_lut (.I0(GND_net), .I1(n17528), .I2(encoder1_position[12]), 
            .I3(n53951), .O(n15010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_12 (.CI(n53951), .I0(n17528), .I1(encoder1_position[12]), 
            .CO(n53952));
    SB_LUT4 add_5172_11_lut (.I0(GND_net), .I1(n17529), .I2(encoder1_position[11]), 
            .I3(n53950), .O(n15011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_11 (.CI(n53950), .I0(n17529), .I1(encoder1_position[11]), 
            .CO(n53951));
    SB_LUT4 add_5172_10_lut (.I0(GND_net), .I1(n17530), .I2(encoder1_position[10]), 
            .I3(n53949), .O(n15012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_10 (.CI(n53949), .I0(n17530), .I1(encoder1_position[10]), 
            .CO(n53950));
    SB_LUT4 add_5172_9_lut (.I0(GND_net), .I1(n17531), .I2(encoder1_position[9]), 
            .I3(n53948), .O(n15013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_9 (.CI(n53948), .I0(n17531), .I1(encoder1_position[9]), 
            .CO(n53949));
    SB_LUT4 dti_counter_2038_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n53495), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5172_8_lut (.I0(GND_net), .I1(n17532), .I2(encoder1_position[8]), 
            .I3(n53947), .O(n15014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n53494), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_8 (.CI(n53947), .I0(n17532), .I1(encoder1_position[8]), 
            .CO(n53948));
    SB_CARRY dti_counter_2038_add_4_8 (.CI(n53494), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n53495));
    SB_LUT4 dti_counter_2038_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n53493), .O(n40_adj_5842)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5172_7_lut (.I0(GND_net), .I1(n17533), .I2(encoder1_position[7]), 
            .I3(n53946), .O(n15015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_7 (.CI(n53946), .I0(n17533), .I1(encoder1_position[7]), 
            .CO(n53947));
    SB_CARRY dti_counter_2038_add_4_7 (.CI(n53493), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n53494));
    SB_LUT4 dti_counter_2038_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n53492), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5172_6_lut (.I0(GND_net), .I1(n17534), .I2(encoder1_position[6]), 
            .I3(n53945), .O(n15016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_6 (.CI(n53945), .I0(n17534), .I1(encoder1_position[6]), 
            .CO(n53946));
    SB_CARRY dti_counter_2038_add_4_6 (.CI(n53492), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n53493));
    SB_LUT4 dti_counter_2038_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n53491), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5172_5_lut (.I0(GND_net), .I1(n17535), .I2(encoder1_position[5]), 
            .I3(n53944), .O(n15017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_5 (.CI(n53944), .I0(n17535), .I1(encoder1_position[5]), 
            .CO(n53945));
    SB_CARRY dti_counter_2038_add_4_5 (.CI(n53491), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n53492));
    SB_LUT4 dti_counter_2038_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n53490), .O(n43_adj_5843)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5769));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5172_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[4]), 
            .I3(n53943), .O(n15018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_4 (.CI(n53943), .I0(encoder1_position[2]), .I1(encoder1_position[4]), 
            .CO(n53944));
    SB_LUT4 add_5172_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[3]), 
            .I3(n53942), .O(n15019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5172_3 (.CI(n53942), .I0(encoder1_position[1]), .I1(encoder1_position[3]), 
            .CO(n53943));
    SB_LUT4 add_5172_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n15020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5172_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5854));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_CARRY add_5172_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n53942));
    SB_LUT4 add_5351_25_lut (.I0(GND_net), .I1(n20274), .I2(encoder1_position[26]), 
            .I3(n53941), .O(n17512)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_4 (.CI(n53490), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n53491));
    SB_LUT4 n71385_bdd_4_lut (.I0(n71385), .I1(duty[6]), .I2(n4937), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n71385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5351_24_lut (.I0(GND_net), .I1(n20275), .I2(encoder1_position[25]), 
            .I3(n53940), .O(n17513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_24 (.CI(n53940), .I0(n20275), .I1(encoder1_position[25]), 
            .CO(n53941));
    SB_LUT4 add_5351_23_lut (.I0(GND_net), .I1(n20276), .I2(encoder1_position[24]), 
            .I3(n53939), .O(n17514)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n53489), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_23 (.CI(n53939), .I0(n20276), .I1(encoder1_position[24]), 
            .CO(n53940));
    SB_LUT4 add_5351_22_lut (.I0(GND_net), .I1(n20277), .I2(encoder1_position[23]), 
            .I3(n53938), .O(n17515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_22 (.CI(n53938), .I0(n20277), .I1(encoder1_position[23]), 
            .CO(n53939));
    SB_LUT4 add_5351_21_lut (.I0(GND_net), .I1(n20278), .I2(encoder1_position[22]), 
            .I3(n53937), .O(n17516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9946_bdd_4_lut_51855 (.I0(n9946), .I1(current[15]), .I2(duty[20]), 
            .I3(n9944), .O(n71379));
    defparam n9946_bdd_4_lut_51855.LUT_INIT = 16'he4aa;
    SB_LUT4 n71379_bdd_4_lut (.I0(n71379), .I1(duty[17]), .I2(n4926), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[17]));
    defparam n71379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9946_bdd_4_lut_51850 (.I0(n9946), .I1(current[15]), .I2(duty[19]), 
            .I3(n9944), .O(n71373));
    defparam n9946_bdd_4_lut_51850.LUT_INIT = 16'he4aa;
    SB_LUT4 n71373_bdd_4_lut (.I0(n71373), .I1(duty[16]), .I2(n4927), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[16]));
    defparam n71373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY dti_counter_2038_add_4_3 (.CI(n53489), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n53490));
    SB_CARRY add_5351_21 (.CI(n53937), .I0(n20278), .I1(encoder1_position[22]), 
            .CO(n53938));
    SB_LUT4 dti_counter_2038_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n53489));
    SB_LUT4 add_5351_20_lut (.I0(GND_net), .I1(n20279), .I2(encoder1_position[21]), 
            .I3(n53936), .O(n17517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_20 (.CI(n53936), .I0(n20279), .I1(encoder1_position[21]), 
            .CO(n53937));
    SB_LUT4 add_5351_19_lut (.I0(GND_net), .I1(n20280), .I2(encoder1_position[20]), 
            .I3(n53935), .O(n17518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_19 (.CI(n53935), .I0(n20280), .I1(encoder1_position[20]), 
            .CO(n53936));
    SB_LUT4 add_5351_18_lut (.I0(GND_net), .I1(n20281), .I2(encoder1_position[19]), 
            .I3(n53934), .O(n17519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_18 (.CI(n53934), .I0(n20281), .I1(encoder1_position[19]), 
            .CO(n53935));
    SB_LUT4 add_5351_17_lut (.I0(GND_net), .I1(n20282), .I2(encoder1_position[18]), 
            .I3(n53933), .O(n17520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_17 (.CI(n53933), .I0(n20282), .I1(encoder1_position[18]), 
            .CO(n53934));
    SB_LUT4 add_5351_16_lut (.I0(GND_net), .I1(n20283), .I2(encoder1_position[17]), 
            .I3(n53932), .O(n17521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_16 (.CI(n53932), .I0(n20283), .I1(encoder1_position[17]), 
            .CO(n53933));
    SB_LUT4 add_5351_15_lut (.I0(GND_net), .I1(n20284), .I2(encoder1_position[16]), 
            .I3(n53931), .O(n17522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_15 (.CI(n53931), .I0(n20284), .I1(encoder1_position[16]), 
            .CO(n53932));
    SB_LUT4 add_5351_14_lut (.I0(GND_net), .I1(n20285), .I2(encoder1_position[15]), 
            .I3(n53930), .O(n17523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_14 (.CI(n53930), .I0(n20285), .I1(encoder1_position[15]), 
            .CO(n53931));
    SB_LUT4 add_5351_13_lut (.I0(GND_net), .I1(n20286), .I2(encoder1_position[14]), 
            .I3(n53929), .O(n17524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_13 (.CI(n53929), .I0(n20286), .I1(encoder1_position[14]), 
            .CO(n53930));
    SB_LUT4 add_5351_12_lut (.I0(GND_net), .I1(n20287), .I2(encoder1_position[13]), 
            .I3(n53928), .O(n17525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_12 (.CI(n53928), .I0(n20287), .I1(encoder1_position[13]), 
            .CO(n53929));
    SB_LUT4 add_5351_11_lut (.I0(GND_net), .I1(n20288), .I2(encoder1_position[12]), 
            .I3(n53927), .O(n17526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_11 (.CI(n53927), .I0(n20288), .I1(encoder1_position[12]), 
            .CO(n53928));
    SB_LUT4 add_5351_10_lut (.I0(GND_net), .I1(n20289), .I2(encoder1_position[11]), 
            .I3(n53926), .O(n17527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n52712), .O(n1242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_4 (.CI(n52705), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n52706));
    SB_CARRY add_5351_10 (.CI(n53926), .I0(n20289), .I1(encoder1_position[11]), 
            .CO(n53927));
    SB_LUT4 add_5351_9_lut (.I0(GND_net), .I1(n20290), .I2(encoder1_position[10]), 
            .I3(n53925), .O(n17528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_9 (.CI(n53925), .I0(n20290), .I1(encoder1_position[10]), 
            .CO(n53926));
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5775));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5773));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5351_8_lut (.I0(GND_net), .I1(n20291), .I2(encoder1_position[9]), 
            .I3(n53924), .O(n17529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_8 (.CI(n53924), .I0(n20291), .I1(encoder1_position[9]), 
            .CO(n53925));
    SB_LUT4 add_5351_7_lut (.I0(GND_net), .I1(n20292), .I2(encoder1_position[8]), 
            .I3(n53923), .O(n17530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_7 (.CI(n53923), .I0(n20292), .I1(encoder1_position[8]), 
            .CO(n53924));
    SB_LUT4 add_5351_6_lut (.I0(GND_net), .I1(n20293), .I2(encoder1_position[7]), 
            .I3(n53922), .O(n17531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_6 (.CI(n53922), .I0(n20293), .I1(encoder1_position[7]), 
            .CO(n53923));
    SB_CARRY add_151_31 (.CI(n52732), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n52733));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n52731), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5351_5_lut (.I0(GND_net), .I1(n20294), .I2(encoder1_position[6]), 
            .I3(n53921), .O(n17532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_5 (.CI(n53921), .I0(n20294), .I1(encoder1_position[6]), 
            .CO(n53922));
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_5351_4_lut (.I0(GND_net), .I1(n20295), .I2(encoder1_position[5]), 
            .I3(n53920), .O(n17533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_4_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dti_counter_2038__i0 (.Q(dti_counter[0]), .C(clk16MHz), .D(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_CARRY add_5351_4 (.CI(n53920), .I0(n20295), .I1(encoder1_position[5]), 
            .CO(n53921));
    SB_LUT4 mux_243_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_91[10]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_5351_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[4]), 
            .I3(n53919), .O(n17534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9946_bdd_4_lut_51845 (.I0(n9946), .I1(current[15]), .I2(duty[18]), 
            .I3(n9944), .O(n71367));
    defparam n9946_bdd_4_lut_51845.LUT_INIT = 16'he4aa;
    SB_CARRY add_5351_3 (.CI(n53919), .I0(encoder1_position[1]), .I1(encoder1_position[4]), 
            .CO(n53920));
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n67567), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5351_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[3]), 
            .I3(GND_net), .O(n17535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5351_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5351_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[3]), 
            .CO(n53919));
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 n71367_bdd_4_lut (.I0(n71367), .I1(duty[15]), .I2(n4928), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[15]));
    defparam n71367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50616_3_lut (.I0(n4), .I1(n305), .I2(n11), .I3(GND_net), 
            .O(n70111));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i50616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50617_3_lut (.I0(n70111), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n70112));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i50617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8_adj_5753));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7), .I3(GND_net), 
            .O(n6_adj_5754));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5753), .I1(n301), .I2(n19_adj_5734), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49046_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n68541));
    defparam i49046_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49025_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n68541), 
            .O(n68520));
    defparam i49025_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51177_4_lut (.I0(n16), .I1(n6_adj_5754), .I2(n19_adj_5734), 
            .I3(n68512), .O(n70672));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51177_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49442_3_lut (.I0(n70112), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n68937));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i49442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51364_4_lut (.I0(n68937), .I1(n70672), .I2(n19_adj_5734), 
            .I3(n68520), .O(n70859));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51364_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51365_3_lut (.I0(n70859), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n70860));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51365_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51261_3_lut (.I0(n70860), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n70756));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51261_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44925_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n294), .I3(GND_net), 
            .O(n64411));
    defparam i44925_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i26_3_lut (.I0(n70756), .I1(n298), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44929_3_lut (.I0(duty[13]), .I1(duty[21]), .I2(n294), .I3(GND_net), 
            .O(n64415));
    defparam i44929_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i45007_4_lut (.I0(duty[15]), .I1(n64411), .I2(duty[20]), .I3(n294), 
            .O(n64493));
    defparam i45007_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i44921_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n64407));
    defparam i44921_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut (.I0(n294), .I1(n64493), .I2(n64415), .I3(n26), 
            .O(n22_adj_5859));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i45005_4_lut (.I0(duty[19]), .I1(n64407), .I2(duty[16]), .I3(n294), 
            .O(n64491));
    defparam i45005_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 n9946_bdd_4_lut_51840 (.I0(n9946), .I1(current[15]), .I2(duty[17]), 
            .I3(n9944), .O(n71361));
    defparam n9946_bdd_4_lut_51840.LUT_INIT = 16'he4aa;
    SB_LUT4 n71361_bdd_4_lut (.I0(n71361), .I1(duty[14]), .I2(n4929), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[14]));
    defparam n71361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i48443_4_lut (.I0(n21_adj_5765), .I1(n19_adj_5766), .I2(n17_adj_5767), 
            .I3(n9_adj_5773), .O(n67938));
    defparam i48443_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49449_3_lut (.I0(n15_adj_5769), .I1(n13_adj_5770), .I2(n11_adj_5771), 
            .I3(GND_net), .O(n68944));
    defparam i49449_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i49374_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n68944), .O(n68869));
    defparam i49374_4_lut.LUT_INIT = 16'h7eff;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i49356_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5769), .O(n68851));
    defparam i49356_4_lut.LUT_INIT = 16'hff7e;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i49481_4_lut (.I0(n9_adj_5773), .I1(n7_adj_5775), .I2(current[2]), 
            .I3(duty[2]), .O(n68976));
    defparam i49481_4_lut.LUT_INIT = 16'heffe;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50285_4_lut (.I0(n15_adj_5769), .I1(n13_adj_5770), .I2(n11_adj_5771), 
            .I3(n68976), .O(n69780));
    defparam i50285_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50255_4_lut (.I0(n21_adj_5765), .I1(n19_adj_5766), .I2(n17_adj_5767), 
            .I3(n69780), .O(n69750));
    defparam i50255_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY add_151_30 (.CI(n52731), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n52732));
    SB_LUT4 add_1190_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n52826), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_24_lut (.I0(GND_net), .I1(GND_net), .I2(n11435), 
            .I3(n52825), .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n52730), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_24 (.CI(n52825), .I0(GND_net), .I1(n11435), .CO(n52826));
    SB_LUT4 add_1190_23_lut (.I0(GND_net), .I1(GND_net), .I2(n11437), 
            .I3(n52824), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_23_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dti_counter_2038__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n30237), 
            .D(n38), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n30237), 
            .D(n39), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n30237), 
            .D(n40_adj_5842), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n30237), 
            .D(n41), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n30237), 
            .D(n42), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n30237), 
            .D(n43_adj_5843), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n30237), 
            .D(n44), .R(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_CARRY add_1190_23 (.CI(n52824), .I0(GND_net), .I1(n11437), .CO(n52825));
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n62946));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n60952));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_1190_22_lut (.I0(GND_net), .I1(GND_net), .I2(n11439), 
            .I3(n52823), .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_22 (.CI(n52823), .I0(GND_net), .I1(n11439), .CO(n52824));
    SB_LUT4 add_1190_21_lut (.I0(GND_net), .I1(GND_net), .I2(n11441), 
            .I3(n52822), .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50927_4_lut (.I0(current[15]), .I1(n23_adj_5763), .I2(duty[12]), 
            .I3(n69750), .O(n70422));
    defparam i50927_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_1190_21 (.CI(n52822), .I0(GND_net), .I1(n11441), .CO(n52823));
    SB_LUT4 add_1190_20_lut (.I0(GND_net), .I1(GND_net), .I2(n11443), 
            .I3(n52821), .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9946_bdd_4_lut_51835 (.I0(n9946), .I1(current[15]), .I2(duty[16]), 
            .I3(n9944), .O(n71355));
    defparam n9946_bdd_4_lut_51835.LUT_INIT = 16'he4aa;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i49382_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n70422), .O(n68877));
    defparam i49382_4_lut.LUT_INIT = 16'h7eff;
    SB_CARRY add_1190_20 (.CI(n52821), .I0(GND_net), .I1(n11443), .CO(n52822));
    SB_LUT4 add_1190_19_lut (.I0(GND_net), .I1(GND_net), .I2(n11445), 
            .I3(n52820), .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50609_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n68877), .O(n70104));
    defparam i50609_4_lut.LUT_INIT = 16'hff7e;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i51185_4_lut (.I0(current[15]), .I1(duty[17]), .I2(duty[18]), 
            .I3(n70104), .O(n70680));
    defparam i51185_4_lut.LUT_INIT = 16'hff7e;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50941_3_lut (.I0(n6_adj_5776), .I1(duty[10]), .I2(n21_adj_5765), 
            .I3(GND_net), .O(n70436));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50941_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50942_3_lut (.I0(n70436), .I1(duty[11]), .I2(n23_adj_5763), 
            .I3(GND_net), .O(n70437));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50942_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50241_4_lut (.I0(current[15]), .I1(n23_adj_5763), .I2(duty[12]), 
            .I3(n67938), .O(n69736));
    defparam i50241_4_lut.LUT_INIT = 16'hffde;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5774), .I1(duty[9]), .I2(n19_adj_5766), 
            .I3(GND_net), .O(n16_adj_5768));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50631_3_lut (.I0(n70437), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n22_adj_5764));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50631_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5777));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i50925_3_lut (.I0(n4_adj_5777), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n70420));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50925_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i48348_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n68869), .O(n67843));
    defparam i48348_4_lut.LUT_INIT = 16'h5adb;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY add_1190_19 (.CI(n52820), .I0(GND_net), .I1(n11445), .CO(n52821));
    SB_LUT4 add_1190_18_lut (.I0(GND_net), .I1(GND_net), .I2(n11447), 
            .I3(n52819), .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_11 (.CI(n52712), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n52713));
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n52704), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_18 (.CI(n52819), .I0(GND_net), .I1(n11447), .CO(n52820));
    SB_CARRY add_151_29 (.CI(n52730), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n52731));
    SB_LUT4 add_1190_17_lut (.I0(GND_net), .I1(GND_net), .I2(n11449), 
            .I3(n52818), .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_17 (.CI(n52818), .I0(GND_net), .I1(n11449), .CO(n52819));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n52729), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n30093), 
            .D(n1251), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 add_1190_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11451), 
            .I3(n52817), .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_16 (.CI(n52817), .I0(GND_net), .I1(n11451), .CO(n52818));
    SB_LUT4 add_1190_15_lut (.I0(GND_net), .I1(GND_net), .I2(n11453), 
            .I3(n52816), .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_15 (.CI(n52816), .I0(GND_net), .I1(n11453), .CO(n52817));
    SB_LUT4 add_1190_14_lut (.I0(GND_net), .I1(GND_net), .I2(n11455), 
            .I3(n52815), .O(n4931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22591_2_lut (.I0(n25253), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n40683));
    defparam i22591_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71355_bdd_4_lut (.I0(n71355), .I1(duty[13]), .I2(n4930), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[13]));
    defparam n71355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 dti_counter_2038_mux_6_i1_4_lut (.I0(n45), .I1(n15_adj_5778), 
            .I2(n40683), .I3(dti_counter[0]), .O(n55));   // verilog/TinyFPGA_B.v(174[23:37])
    defparam dti_counter_2038_mux_6_i1_4_lut.LUT_INIT = 16'ha3a0;
    SB_CARRY add_1190_14 (.CI(n52815), .I0(GND_net), .I1(n11455), .CO(n52816));
    SB_LUT4 add_1190_13_lut (.I0(GND_net), .I1(GND_net), .I2(n11457), 
            .I3(n52814), .O(n4932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_13 (.CI(n52814), .I0(GND_net), .I1(n11457), .CO(n52815));
    SB_LUT4 add_1190_12_lut (.I0(GND_net), .I1(GND_net), .I2(n11459), 
            .I3(n52813), .O(n4933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_28 (.CI(n52729), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n52730));
    SB_CARRY add_1190_12 (.CI(n52813), .I0(GND_net), .I1(n11459), .CO(n52814));
    SB_LUT4 add_1190_11_lut (.I0(GND_net), .I1(GND_net), .I2(n11461), 
            .I3(n52812), .O(n4934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_11 (.CI(n52812), .I0(GND_net), .I1(n11461), .CO(n52813));
    SB_LUT4 add_1190_10_lut (.I0(GND_net), .I1(GND_net), .I2(n11463), 
            .I3(n52811), .O(n4935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_10 (.CI(n52811), .I0(GND_net), .I1(n11463), .CO(n52812));
    SB_LUT4 add_1190_9_lut (.I0(GND_net), .I1(GND_net), .I2(n11465), .I3(n52810), 
            .O(n4936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_9 (.CI(n52810), .I0(GND_net), .I1(n11465), .CO(n52811));
    SB_LUT4 add_1190_8_lut (.I0(GND_net), .I1(GND_net), .I2(n11467), .I3(n52809), 
            .O(n4937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n52728), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_8 (.CI(n52809), .I0(GND_net), .I1(n11467), .CO(n52810));
    SB_LUT4 add_1190_7_lut (.I0(GND_net), .I1(GND_net), .I2(n11469), .I3(n52808), 
            .O(n4938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_7 (.CI(n52808), .I0(GND_net), .I1(n11469), .CO(n52809));
    SB_LUT4 add_1190_6_lut (.I0(GND_net), .I1(GND_net), .I2(n11471), .I3(n52807), 
            .O(n4939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_6 (.CI(n52807), .I0(GND_net), .I1(n11471), .CO(n52808));
    SB_LUT4 add_1190_5_lut (.I0(GND_net), .I1(GND_net), .I2(n11473), .I3(n52806), 
            .O(n4940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_5 (.CI(n52806), .I0(GND_net), .I1(n11473), .CO(n52807));
    SB_LUT4 add_1190_4_lut (.I0(GND_net), .I1(GND_net), .I2(n11475), .I3(n52805), 
            .O(n4941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_4 (.CI(n52805), .I0(GND_net), .I1(n11475), .CO(n52806));
    SB_LUT4 add_1190_3_lut (.I0(GND_net), .I1(GND_net), .I2(n11477), .I3(n52804), 
            .O(n4942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_3 (.CI(n52804), .I0(GND_net), .I1(n11477), .CO(n52805));
    SB_LUT4 add_1190_2_lut (.I0(GND_net), .I1(GND_net), .I2(n10009), .I3(VCC_net), 
            .O(n4943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_23_lut (.I0(GND_net), .I1(n21520), .I2(encoder1_position[23]), 
            .I3(n53891), .O(n20274)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_22_lut (.I0(GND_net), .I1(n21521), .I2(encoder1_position[22]), 
            .I3(n53890), .O(n20275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_22 (.CI(n53890), .I0(n21521), .I1(encoder1_position[22]), 
            .CO(n53891));
    SB_LUT4 add_5385_21_lut (.I0(GND_net), .I1(n21522), .I2(encoder1_position[21]), 
            .I3(n53889), .O(n20276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_21 (.CI(n53889), .I0(n21522), .I1(encoder1_position[21]), 
            .CO(n53890));
    SB_CARRY add_1190_2 (.CI(VCC_net), .I0(GND_net), .I1(n10009), .CO(n52804));
    SB_LUT4 add_5385_20_lut (.I0(GND_net), .I1(n21523), .I2(encoder1_position[20]), 
            .I3(n53888), .O(n20277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_20 (.CI(n53888), .I0(n21523), .I1(encoder1_position[20]), 
            .CO(n53889));
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n30015), .D(GHC_N_391), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n30015), .D(GHB_N_377), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n30015), .D(GHA_N_355), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i22594_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i22594_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5869), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n52711), .O(n1243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22593_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i22593_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n30015), .D(GLA_N_372), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY add_151_27 (.CI(n52728), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n52729));
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n30015), .D(GLB_N_386), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n30015), .D(GLC_N_400), 
            .R(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 add_5385_19_lut (.I0(GND_net), .I1(n21524), .I2(encoder1_position[19]), 
            .I3(n53887), .O(n20278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_19 (.CI(n53887), .I0(n21524), .I1(encoder1_position[19]), 
            .CO(n53888));
    SB_LUT4 add_5385_18_lut (.I0(GND_net), .I1(n21525), .I2(encoder1_position[18]), 
            .I3(n53886), .O(n20279)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_18_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n52727), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_18 (.CI(n53886), .I0(n21525), .I1(encoder1_position[18]), 
            .CO(n53887));
    SB_LUT4 i22714_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i22714_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_151_26 (.CI(n52727), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n52728));
    SB_CARRY add_151_10 (.CI(n52711), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n52712));
    SB_CARRY add_151_3 (.CI(n52704), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n52705));
    SB_LUT4 add_5385_17_lut (.I0(GND_net), .I1(n21526), .I2(encoder1_position[17]), 
            .I3(n53885), .O(n20280)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n52710), .O(n1244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n52726), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_17 (.CI(n53885), .I0(n21526), .I1(encoder1_position[17]), 
            .CO(n53886));
    SB_CARRY add_151_25 (.CI(n52726), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n52727));
    SB_LUT4 add_5385_16_lut (.I0(GND_net), .I1(n21527), .I2(encoder1_position[16]), 
            .I3(n53884), .O(n20281)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_16 (.CI(n53884), .I0(n21527), .I1(encoder1_position[16]), 
            .CO(n53885));
    SB_LUT4 add_5385_15_lut (.I0(GND_net), .I1(n21528), .I2(encoder1_position[15]), 
            .I3(n53883), .O(n20282)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_15 (.CI(n53883), .I0(n21528), .I1(encoder1_position[15]), 
            .CO(n53884));
    SB_LUT4 add_5385_14_lut (.I0(GND_net), .I1(n21529), .I2(encoder1_position[14]), 
            .I3(n53882), .O(n20283)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_14 (.CI(n53882), .I0(n21529), .I1(encoder1_position[14]), 
            .CO(n53883));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n52725), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5385_13_lut (.I0(GND_net), .I1(n21530), .I2(encoder1_position[13]), 
            .I3(n53881), .O(n20284)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n52725), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n52726));
    SB_CARRY add_5385_13 (.CI(n53881), .I0(n21530), .I1(encoder1_position[13]), 
            .CO(n53882));
    SB_LUT4 add_5385_12_lut (.I0(GND_net), .I1(n21531), .I2(encoder1_position[12]), 
            .I3(n53880), .O(n20285)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_12 (.CI(n53880), .I0(n21531), .I1(encoder1_position[12]), 
            .CO(n53881));
    SB_LUT4 add_5385_11_lut (.I0(GND_net), .I1(n21532), .I2(encoder1_position[11]), 
            .I3(n53879), .O(n20286)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_11 (.CI(n53879), .I0(n21532), .I1(encoder1_position[11]), 
            .CO(n53880));
    SB_LUT4 add_5385_10_lut (.I0(GND_net), .I1(n21533), .I2(encoder1_position[10]), 
            .I3(n53878), .O(n20287)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_10 (.CI(n53878), .I0(n21533), .I1(encoder1_position[10]), 
            .CO(n53879));
    SB_LUT4 add_5385_9_lut (.I0(GND_net), .I1(n21534), .I2(encoder1_position[9]), 
            .I3(n53877), .O(n20288)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_9 (.CI(n53877), .I0(n21534), .I1(encoder1_position[9]), 
            .CO(n53878));
    SB_LUT4 add_5385_8_lut (.I0(GND_net), .I1(n21535), .I2(encoder1_position[8]), 
            .I3(n53876), .O(n20289)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_8 (.CI(n53876), .I0(n21535), .I1(encoder1_position[8]), 
            .CO(n53877));
    SB_LUT4 add_5385_7_lut (.I0(GND_net), .I1(n21536), .I2(encoder1_position[7]), 
            .I3(n53875), .O(n20290)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_7 (.CI(n53875), .I0(n21536), .I1(encoder1_position[7]), 
            .CO(n53876));
    SB_LUT4 add_5385_6_lut (.I0(GND_net), .I1(n21537), .I2(encoder1_position[6]), 
            .I3(n53874), .O(n20291)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_6 (.CI(n53874), .I0(n21537), .I1(encoder1_position[6]), 
            .CO(n53875));
    SB_LUT4 add_5385_5_lut (.I0(GND_net), .I1(n21538), .I2(encoder1_position[5]), 
            .I3(n53873), .O(n20292)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_5 (.CI(n53873), .I0(n21538), .I1(encoder1_position[5]), 
            .CO(n53874));
    SB_LUT4 add_5385_4_lut (.I0(GND_net), .I1(n21539), .I2(encoder1_position[4]), 
            .I3(n53872), .O(n20293)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48988_3_lut_4_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(current_limit[5]), .I3(current[5]), .O(n68483));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i48988_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5385_4 (.CI(n53872), .I0(n21539), .I1(encoder1_position[4]), 
            .CO(n53873));
    SB_LUT4 LessThan_14_i12_3_lut_3_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(current_limit[5]), .I3(GND_net), .O(n12_adj_5761));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i12_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_5385_3_lut (.I0(GND_net), .I1(n21540), .I2(encoder1_position[3]), 
            .I3(n53871), .O(n20294)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5385_3 (.CI(n53871), .I0(n21540), .I1(encoder1_position[3]), 
            .CO(n53872));
    SB_LUT4 add_5385_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n20295)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5385_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_51993 (.I0(byte_transmit_counter[3]), 
            .I1(n71220), .I2(n67794), .I3(byte_transmit_counter[4]), .O(n71523));
    defparam byte_transmit_counter_3__bdd_4_lut_51993.LUT_INIT = 16'he4aa;
    SB_LUT4 n71523_bdd_4_lut (.I0(n71523), .I1(n64802), .I2(n7_adj_5847), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n71523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_5385_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n53871));
    SB_LUT4 LessThan_11_i35_rep_50_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n71784));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_50_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51238_3_lut (.I0(n30), .I1(n10_adj_5772), .I2(n68851), .I3(GND_net), 
            .O(n70733));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50629_4_lut (.I0(n70420), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n70124));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50629_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i51392_4_lut (.I0(n70124), .I1(n70733), .I2(n71784), .I3(n67843), 
            .O(n70887));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51392_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51393_3_lut (.I0(n70887), .I1(duty[18]), .I2(current[15]), 
            .I3(GND_net), .O(n70888));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51393_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51366_4_lut (.I0(current[15]), .I1(duty[19]), .I2(duty[20]), 
            .I3(n70680), .O(n70861));
    defparam i51366_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i50281_3_lut (.I0(n22_adj_5764), .I1(n16_adj_5768), .I2(n69736), 
            .I3(GND_net), .O(n69776));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51265_4_lut (.I0(n70888), .I1(duty[20]), .I2(current[15]), 
            .I3(duty[19]), .O(n40));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51265_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i50624_3_lut (.I0(n40), .I1(n69776), .I2(n70861), .I3(GND_net), 
            .O(n70119));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50624_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n52962), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n52961), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n52961), .I0(GND_net), .I1(n2), 
            .CO(n52962));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5739), 
            .I3(n52960), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n52960), .I0(GND_net), .I1(n14_adj_5739), 
            .CO(n52961));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5740), 
            .I3(n52959), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n52959), .I0(GND_net), .I1(n15_adj_5740), 
            .CO(n52960));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5741), 
            .I3(n52958), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1815 (.I0(n70119), .I1(current[15]), .I2(duty[21]), 
            .I3(GND_net), .O(n6_adj_5845));
    defparam i2_3_lut_adj_1815.LUT_INIT = 16'hfefe;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n52958), .I0(GND_net), .I1(n16_adj_5741), 
            .CO(n52959));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5742), 
            .I3(n52957), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n52957), .I0(GND_net), .I1(n17_adj_5742), 
            .CO(n52958));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5743), 
            .I3(n52956), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[31]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[30]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[29]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[28]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[27]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[26]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[25]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[24]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 326[6])
    SB_CARRY unary_minus_16_add_3_9 (.CI(n52956), .I0(GND_net), .I1(n18_adj_5743), 
            .CO(n52957));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5744), 
            .I3(n52955), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n52955), .I0(GND_net), .I1(n19_adj_5744), 
            .CO(n52956));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5745), 
            .I3(n52954), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n52954), .I0(GND_net), .I1(n20_adj_5745), 
            .CO(n52955));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5746), 
            .I3(n52953), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n52953), .I0(GND_net), .I1(n21_adj_5746), 
            .CO(n52954));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5747), 
            .I3(n52952), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n52952), .I0(GND_net), .I1(n22_adj_5747), 
            .CO(n52953));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5748), 
            .I3(n52951), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n52951), .I0(GND_net), .I1(n23_adj_5748), 
            .CO(n52952));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5749), 
            .I3(n52950), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n52950), .I0(GND_net), .I1(n24_adj_5749), 
            .CO(n52951));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n41195), .I1(GND_net), .I2(n25_adj_5750), 
            .I3(VCC_net), .O(n67567)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5750), 
            .CO(n52950));
    SB_LUT4 i7_4_lut (.I0(duty[22]), .I1(duty[23]), .I2(n6_adj_5845), 
            .I3(n260), .O(n9946));
    defparam i7_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n52724), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n52724), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n52725));
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n52723), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n58271));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_CARRY add_151_22 (.CI(n52723), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n52724));
    SB_LUT4 n9946_bdd_4_lut_51830 (.I0(n9946), .I1(current[5]), .I2(duty[8]), 
            .I3(n9944), .O(n71349));
    defparam n9946_bdd_4_lut_51830.LUT_INIT = 16'he4aa;
    SB_LUT4 n71349_bdd_4_lut (.I0(n71349), .I1(duty[5]), .I2(n4938), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n71349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n30093), 
            .D(n1250), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n30093), 
            .D(n1249), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n30093), 
            .D(n1248), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n30093), 
            .D(n1247), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n30093), 
            .D(n1246), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n30093), 
            .D(n1245), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n30093), 
            .D(n1244), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n30093), 
            .D(n1243), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n30093), 
            .D(n1242), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n30093), 
            .D(n1241), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n30093), 
            .D(n1240), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n30093), 
            .D(n1239), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n30093), 
            .D(n1238), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n30093), 
            .D(n1237), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n30093), 
            .D(n1236), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n30093), 
            .D(n1235), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n30093), 
            .D(n1234), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n30093), 
            .D(n1233), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n30093), 
            .D(n1232), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n30093), 
            .D(n1231), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n30093), 
            .D(n1230), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n30093), 
            .D(n1229), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n30093), 
            .D(n1228), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n30093), 
            .D(n1227), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n30093), 
            .D(n1226), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n30093), 
            .D(n1225), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n30093), 
            .D(n1224), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n30093), 
            .D(n1223), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n30093), 
            .D(n1222), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n30093), 
            .D(n1221), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n30093), 
            .D(n1220), .R(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n52722), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n58351));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i49339_2_lut (.I0(displacement[0]), .I1(n15_adj_5808), .I2(GND_net), 
            .I3(GND_net), .O(n67541));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam i49339_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13933_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n59777), .I3(GND_net), .O(n32124));   // verilog/coms.v(130[12] 305[6])
    defparam i13933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13936_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n59777), .I3(GND_net), .O(n32127));   // verilog/coms.v(130[12] 305[6])
    defparam i13936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13939_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n59777), .I3(GND_net), .O(n32130));   // verilog/coms.v(130[12] 305[6])
    defparam i13939_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_9 (.CI(n52710), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n52711));
    SB_CARRY add_151_21 (.CI(n52722), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n52723));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5796), .I3(n52880), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3), .I3(n52879), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n52709), .O(n1245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_8 (.CI(n52709), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n52710));
    SB_LUT4 add_5383_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(encoder1_position[21]), 
            .I3(n53792), .O(n21520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(encoder1_position[20]), 
            .I3(n53791), .O(n21521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_21 (.CI(n53791), .I0(encoder1_position[19]), .I1(encoder1_position[20]), 
            .CO(n53792));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n52879), .I0(encoder0_position_scaled[22]), 
            .I1(n3), .CO(n52880));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5795), .I3(n52878), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n52878), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5795), .CO(n52879));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5814), .I3(n52877), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n52721), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_20 (.CI(n52721), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n52722));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n52720), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(encoder1_position[19]), 
            .I3(n53790), .O(n21522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n52877), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5814), .CO(n52878));
    SB_CARRY add_5383_20 (.CI(n53790), .I0(encoder1_position[18]), .I1(encoder1_position[19]), 
            .CO(n53791));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5813), .I3(n52876), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(encoder1_position[18]), 
            .I3(n53789), .O(n21523)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_19 (.CI(n53789), .I0(encoder1_position[17]), .I1(encoder1_position[18]), 
            .CO(n53790));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n52876), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5813), .CO(n52877));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5812), .I3(n52875), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n52875), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5812), .CO(n52876));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5811), .I3(n52874), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n52874), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5811), .CO(n52875));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5810), .I3(n52873), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n52873), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5810), .CO(n52874));
    SB_LUT4 add_5383_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(encoder1_position[17]), 
            .I3(n53788), .O(n21524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_19 (.CI(n52720), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n52721));
    SB_CARRY add_5383_18 (.CI(n53788), .I0(encoder1_position[16]), .I1(encoder1_position[17]), 
            .CO(n53789));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5794), .I3(n52872), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n52872), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5794), .CO(n52873));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5793), .I3(n52871), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n52871), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5793), .CO(n52872));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5792), .I3(n52870), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(encoder1_position[16]), 
            .I3(n53787), .O(n21525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_17 (.CI(n53787), .I0(encoder1_position[15]), .I1(encoder1_position[16]), 
            .CO(n53788));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n52870), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5792), .CO(n52871));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5738), .I3(n52869), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n52869), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5738), .CO(n52870));
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n52719), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(encoder1_position[15]), 
            .I3(n53786), .O(n21526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_16 (.CI(n53786), .I0(encoder1_position[14]), .I1(encoder1_position[15]), 
            .CO(n53787));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n52868), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n52868), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n52869));
    SB_CARRY add_151_18 (.CI(n52719), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n52720));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n52718), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n52718), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n52719));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n52708), .O(n1246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(encoder1_position[14]), 
            .I3(n53785), .O(n21527)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5737), .I3(n52867), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n52867), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5737), .CO(n52868));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n52717), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n52704));
    SB_CARRY add_151_16 (.CI(n52717), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n52718));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5736), .I3(n52866), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n52866), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5736), .CO(n52867));
    SB_CARRY add_151_7 (.CI(n52708), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n52709));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n52716), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n52707), .O(n1247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_15 (.CI(n53785), .I0(encoder1_position[13]), .I1(encoder1_position[14]), 
            .CO(n53786));
    SB_LUT4 add_5383_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(encoder1_position[13]), 
            .I3(n53784), .O(n21528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5735), .I3(n52865), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n52865), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5735), .CO(n52866));
    SB_CARRY add_151_15 (.CI(n52716), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n52717));
    SB_CARRY add_5383_14 (.CI(n53784), .I0(encoder1_position[12]), .I1(encoder1_position[13]), 
            .CO(n53785));
    SB_LUT4 add_5383_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(encoder1_position[12]), 
            .I3(n53783), .O(n21529)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_13 (.CI(n53783), .I0(encoder1_position[11]), .I1(encoder1_position[12]), 
            .CO(n53784));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18), .I3(n52864), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n52864), .I0(encoder0_position_scaled[7]), 
            .I1(n18), .CO(n52865));
    SB_CARRY add_151_6 (.CI(n52707), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n52708));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n52715), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n52863), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(encoder1_position[11]), 
            .I3(n53782), .O(n21530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_12 (.CI(n53782), .I0(encoder1_position[10]), .I1(encoder1_position[11]), 
            .CO(n53783));
    SB_LUT4 add_5383_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(encoder1_position[10]), 
            .I3(n53781), .O(n21531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_5383_11 (.CI(n53781), .I0(encoder1_position[9]), .I1(encoder1_position[10]), 
            .CO(n53782));
    SB_LUT4 add_5383_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(encoder1_position[9]), 
            .I3(n53780), .O(n21532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_10 (.CI(n53780), .I0(encoder1_position[8]), .I1(encoder1_position[9]), 
            .CO(n53781));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n52863), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n52864));
    SB_LUT4 add_5383_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(encoder1_position[8]), 
            .I3(n53779), .O(n21533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_9 (.CI(n53779), .I0(encoder1_position[7]), .I1(encoder1_position[8]), 
            .CO(n53780));
    SB_LUT4 add_5383_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(encoder1_position[7]), 
            .I3(n53778), .O(n21534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_8 (.CI(n53778), .I0(encoder1_position[6]), .I1(encoder1_position[7]), 
            .CO(n53779));
    SB_LUT4 add_5383_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(encoder1_position[6]), 
            .I3(n53777), .O(n21535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_7 (.CI(n53777), .I0(encoder1_position[5]), .I1(encoder1_position[6]), 
            .CO(n53778));
    SB_LUT4 add_5383_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(encoder1_position[5]), 
            .I3(n53776), .O(n21536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_6 (.CI(n53776), .I0(encoder1_position[4]), .I1(encoder1_position[5]), 
            .CO(n53777));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n52862), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[4]), 
            .I3(n53775), .O(n21537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n52862), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n52863));
    SB_CARRY add_5383_5 (.CI(n53775), .I0(encoder1_position[3]), .I1(encoder1_position[4]), 
            .CO(n53776));
    SB_LUT4 add_5383_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[3]), 
            .I3(n53774), .O(n21538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_4 (.CI(n53774), .I0(encoder1_position[2]), .I1(encoder1_position[3]), 
            .CO(n53775));
    SB_LUT4 add_5383_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n53773), .O(n21539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_3 (.CI(n53773), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n53774));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n52861), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n21540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_91[1]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13605_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n30673), 
            .I3(GND_net), .O(n31796));   // verilog/coms.v(130[12] 305[6])
    defparam i13605_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13943_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n59777), .I3(GND_net), .O(n32134));   // verilog/coms.v(130[12] 305[6])
    defparam i13943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13946_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n59777), .I3(GND_net), .O(n32137));   // verilog/coms.v(130[12] 305[6])
    defparam i13946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13958_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n59779), .I3(GND_net), .O(n32149));   // verilog/coms.v(130[12] 305[6])
    defparam i13958_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_91[2]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i3_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_5383_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n53773));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n52861), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n52862));
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_91[3]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_91[4]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n9946_bdd_4_lut_51825 (.I0(n9946), .I1(current[15]), .I2(duty[15]), 
            .I3(n9944), .O(n71337));
    defparam n9946_bdd_4_lut_51825.LUT_INIT = 16'he4aa;
    SB_LUT4 n71337_bdd_4_lut (.I0(n71337), .I1(duty[12]), .I2(n4931), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[12]));
    defparam n71337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5734));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45086_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64581));
    defparam i45086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45087_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64582));
    defparam i45087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45090_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64585));
    defparam i45090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45089_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64584));
    defparam i45089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45386_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64881));
    defparam i45386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45387_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64882));
    defparam i45387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45084_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64579));
    defparam i45084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45083_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64578));
    defparam i45083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_91[5]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13949_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n59777), .I3(GND_net), .O(n32140));   // verilog/coms.v(130[12] 305[6])
    defparam i13949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5735));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5736));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13952_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n59777), .I3(GND_net), .O(n32143));   // verilog/coms.v(130[12] 305[6])
    defparam i13952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5737));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_91[11]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_91[12]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5738));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5792));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_91[13]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5793));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_91[14]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n23_adj_5860), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5233), .I3(r_SM_Main_adj_5942[0]), .O(n63671));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfeff;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5794));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_91[15]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5810));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63671), .O(n61776));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_91[16]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_243_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_91[6]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5811));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5812));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5813));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_91[17]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5814));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5795));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5796));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_91[18]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_91[19]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_91[20]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_91[21]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_91[22]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_91[23]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13596_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n30673), 
            .I3(GND_net), .O(n31787));   // verilog/coms.v(130[12] 305[6])
    defparam i13596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23141_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n39602), .O(n41236));
    defparam i23141_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i13491_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n30039), .I3(GND_net), .O(n31682));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13593_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n30673), 
            .I3(GND_net), .O(n31784));   // verilog/coms.v(130[12] 305[6])
    defparam i13593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14059_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[0]), 
            .I2(n10_adj_5846), .I3(n27930), .O(n32250));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14059_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13502_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n25082), .I3(GND_net), .O(n31693));   // verilog/coms.v(130[12] 305[6])
    defparam i13502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13504_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n25151), .I3(GND_net), .O(n31695));   // verilog/coms.v(130[12] 305[6])
    defparam i13504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13581_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n30671), 
            .I3(GND_net), .O(n31772));   // verilog/coms.v(130[12] 305[6])
    defparam i13581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13575_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n30671), 
            .I3(GND_net), .O(n31766));   // verilog/coms.v(130[12] 305[6])
    defparam i13575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n4_adj_5781), .I1(r_SM_Main[1]), .I2(n6_adj_5865), 
            .I3(r_Bit_Index[0]), .O(n63569));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63569), .O(n63575));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1820 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63575), .O(n63581));
    defparam i1_4_lut_adj_1820.LUT_INIT = 16'hfffe;
    SB_LUT4 i14095_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n63581), 
            .I3(n27), .O(n32286));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14095_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13508_3_lut (.I0(current[0]), .I1(data_adj_5926[0]), .I2(n30062), 
            .I3(GND_net), .O(n31699));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14108_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[0]), .I2(n11_adj_5784), 
            .I3(state_7__N_4319), .O(n32299));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14108_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13961_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n59779), .I3(GND_net), .O(n32152));   // verilog/coms.v(130[12] 305[6])
    defparam i13961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13516_3_lut (.I0(b_prev_adj_5789), .I1(b_new_adj_5906[1]), 
            .I2(debounce_cnt_N_3833_adj_5790), .I3(GND_net), .O(n31707));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13517_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3178), .I3(GND_net), 
            .O(n31708));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13566_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n30671), 
            .I3(GND_net), .O(n31757));   // verilog/coms.v(130[12] 305[6])
    defparam i13566_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13563_3_lut (.I0(\data_in_frame[2] [7]), .I1(rx_data[7]), .I2(n30669), 
            .I3(GND_net), .O(n31754));   // verilog/coms.v(130[12] 305[6])
    defparam i13563_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13560_3_lut (.I0(\data_in_frame[2] [6]), .I1(rx_data[6]), .I2(n30669), 
            .I3(GND_net), .O(n31751));   // verilog/coms.v(130[12] 305[6])
    defparam i13560_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13557_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n30669), 
            .I3(GND_net), .O(n31748));   // verilog/coms.v(130[12] 305[6])
    defparam i13557_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14253_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n25151), .I3(GND_net), .O(n32444));   // verilog/coms.v(130[12] 305[6])
    defparam i14253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14254_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n25151), .I3(GND_net), .O(n32445));   // verilog/coms.v(130[12] 305[6])
    defparam i14254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14255_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n25151), .I3(GND_net), .O(n32446));   // verilog/coms.v(130[12] 305[6])
    defparam i14255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14256_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n25151), .I3(GND_net), .O(n32447));   // verilog/coms.v(130[12] 305[6])
    defparam i14256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14257_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n25151), .I3(GND_net), .O(n32448));   // verilog/coms.v(130[12] 305[6])
    defparam i14257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14258_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n25151), .I3(GND_net), .O(n32449));   // verilog/coms.v(130[12] 305[6])
    defparam i14258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14259_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n25151), .I3(GND_net), .O(n32450));   // verilog/coms.v(130[12] 305[6])
    defparam i14259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14260_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n25151), .I3(GND_net), .O(n32451));   // verilog/coms.v(130[12] 305[6])
    defparam i14260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14261_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n25151), .I3(GND_net), .O(n32452));   // verilog/coms.v(130[12] 305[6])
    defparam i14261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14263_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n25151), .I3(GND_net), .O(n32454));   // verilog/coms.v(130[12] 305[6])
    defparam i14263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19776_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n25151), .I3(GND_net), .O(n32455));
    defparam i19776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19771_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n25151), .I3(GND_net), .O(n37917));
    defparam i19771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14266_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n25151), .I3(GND_net), .O(n32457));   // verilog/coms.v(130[12] 305[6])
    defparam i14266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14267_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n25151), .I3(GND_net), .O(n32458));   // verilog/coms.v(130[12] 305[6])
    defparam i14267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20097_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n25151), .I3(GND_net), .O(n32459));
    defparam i20097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19930_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n25151), .I3(GND_net), .O(n32460));
    defparam i19930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14270_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n25151), .I3(GND_net), .O(n32461));   // verilog/coms.v(130[12] 305[6])
    defparam i14270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14271_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n25151), .I3(GND_net), .O(n32462));   // verilog/coms.v(130[12] 305[6])
    defparam i14271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13554_3_lut (.I0(\data_in_frame[2] [4]), .I1(rx_data[4]), .I2(n30669), 
            .I3(GND_net), .O(n31745));   // verilog/coms.v(130[12] 305[6])
    defparam i13554_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19189_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n25082), .I3(GND_net), .O(n32467));
    defparam i19189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14277_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n25082), .I3(GND_net), .O(n32468));   // verilog/coms.v(130[12] 305[6])
    defparam i14277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14278_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n25082), .I3(GND_net), .O(n32469));   // verilog/coms.v(130[12] 305[6])
    defparam i14278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14279_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n25082), .I3(GND_net), .O(n32470));   // verilog/coms.v(130[12] 305[6])
    defparam i14279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19295_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n25082), .I3(GND_net), .O(n32471));
    defparam i19295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14281_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n25082), .I3(GND_net), .O(n32472));   // verilog/coms.v(130[12] 305[6])
    defparam i14281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14283_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n25082), .I3(GND_net), .O(n32474));   // verilog/coms.v(130[12] 305[6])
    defparam i14283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14284_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n25082), .I3(GND_net), .O(n32475));   // verilog/coms.v(130[12] 305[6])
    defparam i14284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14286_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n25082), .I3(GND_net), .O(n32477));   // verilog/coms.v(130[12] 305[6])
    defparam i14286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14287_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n25082), .I3(GND_net), .O(n32478));   // verilog/coms.v(130[12] 305[6])
    defparam i14287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14288_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n25082), .I3(GND_net), .O(n32479));   // verilog/coms.v(130[12] 305[6])
    defparam i14288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14289_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n25082), .I3(GND_net), .O(n32480));   // verilog/coms.v(130[12] 305[6])
    defparam i14289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14290_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n25082), .I3(GND_net), .O(n32481));   // verilog/coms.v(130[12] 305[6])
    defparam i14290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14291_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n25082), .I3(GND_net), .O(n32482));   // verilog/coms.v(130[12] 305[6])
    defparam i14291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14292_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n25082), .I3(GND_net), .O(n32483));   // verilog/coms.v(130[12] 305[6])
    defparam i14292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14293_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n25082), .I3(GND_net), .O(n32484));   // verilog/coms.v(130[12] 305[6])
    defparam i14293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18956_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n25082), .I3(GND_net), .O(n32487));
    defparam i18956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18957_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n25082), .I3(GND_net), .O(n32488));
    defparam i18957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18958_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n25082), .I3(GND_net), .O(n32489));
    defparam i18958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13551_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n30669), 
            .I3(GND_net), .O(n31742));   // verilog/coms.v(130[12] 305[6])
    defparam i13551_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n60082));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n60081));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n31455));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n60080));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n60076));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n60077));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n31451));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n60075));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n60072));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n60073));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n31447));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n60078));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n60079));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n60071));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n31443));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n60074));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset), .I1(n39602), .I2(n8), .I3(GND_net), 
            .O(n30698));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n39602), .I2(GND_net), .I3(GND_net), 
            .O(n39603));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_1836 (.I0(n15_adj_5778), .I1(n25253), .I2(dti), 
            .I3(GND_net), .O(n29991));
    defparam i1_2_lut_3_lut_adj_1836.LUT_INIT = 16'hbaba;
    SB_LUT4 i14011_3_lut_4_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n39603), .I3(n8), .O(n32202));   // verilog/coms.v(130[12] 305[6])
    defparam i14011_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i14605_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2887));   // verilog/coms.v(130[12] 305[6])
    defparam i14605_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14379_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n30039), .I3(GND_net), .O(n32570));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13548_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n30669), 
            .I3(GND_net), .O(n31739));   // verilog/coms.v(130[12] 305[6])
    defparam i13548_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13545_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n30669), 
            .I3(GND_net), .O(n31736));   // verilog/coms.v(130[12] 305[6])
    defparam i13545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14382_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n30039), .I3(GND_net), .O(n32573));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14383_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n338), 
            .I2(n30039), .I3(GND_net), .O(n32574));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14384_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n30039), .I3(GND_net), .O(n32575));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14385_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n30039), .I3(GND_net), .O(n32576));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14386_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n341), 
            .I2(n30039), .I3(GND_net), .O(n32577));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14387_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n30039), .I3(GND_net), .O(n32578));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14388_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n30039), .I3(GND_net), .O(n32579));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14389_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n30039), .I3(GND_net), .O(n32580));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14390_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n30039), .I3(GND_net), .O(n32581));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14391_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n30039), .I3(GND_net), .O(n32582));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14392_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n30039), .I3(GND_net), .O(n32583));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14393_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n30039), .I3(GND_net), .O(n32584));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14394_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n30039), .I3(GND_net), .O(n32585));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14395_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n30039), .I3(GND_net), .O(n32586));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1837 (.I0(n15_adj_5778), .I1(n25253), .I2(dti), 
            .I3(GND_net), .O(n30237));
    defparam i1_2_lut_3_lut_adj_1837.LUT_INIT = 16'heaea;
    SB_LUT4 i14396_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n30039), .I3(GND_net), .O(n32587));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14397_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n30039), .I3(GND_net), .O(n32588));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14398_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n30039), .I3(GND_net), .O(n32589));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14399_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n30039), .I3(GND_net), .O(n32590));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14400_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n30039), .I3(GND_net), .O(n32591));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14401_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n30039), .I3(GND_net), .O(n32592));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14402_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n30039), .I3(GND_net), .O(n32593));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13463_2_lut_3_lut (.I0(n15_adj_5778), .I1(n25253), .I2(dti), 
            .I3(GND_net), .O(n31653));   // verilog/TinyFPGA_B.v(174[23:37])
    defparam i13463_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i14403_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n30039), .I3(GND_net), .O(n32594));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(r_SM_Main[1]), .I1(n6_adj_5865), .I2(r_Bit_Index[0]), 
            .I3(n4_adj_5781), .O(n63533));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_1839 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63533), .O(n63539));
    defparam i1_4_lut_adj_1839.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63539), .O(n63545));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 i14407_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n63545), 
            .I3(n27), .O(n32598));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14407_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63623), .O(n63629));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1842 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63629), .O(n63635));
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_LUT4 i14408_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n63635), 
            .I3(n27), .O(n32599));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14408_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1843 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63587), .O(n63593));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1844 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63593), .O(n63599));
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'hfffe;
    SB_LUT4 i14409_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n63599), 
            .I3(n27), .O(n32600));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14409_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1845 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63641), .O(n63647));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1846 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63647), .O(n63653));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 i14412_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n63653), 
            .I3(n27), .O(n32603));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14412_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1847 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63551), .O(n63557));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63557), .O(n63563));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'hfffe;
    SB_LUT4 i14413_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n63563), 
            .I3(n27), .O(n32604));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14413_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5554_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5554_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63605), .O(n63611));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i5552_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5552_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63611), .O(n63617));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i14414_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n63617), 
            .I3(n27), .O(n32605));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14414_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5556_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i5556_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5558_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i5558_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(o_Rx_DV_N_3488[12]), .I1(n5230), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n63515), .O(n63521));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1852 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5860), 
            .I3(n63521), .O(n63527));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 i14415_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n63527), 
            .I3(n27), .O(n32606));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14415_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14218_3_lut (.I0(\data_in_frame[22] [7]), .I1(rx_data[7]), 
            .I2(n30709), .I3(GND_net), .O(n32409));   // verilog/coms.v(130[12] 305[6])
    defparam i14218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14215_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n30709), .I3(GND_net), .O(n32406));   // verilog/coms.v(130[12] 305[6])
    defparam i14215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14212_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n30709), .I3(GND_net), .O(n32403));   // verilog/coms.v(130[12] 305[6])
    defparam i14212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48686_4_lut (.I0(data_ready), .I1(n6916), .I2(n24_adj_5856), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n67710));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i48686_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i49144_2_lut (.I0(n24_adj_5856), .I1(n6916), .I2(GND_net), 
            .I3(GND_net), .O(n67713));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i49144_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n67713), .I1(n67710), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5848), .O(n58271));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i14205_3_lut (.I0(\data_in_frame[22] [4]), .I1(rx_data[4]), 
            .I2(n30709), .I3(GND_net), .O(n32396));   // verilog/coms.v(130[12] 305[6])
    defparam i14205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14202_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n30709), .I3(GND_net), .O(n32393));   // verilog/coms.v(130[12] 305[6])
    defparam i14202_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14199_3_lut (.I0(\data_in_frame[22] [2]), .I1(rx_data[2]), 
            .I2(n30709), .I3(GND_net), .O(n32390));   // verilog/coms.v(130[12] 305[6])
    defparam i14199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14196_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n30709), .I3(GND_net), .O(n32387));   // verilog/coms.v(130[12] 305[6])
    defparam i14196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[21] [5]), .I1(n30619), .I2(n30708), 
            .I3(rx_data[5]), .O(n59309));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1853 (.I0(\data_in_frame[21] [4]), .I1(n30619), 
            .I2(n30708), .I3(rx_data[4]), .O(n59255));
    defparam i12_4_lut_adj_1853.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[21] [3]), .I1(n61124), .I2(n30708), 
            .I3(rx_data[3]), .O(n59265));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14_4_lut_adj_1854 (.I0(\data_in_frame[21] [2]), .I1(n61124), 
            .I2(n30708), .I3(rx_data[2]), .O(n59263));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1854.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14172_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n30708), .I3(GND_net), .O(n32363));   // verilog/coms.v(130[12] 305[6])
    defparam i14172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13629_3_lut_4_lut (.I0(n1755), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n31820));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13629_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i13627_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n31818));   // verilog/coms.v(130[12] 305[6])
    defparam i13627_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21506_4_lut (.I0(n67702), .I1(n67701), .I2(rx_data[0]), .I3(\data_in_frame[21] [0]), 
            .O(n39619));   // verilog/coms.v(94[13:20])
    defparam i21506_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i21507_3_lut (.I0(n39619), .I1(\data_in_frame[21] [0]), .I2(reset), 
            .I3(GND_net), .O(n32632));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i21507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1855 (.I0(r_SM_Main_adj_5942[0]), .I1(o_Rx_DV_N_3488[24]), 
            .I2(n27), .I3(GND_net), .O(n14_adj_5851));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut_adj_1855.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut_adj_1856 (.I0(n29), .I1(o_Rx_DV_N_3488[12]), .I2(n23_adj_5860), 
            .I3(n5233), .O(n15_adj_5850));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut_adj_1856.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut_adj_1857 (.I0(n15_adj_5850), .I1(n1), .I2(n14_adj_5851), 
            .I3(r_SM_Main_adj_5942[1]), .O(n71737));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut_adj_1857.LUT_INIT = 16'h8000;
    SB_LUT4 i14449_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[1]), 
            .I2(n10_adj_5846), .I3(n27881), .O(n32640));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14449_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14453_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[2]), 
            .I2(n4_adj_5779), .I3(n27930), .O(n32644));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14453_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14454_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[3]), 
            .I2(n4_adj_5779), .I3(n27881), .O(n32645));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14454_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14458_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[4]), 
            .I2(n4_adj_5780), .I3(n27930), .O(n32649));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14459_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[5]), 
            .I2(n4_adj_5780), .I3(n27881), .O(n32650));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14459_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51463_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n40695), .I3(GND_net), .O(n30093));
    defparam i51463_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i14460_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[6]), 
            .I2(n40902), .I3(n27930), .O(n32651));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14460_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i49037_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n67604));
    defparam i49037_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i22703_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n40695), .I3(GND_net), .O(n40795));
    defparam i22703_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1858 (.I0(n8_adj_5815), .I1(n39602), .I2(GND_net), 
            .I3(GND_net), .O(n30621));
    defparam i1_2_lut_adj_1858.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14115_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n30702), .I3(GND_net), .O(n32306));   // verilog/coms.v(130[12] 305[6])
    defparam i14115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1859 (.I0(\data_in_frame[18] [6]), .I1(n30623), 
            .I2(n30702), .I3(rx_data[6]), .O(n59173));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1859.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14109_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n30702), .I3(GND_net), .O(n32300));   // verilog/coms.v(130[12] 305[6])
    defparam i14109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14472_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5919[7]), 
            .I2(n40902), .I3(n27881), .O(n32663));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14472_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14474_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[1]), .I2(n5_adj_5783), 
            .I3(n27938), .O(n32665));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14474_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14475_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[2]), .I2(n5_adj_5809), 
            .I3(n27938), .O(n32666));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14475_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14476_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[3]), .I2(n40832), 
            .I3(n27938), .O(n32667));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14476_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14477_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[4]), .I2(n5_adj_5797), 
            .I3(n27925), .O(n32668));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14477_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14478_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[5]), .I2(n5_adj_5783), 
            .I3(n27925), .O(n32669));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14478_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14479_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[6]), .I2(n5_adj_5809), 
            .I3(n27925), .O(n32670));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14479_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14480_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[7]), .I2(n40832), 
            .I3(n27925), .O(n32671));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14480_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14481_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[8]), .I2(n5_adj_5797), 
            .I3(n27891), .O(n32672));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14481_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14482_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[9]), .I2(n5_adj_5783), 
            .I3(n27891), .O(n32673));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14482_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14483_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[10]), .I2(n5_adj_5809), 
            .I3(n27891), .O(n32674));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14483_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14484_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[11]), .I2(n40832), 
            .I3(n27891), .O(n32675));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14484_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14485_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[12]), .I2(n5_adj_5797), 
            .I3(n27916), .O(n32676));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14485_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14486_4_lut (.I0(CS_MISO_c), .I1(data_adj_5926[15]), .I2(n40832), 
            .I3(n27916), .O(n32677));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14486_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1860 (.I0(n3489), .I1(n89), .I2(reset), 
            .I3(n76), .O(n30708));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1860.LUT_INIT = 16'h0008;
    SB_LUT4 i14099_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n30702), .I3(GND_net), .O(n32290));   // verilog/coms.v(130[12] 305[6])
    defparam i14099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1861 (.I0(\data_in_frame[18] [2]), .I1(n30623), 
            .I2(n30702), .I3(rx_data[2]), .O(n59177));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1861.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_adj_1862 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n60086));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_1862.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1863 (.I0(\data_in_frame[18] [1]), .I1(n30623), 
            .I2(n30702), .I3(rx_data[1]), .O(n59181));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1863.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14087_4_lut (.I0(n63257), .I1(r_Bit_Index[0]), .I2(n60927), 
            .I3(n30084), .O(n32278));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i14087_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i12_4_lut_adj_1864 (.I0(\data_in_frame[18] [0]), .I1(n30623), 
            .I2(n30702), .I3(rx_data[0]), .O(n59185));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1864.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14081_4_lut (.I0(n63255), .I1(r_Bit_Index_adj_5944[0]), .I2(n60925), 
            .I3(n30087), .O(n32272));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i14081_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i12_4_lut_adj_1865 (.I0(\data_in_frame[17] [7]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[7]), .O(n59313));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1865.LUT_INIT = 16'h3a0a;
    SB_LUT4 i21521_4_lut (.I0(n67698), .I1(n67697), .I2(rx_data[6]), .I3(\data_in_frame[17] [6]), 
            .O(n39634));   // verilog/coms.v(94[13:20])
    defparam i21521_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i21522_3_lut (.I0(n39634), .I1(\data_in_frame[17] [6]), .I2(reset), 
            .I3(GND_net), .O(n32704));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i21522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1866 (.I0(\data_in_frame[17] [5]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[5]), .O(n59315));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1866.LUT_INIT = 16'h3a0a;
    SB_LUT4 i13814_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n59773), 
            .I3(GND_net), .O(n32005));   // verilog/coms.v(130[12] 305[6])
    defparam i13814_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1867 (.I0(\data_in_frame[16] [7]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[7]), .O(n59189));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1867.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n59931));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n59925));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n59924));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h4500;
    SB_LUT4 i12_4_lut_adj_1871 (.I0(\data_in_frame[16] [6]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[6]), .O(n59193));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1871.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1872 (.I0(\data_in_frame[16] [5]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[5]), .O(n59197));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1872.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1873 (.I0(\data_in_frame[16] [4]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[4]), .O(n59201));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1873.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1874 (.I0(\data_in_frame[16] [3]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[3]), .O(n59203));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1874.LUT_INIT = 16'h3a0a;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5750));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5749));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n30080), .O(n55993));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5748));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5747));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5746));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5745));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5744));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n59923));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n59922));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h4500;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5743));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5742));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5741));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n59921));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h4500;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5740));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5739));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13818_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n59773), 
            .I3(GND_net), .O(n32009));   // verilog/coms.v(130[12] 305[6])
    defparam i13818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n59933));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n59920));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n59919));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n59918));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n59917));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n59916));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h4500;
    SB_LUT4 i48716_2_lut (.I0(n71628), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67794));
    defparam i48716_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n59915));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n59914));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n59913));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n59912));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n59911));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n59934));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n60050));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h4500;
    SB_LUT4 i2_2_lut (.I0(hall2), .I1(commutation_state_7__N_27[2]), .I2(GND_net), 
            .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n60049));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n60048));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h4500;
    SB_LUT4 i1_3_lut_adj_1893 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1893.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n60047));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n59910));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h4500;
    SB_LUT4 i51696_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5869));
    defparam i51696_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n60046));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n59932));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h4500;
    SB_LUT4 i5_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n60045));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h4500;
    SB_LUT4 i12923_2_lut (.I0(n30015), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n31122));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i12923_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51422_4_lut (.I0(commutation_state[1]), .I1(n25253), .I2(dti), 
            .I3(commutation_state[2]), .O(n30015));
    defparam i51422_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n59909));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n59908));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n59907));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n59906));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n59905));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n59904));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n59903));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5848));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1331), .I3(n40695), .O(n24_adj_5856));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 mux_1677_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n10009));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n59902));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n11477));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n11475));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n11473));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n11471));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n11469));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n59901));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n59900));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n59899));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h4500;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[2]), .O(n63549));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_3_lut_4_lut_adj_1910 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_Bit_Index[0]), .O(n63621));
    defparam i1_3_lut_4_lut_adj_1910.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n31492));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n11467));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n11465));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n11463));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n59898));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n11461));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n60044));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n31490));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n11459));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n11457));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n11455));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n59897));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n11453));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n59896));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1917 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n60043));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1917.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n11451));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13196_4_lut (.I0(n30093), .I1(n1331), .I2(n67604), .I3(n40795), 
            .O(n31358));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i13196_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n60042));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n11449));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n60041));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n60040));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n60039));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n11447));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n60038));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n11445));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n60037));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n11443));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n11441));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n11439));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i41511_3_lut (.I0(n4_adj_5867), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n60952));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i41511_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n59936));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h4500;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n62946));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n60036));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h4500;
    SB_LUT4 i13626_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n31817));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n60035));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h4500;
    SB_LUT4 i13628_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n31819));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13628_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 LessThan_1178_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5839));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1800(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .n1757(n1757), 
            .GND_net(GND_net), .n1759(n1759), .n1761(n1761), .n1763(n1763), 
            .n1765(n1765), .n1767(n1767), .n1769(n1769), .n1771(n1771), 
            .n1773(n1773), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net), .\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), 
            .n31820(n31820), .n1755(n1755), .n31819(n31819), .a_prev(a_prev), 
            .n31817(n31817), .b_prev(b_prev), .position_31__N_3836(position_31__N_3836), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 i48363_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n67858));   // verilog/uart_rx.v(119[17:57])
    defparam i48363_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_3_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n35072), .I3(GND_net), .O(n25082));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i13630_3_lut (.I0(a_prev_adj_5788), .I1(a_new_adj_5905[1]), 
            .I2(debounce_cnt_N_3833_adj_5790), .I3(GND_net), .O(n31821));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n60034));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n60033));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n60032));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n60031));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1931 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n59895));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1931.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n59894));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n59893));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n31484));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n59892));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n59891));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n59890));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n59889));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h4500;
    SB_LUT4 i13515_3_lut_4_lut (.I0(n1805), .I1(b_prev_adj_5789), .I2(a_new_adj_5905[1]), 
            .I3(position_31__N_3836_adj_5791), .O(n31706));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13515_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i13514_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5942[1]), 
            .I2(r_SM_Main_adj_5942[2]), .I3(n6_adj_5849), .O(n31705));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13514_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n60030));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n60029));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1941 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n59888));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1941.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_3_lut_adj_1942 (.I0(hall1), .I1(hall2), .I2(n24006), 
            .I3(GND_net), .O(n4_adj_5867));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_1942.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n59887));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n59886));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n60028));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n59885));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n31475));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n31474));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n59884));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n59883));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n31471));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n31470));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n59882));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n59881));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h4500;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5952[0]), .I1(n67782), .I2(n6720), 
            .I3(n10_adj_5782), .O(n8_adj_5866));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n40695), .O(n58351));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 i13665_3_lut (.I0(current[11]), .I1(data_adj_5926[11]), .I2(n30062), 
            .I3(GND_net), .O(n31856));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13666_3_lut (.I0(current[10]), .I1(data_adj_5926[10]), .I2(n30062), 
            .I3(GND_net), .O(n31857));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n31467));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h4500;
    SB_LUT4 i13667_3_lut (.I0(current[9]), .I1(data_adj_5926[9]), .I2(n30062), 
            .I3(GND_net), .O(n31858));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13668_3_lut (.I0(current[8]), .I1(data_adj_5926[8]), .I2(n30062), 
            .I3(GND_net), .O(n31859));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13669_3_lut (.I0(current[7]), .I1(data_adj_5926[7]), .I2(n30062), 
            .I3(GND_net), .O(n31860));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13670_3_lut (.I0(current[6]), .I1(data_adj_5926[6]), .I2(n30062), 
            .I3(GND_net), .O(n31861));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n59880));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h4500;
    SB_LUT4 i13671_3_lut (.I0(current[5]), .I1(data_adj_5926[5]), .I2(n30062), 
            .I3(GND_net), .O(n31862));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13672_3_lut (.I0(current[4]), .I1(data_adj_5926[4]), .I2(n30062), 
            .I3(GND_net), .O(n31863));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n59879));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h4500;
    SB_LUT4 i13673_3_lut (.I0(current[3]), .I1(data_adj_5926[3]), .I2(n30062), 
            .I3(GND_net), .O(n31864));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5562_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5562_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i13674_3_lut (.I0(current[2]), .I1(data_adj_5926[2]), .I2(n30062), 
            .I3(GND_net), .O(n31865));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n59878));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h4500;
    SB_LUT4 i13675_3_lut (.I0(current[1]), .I1(data_adj_5926[1]), .I2(n30062), 
            .I3(GND_net), .O(n31866));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n60027));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h4500;
    SB_LUT4 i13676_3_lut (.I0(baudrate[31]), .I1(data_adj_5919[7]), .I2(n30137), 
            .I3(GND_net), .O(n31867));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n59873));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h4500;
    SB_LUT4 i13677_3_lut (.I0(baudrate[30]), .I1(data_adj_5919[6]), .I2(n30137), 
            .I3(GND_net), .O(n31868));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n59877));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n31461));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h4500;
    SB_LUT4 i5560_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5560_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i13678_3_lut (.I0(baudrate[29]), .I1(data_adj_5919[5]), .I2(n30137), 
            .I3(GND_net), .O(n31869));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n31460));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h4500;
    SB_LUT4 i13679_3_lut (.I0(baudrate[28]), .I1(data_adj_5919[4]), .I2(n30137), 
            .I3(GND_net), .O(n31870));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13680_3_lut (.I0(baudrate[27]), .I1(data_adj_5919[3]), .I2(n30137), 
            .I3(GND_net), .O(n31871));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n59876));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h4500;
    SB_LUT4 i13681_3_lut (.I0(baudrate[26]), .I1(data_adj_5919[2]), .I2(n30137), 
            .I3(GND_net), .O(n31872));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n59875));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h4500;
    SB_LUT4 i13682_3_lut (.I0(baudrate[25]), .I1(data_adj_5919[1]), .I2(n30137), 
            .I3(GND_net), .O(n31873));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n60026));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n60025));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h4500;
    SB_LUT4 i13683_3_lut (.I0(baudrate[24]), .I1(data_adj_5919[0]), .I2(n30137), 
            .I3(GND_net), .O(n31874));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n60024));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n60023));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n60022));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n60021));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n60020));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n60019));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n60018));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n60017));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n60016));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n60015));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n60014));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n60013));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n60012));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n60011));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n60010));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n60009));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n60008));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n60007));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n60006));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n60005));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n60004));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n60003));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n60002));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n60001));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n60000));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n59999));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n59998));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n59997));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n59996));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n59995));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n59994));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n59993));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n59992));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n59991));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n59990));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n59989));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n59988));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n59987));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n59986));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h4500;
    SB_LUT4 n9946_bdd_4_lut_51815 (.I0(n9946), .I1(current[11]), .I2(duty[14]), 
            .I3(n9944), .O(n71313));
    defparam n9946_bdd_4_lut_51815.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n59985));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n59984));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n59983));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n59982));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n59981));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n59980));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n59979));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n59978));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n59977));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2016 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n59976));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2016.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n59975));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2018 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n59974));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2018.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n59973));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h4500;
    SB_LUT4 i13715_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3178), .I3(GND_net), 
            .O(n31906));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2020 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n59972));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2020.LUT_INIT = 16'h4500;
    SB_LUT4 i13716_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3178), .I3(GND_net), 
            .O(n31907));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n60051));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h4500;
    SB_LUT4 i13717_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3178), .I3(GND_net), 
            .O(n31908));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n59971));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2023 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n59970));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2023.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n59935));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h4500;
    SB_LUT4 i13718_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3178), .I3(GND_net), 
            .O(n31909));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n59969));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h4500;
    SB_LUT4 i13719_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3178), .I3(GND_net), 
            .O(n31910));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2026 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n59968));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2026.LUT_INIT = 16'h4500;
    SB_LUT4 i13720_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3178), .I3(GND_net), 
            .O(n31911));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n59967));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h4500;
    SB_LUT4 i48719_2_lut_3_lut (.I0(n3489), .I1(n89), .I2(n76), .I3(GND_net), 
            .O(n67701));
    defparam i48719_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 n71313_bdd_4_lut (.I0(n71313), .I1(duty[11]), .I2(n4932), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[11]));
    defparam n71313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13721_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3178), .I3(GND_net), 
            .O(n31912));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n59966));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h4500;
    SB_LUT4 i48720_2_lut_3_lut (.I0(n3489), .I1(n89), .I2(n65), .I3(GND_net), 
            .O(n67697));
    defparam i48720_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i13722_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3178), .I3(GND_net), 
            .O(n31913));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n59965));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n59964));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h4500;
    SB_LUT4 i13723_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3178), .I3(GND_net), 
            .O(n31914));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n59963));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n59962));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n59961));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2034 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n59960));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2034.LUT_INIT = 16'h4500;
    SB_LUT4 i13724_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3178), .I3(GND_net), 
            .O(n31915));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2035 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n59959));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2035.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2036 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n59958));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2036.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2037 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n59957));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2037.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n59956));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n59955));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n59954));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2041 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n59953));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2041.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n59952));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n59951));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n59950));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n59949));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n59948));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n59947));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2048 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n59946));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2048.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2049 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n59874));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2049.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2050 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n59945));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2050.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n59944));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2052 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n59943));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2052.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n59942));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2054 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n59941));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2054.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n59940));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n59939));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n59938));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n59937));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h4500;
    SB_LUT4 mux_1677_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n11437));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n11435));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n59930));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h4500;
    SB_LUT4 i13964_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n59779), .I3(GND_net), .O(n32155));   // verilog/coms.v(130[12] 305[6])
    defparam i13964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9946_bdd_4_lut_51796 (.I0(n9946), .I1(current[4]), .I2(duty[7]), 
            .I3(n9944), .O(n71307));
    defparam n9946_bdd_4_lut_51796.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2060 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n59929));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2060.LUT_INIT = 16'h4500;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n59928));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h4500;
    SB_LUT4 i45215_3_lut (.I0(n4923), .I1(duty[20]), .I2(n9946), .I3(GND_net), 
            .O(n64710));
    defparam i45215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45217_3_lut (.I0(n64710), .I1(n64705), .I2(n9944), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i45217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45212_3_lut (.I0(n4922), .I1(duty[21]), .I2(n9946), .I3(GND_net), 
            .O(n64707));
    defparam i45212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45214_3_lut (.I0(n64707), .I1(n64705), .I2(n9944), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i45214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45210_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n9946), 
            .I3(GND_net), .O(n64705));
    defparam i45210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45209_3_lut (.I0(n4921), .I1(duty[22]), .I2(n9946), .I3(GND_net), 
            .O(n64704));
    defparam i45209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45211_3_lut (.I0(n64704), .I1(n64705), .I2(n9944), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i45211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_2062 (.I0(dti_counter[2]), .I1(dti_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5853));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut_adj_2062.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_2063 (.I0(dti_counter[6]), .I1(dti_counter[7]), 
            .I2(dti_counter[1]), .I3(dti_counter[5]), .O(n14_adj_5852));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_2063.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_2064 (.I0(dti_counter[0]), .I1(n14_adj_5852), .I2(n10_adj_5853), 
            .I3(dti_counter[3]), .O(n25253));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_2064.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2065 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5864));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2065.LUT_INIT = 16'h7bde;
    SB_LUT4 n71307_bdd_4_lut (.I0(n71307), .I1(duty[4]), .I2(n4939), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n71307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n59927));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h4500;
    SB_LUT4 i2_3_lut_adj_2067 (.I0(commutation_state[0]), .I1(n4_adj_5864), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5778));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut_adj_2067.LUT_INIT = 16'hdede;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n59926));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h4500;
    SB_LUT4 i51662_2_lut (.I0(n25253), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i51662_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i13967_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n59779), .I3(GND_net), .O(n32158));   // verilog/coms.v(130[12] 305[6])
    defparam i13967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13602_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n30673), 
            .I3(GND_net), .O(n31793));   // verilog/coms.v(130[12] 305[6])
    defparam i13602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13971_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n59779), .I3(GND_net), .O(n32162));   // verilog/coms.v(130[12] 305[6])
    defparam i13971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9946_bdd_4_lut_51791 (.I0(n9946), .I1(current[10]), .I2(duty[13]), 
            .I3(n9944), .O(n71301));
    defparam n9946_bdd_4_lut_51791.LUT_INIT = 16'he4aa;
    SB_LUT4 i13974_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n59779), .I3(GND_net), .O(n32165));   // verilog/coms.v(130[12] 305[6])
    defparam i13974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13977_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n59779), .I3(GND_net), .O(n32168));   // verilog/coms.v(130[12] 305[6])
    defparam i13977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13980_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n59779), .I3(GND_net), .O(n32171));   // verilog/coms.v(130[12] 305[6])
    defparam i13980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n71301_bdd_4_lut (.I0(n71301), .I1(duty[10]), .I2(n4933), 
            .I3(n9944), .O(pwm_setpoint_23__N_3[10]));
    defparam n71301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5774));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5776));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5772));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_4_lut_adj_2069 (.I0(n260), .I1(n64491), .I2(duty[23]), 
            .I3(n22_adj_5859), .O(n9944));
    defparam i1_4_lut_4_lut_adj_2069.LUT_INIT = 16'h1505;
    SB_LUT4 i49017_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n68512));
    defparam i49017_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n9946_bdd_4_lut_51786 (.I0(n9946), .I1(current[3]), .I2(duty[6]), 
            .I3(n9944), .O(n71295));
    defparam n9946_bdd_4_lut_51786.LUT_INIT = 16'he4aa;
    SB_LUT4 n71295_bdd_4_lut (.I0(n71295), .I1(duty[3]), .I2(n4940), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n71295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_2070 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(n55567), .I3(\data_out_frame[18] [5]), .O(n55781));
    defparam i2_3_lut_4_lut_adj_2070.LUT_INIT = 16'h6996;
    SB_LUT4 i45315_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64810));
    defparam i45315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45316_4_lut (.I0(n64810), .I1(n30323), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64811));
    defparam i45316_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45314_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64809));
    defparam i45314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_2071 (.I0(n8), .I1(n39602), .I2(GND_net), .I3(GND_net), 
            .O(n30629));
    defparam i1_2_lut_adj_2071.LUT_INIT = 16'hbbbb;
    SB_LUT4 i48699_2_lut (.I0(n71574), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67793));
    defparam i48699_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_2072 (.I0(\data_in_frame[16] [2]), .I1(n30629), 
            .I2(n30698), .I3(rx_data[2]), .O(n59095));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2072.LUT_INIT = 16'h3a0a;
    SB_LUT4 i45321_3_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n64816));
    defparam i45321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45320_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[6] [7]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n64815));
    defparam i45320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45322_4_lut (.I0(n64816), .I1(n30278), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64817));
    defparam i45322_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48379_3_lut_4_lut (.I0(r_Clock_Count_adj_5943[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5943[2]), .O(n67874));   // verilog/uart_tx.v(117[17:57])
    defparam i48379_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1181_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5943[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5831));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 n9946_bdd_4_lut_51781 (.I0(n9946), .I1(current[9]), .I2(duty[12]), 
            .I3(n9944), .O(n71265));
    defparam n9946_bdd_4_lut_51781.LUT_INIT = 16'he4aa;
    SB_LUT4 n71265_bdd_4_lut (.I0(n71265), .I1(duty[9]), .I2(n4934), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n71265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9946_bdd_4_lut_51757 (.I0(n9946), .I1(current[2]), .I2(duty[5]), 
            .I3(n9944), .O(n71253));
    defparam n9946_bdd_4_lut_51757.LUT_INIT = 16'he4aa;
    SB_LUT4 n71253_bdd_4_lut (.I0(n71253), .I1(duty[2]), .I2(n4941), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n71253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9946_bdd_4_lut_51748 (.I0(n9946), .I1(current[8]), .I2(duty[11]), 
            .I3(n9944), .O(n71229));
    defparam n9946_bdd_4_lut_51748.LUT_INIT = 16'he4aa;
    SB_LUT4 n71229_bdd_4_lut (.I0(n71229), .I1(duty[8]), .I2(n4935), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n71229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_14_i21_2_lut (.I0(current[10]), .I1(current_limit[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5756));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9946_bdd_4_lut_51728 (.I0(n9946), .I1(current[7]), .I2(duty[10]), 
            .I3(n9944), .O(n71223));
    defparam n9946_bdd_4_lut_51728.LUT_INIT = 16'he4aa;
    SB_LUT4 n71223_bdd_4_lut (.I0(n71223), .I1(duty[7]), .I2(n4936), .I3(n9944), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n71223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5759));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n64578), .I2(n64579), .I3(byte_transmit_counter[1]), .O(n71217));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71217_bdd_4_lut (.I0(n71217), .I1(n64882), .I2(n64881), .I3(byte_transmit_counter[1]), 
            .O(n71220));
    defparam n71217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[1]), .I3(neopxl_color[3]), .O(n71655));
    defparam color_bit_N_502_1__bdd_4_lut_4_lut.LUT_INIT = 16'he6a2;
    SB_LUT4 i51426_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[4] [3]), .I2(n30673), 
            .I3(GND_net), .O(n59473));   // verilog/coms.v(94[13:20])
    defparam i51426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_91[7]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_91[8]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5757));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    TLI4970 tli (.clk16MHz(clk16MHz), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n30062(n30062), .\current[15] (current[15]), .n31866(n31866), 
            .\current[1] (current[1]), .n31865(n31865), .\current[2] (current[2]), 
            .n31864(n31864), .\current[3] (current[3]), .n31863(n31863), 
            .\current[4] (current[4]), .n31862(n31862), .\current[5] (current[5]), 
            .n31861(n31861), .\current[6] (current[6]), .n31860(n31860), 
            .\current[7] (current[7]), .n31859(n31859), .\current[8] (current[8]), 
            .n31858(n31858), .\current[9] (current[9]), .n31857(n31857), 
            .\current[10] (current[10]), .n31856(n31856), .\current[11] (current[11]), 
            .\data[15] (data_adj_5926[15]), .\data[12] (data_adj_5926[12]), 
            .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .n32677(n32677), .n32676(n32676), 
            .n32675(n32675), .\data[11] (data_adj_5926[11]), .n32674(n32674), 
            .\data[10] (data_adj_5926[10]), .n32673(n32673), .\data[9] (data_adj_5926[9]), 
            .n32672(n32672), .\data[8] (data_adj_5926[8]), .n32671(n32671), 
            .\data[7] (data_adj_5926[7]), .n32670(n32670), .\data[6] (data_adj_5926[6]), 
            .n32669(n32669), .\data[5] (data_adj_5926[5]), .n32668(n32668), 
            .\data[4] (data_adj_5926[4]), .n32667(n32667), .\data[3] (data_adj_5926[3]), 
            .n32666(n32666), .\data[2] (data_adj_5926[2]), .n32665(n32665), 
            .\data[1] (data_adj_5926[1]), .n32299(n32299), .\data[0] (data_adj_5926[0]), 
            .n31699(n31699), .\current[0] (current[0]), .n27916(n27916), 
            .n27891(n27891), .n11(n11_adj_5784), .n27938(n27938), .n5(n5_adj_5783), 
            .n5_adj_25(n5_adj_5809), .n40832(n40832), .n27925(n27925), 
            .n5_adj_26(n5_adj_5797), .state_7__N_4319(state_7__N_4319)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(406[11] 412[4])
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(325[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_2073 (.I0(\data_out_frame[24] [3]), .I1(n55267), 
            .I2(n60414), .I3(n55802), .O(n60514));
    defparam i1_2_lut_4_lut_adj_2073.LUT_INIT = 16'h9669;
    SB_LUT4 i14008_3_lut (.I0(\data_in_frame[16] [0]), .I1(rx_data[0]), 
            .I2(n30698), .I3(GND_net), .O(n32199));   // verilog/coms.v(130[12] 305[6])
    defparam i14008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13837_4_lut_4_lut (.I0(n30217), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n32028));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13837_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5758));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5752), .I3(n15_adj_5808), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_91[9]), 
            .I2(n15_adj_5785), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5762));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i50601_3_lut (.I0(n4_adj_5762), .I1(current_limit[2]), .I2(current[2]), 
            .I3(GND_net), .O(n70096));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i50601_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_2074 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n60609));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_2074.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_2075 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(Kp_23__N_869), .I3(Kp_23__N_715), .O(n60538));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_2075.LUT_INIT = 16'h6996;
    SB_LUT4 i50602_3_lut (.I0(n70096), .I1(current_limit[3]), .I2(current[3]), 
            .I3(GND_net), .O(n37892));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i50602_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_2076 (.I0(state[0]), .I1(bit_ctr[3]), .I2(n40859), 
            .I3(bit_ctr[4]), .O(n4_adj_5844));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_4_lut_adj_2076.LUT_INIT = 16'hd555;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1800(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .\a_new[1] (a_new_adj_5905[1]), 
            .encoder1_position({encoder1_position}), .GND_net(GND_net), 
            .\b_new[1] (b_new_adj_5906[1]), .b_prev(b_prev_adj_5789), .VCC_net(VCC_net), 
            .n31821(n31821), .a_prev(a_prev_adj_5788), .position_31__N_3836(position_31__N_3836_adj_5791), 
            .n31707(n31707), .n31706(n31706), .n1805(n1805), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5790)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i1_4_lut_4_lut_adj_2077 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2834), .O(n25_adj_5855));   // verilog/TinyFPGA_B.v(378[7:11])
    defparam i1_4_lut_4_lut_adj_2077.LUT_INIT = 16'h5450;
    coms neopxl_color_23__I_0 (.reset(reset), .rx_data({rx_data}), .\data_in_frame[6] ({\data_in_frame[6] [7], 
         Open_2, Open_3, Open_4, \data_in_frame[6] [3:0]}), .n2887(n2887), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .clk16MHz(clk16MHz), 
         .n59931(n59931), .n59925(n59925), .n59095(n59095), .VCC_net(VCC_net), 
         .\data_in_frame[16] ({\data_in_frame[16] }), .n59924(n59924), .n32202(n32202), 
         .n59923(n59923), .n59922(n59922), .n59921(n59921), .n59933(n59933), 
         .n59920(n59920), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n59919(n59919), .n59918(n59918), .n59917(n59917), .n59916(n59916), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .n59915(n59915), .n59914(n59914), 
         .n59913(n59913), .n59912(n59912), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n59911(n59911), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n59934(n59934), .n32199(n32199), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n60050(n60050), .n59473(n59473), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n60049(n60049), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n60048(n60048), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n60047(n60047), .n59910(n59910), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n60046(n60046), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n59932(n59932), .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .byte_transmit_counter({Open_5, Open_6, Open_7, byte_transmit_counter[4:0]}), 
         .GND_net(GND_net), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[1][6] (\data_out_frame[1] [6]), 
         .n60045(n60045), .n59909(n59909), .n59908(n59908), .n59907(n59907), 
         .n59906(n59906), .n59905(n59905), .n59904(n59904), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n59903(n59903), .n59902(n59902), .n59901(n59901), .n59900(n59900), 
         .n59899(n59899), .n31492(n31492), .n59898(n59898), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n60044(n60044), .n31490(n31490), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .n59897(n59897), .n59896(n59896), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n60043(n60043), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n67793(n67793), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .n60042(n60042), .\data_in_frame[2] ({\data_in_frame[2] [7:1], 
         Open_8}), .deadband({deadband}), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .IntegralLimit({IntegralLimit}), .\data_in_frame[3] ({Open_9, Open_10, 
         Open_11, Open_12, Open_13, Open_14, Open_15, \data_in_frame[3] [0]}), 
         .\Kp[0] (Kp[0]), .\data_in_frame[5] ({\data_in_frame[5] }), .\Ki[0] (Ki[0]), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .PWMLimit({PWMLimit}), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .n60041(n60041), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n60040(n60040), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n60039(n60039), 
         .n60038(n60038), .n60037(n60037), .n59936(n59936), .n60036(n60036), 
         .n60035(n60035), .n60034(n60034), .n32171(n32171), .\data_in_frame[14] ({\data_in_frame[14] }), 
         .n60033(n60033), .n32168(n32168), .n60032(n60032), .n32165(n32165), 
         .n60031(n60031), .n59895(n59895), .n59894(n59894), .n59893(n59893), 
         .n31484(n31484), .n59892(n59892), .n59891(n59891), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .n59890(n59890), .n59889(n59889), .n32162(n32162), .n60030(n60030), 
         .n31793(n31793), .n60029(n60029), .n32158(n32158), .n59888(n59888), 
         .n59887(n59887), .n59886(n59886), .n60028(n60028), .n59885(n59885), 
         .n31475(n31475), .n31474(n31474), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n59884(n59884), .n59883(n59883), .n31471(n31471), .n31470(n31470), 
         .n32155(n32155), .n59882(n59882), .n59881(n59881), .n31467(n31467), 
         .n59880(n59880), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n59879(n59879), .n59878(n59878), .n60027(n60027), .n59873(n59873), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .n59877(n59877), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n31461(n31461), 
         .n60134(n60134), .n32152(n32152), .n31460(n31460), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n59876(n59876), .n59875(n59875), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n60514(n60514), .\data_out_frame[26] ({\data_out_frame[26] }), 
         .n60082(n60082), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .n32149(n32149), 
         .n60026(n60026), .LED_c(LED_c), .n60081(n60081), .\Ki[15] (Ki[15]), 
         .\FRAME_MATCHER.i_31__N_2513 (\FRAME_MATCHER.i_31__N_2513 ), .n35072(n35072), 
         .n31455(n31455), .\Ki[14] (Ki[14]), .\Ki[13] (Ki[13]), .setpoint({setpoint}), 
         .\Ki[12] (Ki[12]), .n32146(n32146), .n60080(n60080), .n60076(n60076), 
         .\Ki[11] (Ki[11]), .n60077(n60077), .\Ki[10] (Ki[10]), .n31451(n31451), 
         .\Ki[9] (Ki[9]), .n64802(n64802), .\Ki[8] (Ki[8]), .\Ki[7] (Ki[7]), 
         .n60075(n60075), .n60025(n60025), .\data_out_frame[27] ({\data_out_frame[27] }), 
         .n60072(n60072), .\Ki[6] (Ki[6]), .n60073(n60073), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .\encoder0_position_scaled[21] (encoder0_position_scaled[21]), .n31447(n31447), 
         .n32143(n32143), .n60078(n60078), .n60079(n60079), .n32140(n32140), 
         .\Ki[5] (Ki[5]), .\Ki[4] (Ki[4]), .\Ki[3] (Ki[3]), .\Ki[2] (Ki[2]), 
         .n60071(n60071), .n55748(n55748), .\Ki[1] (Ki[1]), .\Kp[15] (Kp[15]), 
         .n60024(n60024), .n55746(n55746), .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), 
         .\Kp[14] (Kp[14]), .n31443(n31443), .n60074(n60074), .n60414(n60414), 
         .n55760(n55760), .n60523(n60523), .\Kp[13] (Kp[13]), .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), 
         .\Kp[12] (Kp[12]), .\Kp[11] (Kp[11]), .n55781(n55781), .n32137(n32137), 
         .\Kp[10] (Kp[10]), .n32134(n32134), .n60150(n60150), .n31796(n31796), 
         .n60023(n60023), .n32130(n32130), .n32127(n32127), .n32124(n32124), 
         .n55267(n55267), .n55737(n55737), .\Kp[9] (Kp[9]), .n60022(n60022), 
         .\Kp[8] (Kp[8]), .n60021(n60021), .\Kp[7] (Kp[7]), .\Kp[6] (Kp[6]), 
         .n71628(n71628), .\data_out_frame[8][2] (\data_out_frame[8] [2]), 
         .\FRAME_MATCHER.i[2] (\FRAME_MATCHER.i [2]), .\FRAME_MATCHER.i[1] (\FRAME_MATCHER.i [1]), 
         .\data_in_frame[3][5] (\data_in_frame[3] [5]), .\Kp[5] (Kp[5]), 
         .\data_in_frame[21][7] (\data_in_frame[21] [7]), .\data_in_frame[17] ({\data_in_frame[17] [7], 
         Open_16, \data_in_frame[17] [5], Open_17, Open_18, Open_19, 
         Open_20, Open_21}), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .\data_in_frame[18] ({Open_22, \data_in_frame[18] [6], Open_23, 
         Open_24, Open_25, \data_in_frame[18] [2], Open_26, Open_27}), 
         .\data_in_frame[21][1] (\data_in_frame[21] [1]), .\data_in_frame[21][2] (\data_in_frame[21] [2]), 
         .\data_in_frame[21][4] (\data_in_frame[21] [4]), .\data_in_frame[21][0] (\data_in_frame[21] [0]), 
         .\data_in_frame[18][7] (\data_in_frame[18] [7]), .\Kp[4] (Kp[4]), 
         .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .\data_in_frame[21][3] (\data_in_frame[21] [3]), 
         .n31802(n31802), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .\Kp[3] (Kp[3]), .\Kp[2] (Kp[2]), .\Kp[1] (Kp[1]), .n60020(n60020), 
         .\data_in_frame[18][1] (\data_in_frame[18] [1]), .\data_in_frame[18][3] (\data_in_frame[18] [3]), 
         .n60019(n60019), .n32068(n32068), .n32065(n32065), .n32062(n32062), 
         .n60018(n60018), .n71574(n71574), .control_mode({Open_28, Open_29, 
         control_mode[5:4], Open_30, Open_31, Open_32, Open_33}), 
         .n62692(n62692), .n30673(n30673), .n32059(n32059), .n32056(n32056), 
         .n32053(n32053), .n32050(n32050), .n32047(n32047), .n32044(n32044), 
         .n32041(n32041), .n32038(n32038), .n31806(n31806), .\control_mode[6] (control_mode[6]), 
         .\control_mode[7] (control_mode[7]), .n31811(n31811), .n31853(n31853), 
         .n31916(n31916), .n31919(n31919), .n31922(n31922), .n31925(n31925), 
         .n32018(n32018), .n32015(n32015), .n60609(n60609), .n32012(n32012), 
         .n32009(n32009), .n32005(n32005), .n60017(n60017), .\data_in_frame[6][6] (\data_in_frame[6] [6]), 
         .\data_in_frame[17][6] (\data_in_frame[17] [6]), .\data_in_frame[18][0] (\data_in_frame[18] [0]), 
         .DE_c(DE_c), .n60016(n60016), .n60015(n60015), .n60014(n60014), 
         .n60013(n60013), .n60012(n60012), .n60011(n60011), .n60010(n60010), 
         .n60009(n60009), .n60008(n60008), .\data_out_frame[8][1] (\data_out_frame[8] [1]), 
         .n60007(n60007), .n60006(n60006), .\data_out_frame[8][3] (\data_out_frame[8] [3]), 
         .n60005(n60005), .\data_out_frame[8][4] (\data_out_frame[8] [4]), 
         .n60004(n60004), .\data_out_frame[8][5] (\data_out_frame[8] [5]), 
         .n60003(n60003), .\data_out_frame[8][6] (\data_out_frame[8] [6]), 
         .n60002(n60002), .\data_out_frame[8][7] (\data_out_frame[8] [7]), 
         .n60001(n60001), .n60000(n60000), .n59999(n59999), .n59998(n59998), 
         .n59997(n59997), .n59996(n59996), .n59995(n59995), .n59994(n59994), 
         .n59993(n59993), .n59992(n59992), .n59991(n59991), .n59990(n59990), 
         .n59989(n59989), .n59988(n59988), .n59987(n59987), .n59986(n59986), 
         .n59985(n59985), .n59984(n59984), .n59983(n59983), .n59982(n59982), 
         .n59981(n59981), .n59980(n59980), .n59979(n59979), .n59978(n59978), 
         .n59977(n59977), .n59976(n59976), .n59975(n59975), .n59974(n59974), 
         .n59973(n59973), .n59972(n59972), .n60051(n60051), .n59971(n59971), 
         .n59970(n59970), .n59935(n59935), .n59969(n59969), .n59968(n59968), 
         .n59967(n59967), .n59966(n59966), .n59965(n59965), .n59964(n59964), 
         .n59963(n59963), .n59962(n59962), .n59961(n59961), .n59960(n59960), 
         .n59959(n59959), .n59958(n59958), .n59957(n59957), .n59956(n59956), 
         .n59955(n59955), .n59954(n59954), .n59953(n59953), .n59952(n59952), 
         .n59951(n59951), .n59950(n59950), .n59949(n59949), .n59948(n59948), 
         .n59947(n59947), .n59946(n59946), .n59874(n59874), .n59945(n59945), 
         .n59944(n59944), .n59943(n59943), .n59942(n59942), .n59941(n59941), 
         .n59940(n59940), .n31818(n31818), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n59939(n59939), .n59938(n59938), .n59937(n59937), .n59930(n59930), 
         .displacement({displacement}), .n59929(n59929), .\data_in_frame[1] ({\data_in_frame[1] [7:4], 
         Open_34, Open_35, Open_36, Open_37}), .n59928(n59928), .\data_in_frame[22] ({Open_38, 
         \data_in_frame[22] [6], Open_39, \data_in_frame[22] [4], Open_40, 
         \data_in_frame[22] [2:1], Open_41}), .\data_in_frame[22][3] (\data_in_frame[22] [3]), 
         .\data_in_frame[22][7] (\data_in_frame[22] [7]), .Kp_23__N_715(Kp_23__N_715), 
         .n60538(n60538), .Kp_23__N_869(Kp_23__N_869), .n3489(n3489), 
         .n59927(n59927), .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), 
         .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), .n59203(n59203), 
         .n39602(n39602), .n61124(n61124), .n76(n76), .n59201(n59201), 
         .n59197(n59197), .n59193(n59193), .n59189(n59189), .n59315(n59315), 
         .n32704(n32704), .n59313(n59313), .n59185(n59185), .n59181(n59181), 
         .n59177(n59177), .n32290(n32290), .n32300(n32300), .\data_in_frame[18][5] (\data_in_frame[18] [5]), 
         .n59173(n59173), .n32306(n32306), .n32632(n32632), .n32363(n32363), 
         .n59263(n59263), .n59265(n59265), .n59255(n59255), .n59309(n59309), 
         .\data_in_frame[21][5] (\data_in_frame[21] [5]), .n32387(n32387), 
         .n32390(n32390), .n32393(n32393), .n32396(n32396), .n32403(n32403), 
         .\data_in_frame[22][5] (\data_in_frame[22] [5]), .n32406(n32406), 
         .n32409(n32409), .n31736(n31736), .n31739(n31739), .n31742(n31742), 
         .n32489(n32489), .neopxl_color({neopxl_color}), .n32488(n32488), 
         .n32487(n32487), .n32484(n32484), .n32483(n32483), .n32482(n32482), 
         .n32481(n32481), .n32480(n32480), .n32479(n32479), .n32478(n32478), 
         .n32477(n32477), .n32475(n32475), .n32474(n32474), .n32472(n32472), 
         .n32471(n32471), .n32470(n32470), .n32469(n32469), .n32468(n32468), 
         .n32467(n32467), .\control_mode[1] (control_mode[1]), .n31745(n31745), 
         .n32462(n32462), .n32461(n32461), .n32460(n32460), .n32459(n32459), 
         .n32458(n32458), .current_limit({current_limit}), .n32457(n32457), 
         .n37917(n37917), .n32455(n32455), .n30619(n30619), .n59926(n59926), 
         .n32454(n32454), .n32452(n32452), .n32451(n32451), .n32450(n32450), 
         .n32449(n32449), .n32448(n32448), .n32447(n32447), .n32446(n32446), 
         .n32445(n32445), .n32444(n32444), .n31748(n31748), .n31751(n31751), 
         .n31754(n31754), .n31757(n31757), .n67702(n67702), .n59777(n59777), 
         .n31766(n31766), .n31772(n31772), .n31695(n31695), .\control_mode[0] (control_mode[0]), 
         .n31693(n31693), .n31784(n31784), .n31787(n31787), .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), 
         .ID({ID}), .n55567(n55567), .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), 
         .n71580(n71580), .n55802(n55802), .n30671(n30671), .n25151(n25151), 
         .pwm_setpoint({pwm_setpoint}), .n25082(n25082), .n8(n8), .rx_data_ready(rx_data_ready), 
         .n65(n65), .n30627(n30627), .n59773(n59773), .n67698(n67698), 
         .n89(n89), .n30669(n30669), .tx_active(tx_active), .control_update(control_update), 
         .n30039(n30039), .n30709(n30709), .n30708(n30708), .n15(n15_adj_5808), 
         .n30702(n30702), .n15_adj_6(n15_adj_5785), .n15_adj_7(n15_adj_5752), 
         .\current[15] (current[15]), .n7(n7_adj_5847), .n64811(n64811), 
         .n64809(n64809), .n30700(n30700), .n59779(n59779), .n28460(n28460), 
         .encoder1_position_scaled({encoder1_position_scaled}), .n41236(n41236), 
         .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), 
         .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), 
         .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), .\encoder0_position_scaled[2] (encoder0_position_scaled[2]), 
         .\encoder0_position_scaled[1] (encoder0_position_scaled[1]), .n6(n6_adj_5861), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), 
         .n8_adj_8(n8_adj_5815), .n30621(n30621), .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), 
         .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), 
         .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), 
         .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), .\encoder0_position_scaled[23] (encoder0_position_scaled[23]), 
         .n39603(n39603), .\current[7] (current[7]), .\current[6] (current[6]), 
         .\current[5] (current[5]), .n30623(n30623), .\current[4] (current[4]), 
         .\current[3] (current[3]), .\current[2] (current[2]), .n59772(n59772), 
         .n30323(n30323), .\current[1] (current[1]), .n30278(n30278), 
         .n64817(n64817), .n64815(n64815), .\current[0] (current[0]), 
         .\current[11] (current[11]), .\current[10] (current[10]), .\current[9] (current[9]), 
         .\current[8] (current[8]), .n64584(n64584), .n64585(n64585), 
         .n64582(n64582), .n64581(n64581), .n1(n1), .tx_o(tx_o), .\tx_data[0] (tx_data[0]), 
         .r_SM_Main({r_SM_Main_adj_5942}), .\r_Bit_Index[0] (r_Bit_Index_adj_5944[0]), 
         .n59789(n59789), .n63279(n63279), .n27(n27), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
         .r_Clock_Count({r_Clock_Count_adj_5943}), .n32272(n32272), .n71737(n71737), 
         .n30087(n30087), .n31705(n31705), .n5233(n5233), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
         .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n29(n29), .n23(n23_adj_5860), 
         .n61776(n61776), .n6_adj_9(n6_adj_5849), .n60925(n60925), .n63255(n63255), 
         .tx_enable(tx_enable), .baudrate({baudrate}), .n27889(n27889), 
         .r_SM_Main_adj_23({r_SM_Main}), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
         .r_Clock_Count_adj_24({r_Clock_Count}), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .\r_Bit_Index[0]_adj_21 (r_Bit_Index[0]), 
         .n59798(n59798), .n63269(n63269), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .n5230(n5230), .n32278(n32278), 
         .n55993(n55993), .n30084(n30084), .n32606(n32606), .n32605(n32605), 
         .n32604(n32604), .n32603(n32603), .n32600(n32600), .n32599(n32599), 
         .n32598(n32598), .n32286(n32286), .n60086(n60086), .n4(n4_adj_5781), 
         .n6_adj_22(n6_adj_5865), .n30080(n30080), .n60927(n60927), .n63257(n63257), 
         .n63621(n63621), .n63605(n63605), .n63549(n63549), .n63515(n63515), 
         .n63551(n63551), .n63641(n63641), .n63587(n63587), .n63623(n63623)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i1956_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1331), .I3(n40695), .O(n6916));   // verilog/TinyFPGA_B.v(363[5] 389[12])
    defparam i1956_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2078 (.I0(n3489), .I1(n89), .I2(reset), 
            .I3(n65), .O(n30700));   // verilog/TinyFPGA_B.v(360[10] 390[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2078.LUT_INIT = 16'h0008;
    EEPROM eeprom (.clk16MHz(clk16MHz), .GND_net(GND_net), .\state_7__N_3918[0] (state_7__N_3918[0]), 
           .ID({ID}), .baudrate({baudrate}), .n31874(n31874), .n31873(n31873), 
           .n31872(n31872), .n31871(n31871), .n31870(n31870), .n31869(n31869), 
           .n31868(n31868), .n31867(n31867), .data_ready(data_ready), 
           .data({data_adj_5919}), .n30137(n30137), .scl_enable(scl_enable), 
           .VCC_net(VCC_net), .scl(scl), .sda_enable(sda_enable), .n32663(n32663), 
           .n32651(n32651), .n32650(n32650), .n32649(n32649), .n32645(n32645), 
           .n32644(n32644), .n32640(n32640), .n6720(n6720), .n32250(n32250), 
           .n8(n8_adj_5866), .\state[0] (state_adj_5952[0]), .\state_7__N_4126[3] (state_7__N_4126[3]), 
           .n4(n4_adj_5779), .n4_adj_4(n4_adj_5780), .n40902(n40902), 
           .sda_out(sda_out), .n10(n10_adj_5846), .n10_adj_5(n10_adj_5782), 
           .n27930(n27930), .n27881(n27881), .n67782(n67782)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(392[10] 404[6])
    pwm PWM (.pwm_setpoint({pwm_setpoint}), .GND_net(GND_net), .n2887(n2887), 
        .pwm_out(pwm_out), .clk32MHz(clk32MHz), .VCC_net(VCC_net), .reset(reset)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i13821_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n59773), 
            .I3(GND_net), .O(n32012));   // verilog/coms.v(130[12] 305[6])
    defparam i13821_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.\Ki[4] (Ki[4]), .n335({n336, n337, n338, 
            n339, n340, n341, n342, n343, n344, n345, n346, 
            n347, n348, n349, n350, n351, n352, n353, n354, 
            n355, n356, n357, n358, n359}), .GND_net(GND_net), .\Ki[5] (Ki[5]), 
            .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .setpoint({setpoint}), .motor_state({Open_42, 
            Open_43, Open_44, Open_45, Open_46, Open_47, Open_48, 
            Open_49, Open_50, Open_51, Open_52, Open_53, Open_54, 
            motor_state[10:1], Open_55}), .IntegralLimit({IntegralLimit}), 
            .\Ki[9] (Ki[9]), .\Kp[8] (Kp[8]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
            .\Ki[8] (Ki[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Ki[1] (Ki[1]), 
            .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Kp[11] (Kp[11]), 
            .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Ki[12] (Ki[12]), .\Kp[2] (Kp[2]), .\Ki[13] (Ki[13]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .\Kp[7] (Kp[7]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .VCC_net(VCC_net), .\Kp[14] (Kp[14]), 
            .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), .n32594(n32594), 
            .n32593(n32593), .n32592(n32592), .n32591(n32591), .n32590(n32590), 
            .n32589(n32589), .n32588(n32588), .n32587(n32587), .n32586(n32586), 
            .n32585(n32585), .n32584(n32584), .n32583(n32583), .n32582(n32582), 
            .n32581(n32581), .n32580(n32580), .n32579(n32579), .n32578(n32578), 
            .n32577(n32577), .n32576(n32576), .n32575(n32575), .n32574(n32574), 
            .n32573(n32573), .n32570(n32570), .n31682(n31682), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\encoder1_position_scaled[0] (encoder1_position_scaled[0]), .n15(n15_adj_5785), 
            .n67541(n67541), .n15_adj_1(n15_adj_5752), .\motor_state[20] (motor_state[20]), 
            .\motor_state[19] (motor_state[19]), .\motor_state[18] (motor_state[18]), 
            .\motor_state[17] (motor_state[17]), .\motor_state[16] (motor_state[16]), 
            .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .\motor_state[11] (motor_state[11]), .\Kp[15] (Kp[15]), .deadband({deadband}), 
            .PWMLimit({PWMLimit}), .n41195(n41195), .\control_mode[0] (control_mode[0]), 
            .\control_mode[7] (control_mode[7]), .\control_mode[6] (control_mode[6]), 
            .n62692(n62692), .\control_mode[1] (control_mode[1]), .n43(n43)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, n67418, GND_net, 
            bit_ctr, n40859, n54840, \color_bit_N_502[1] , n30217, 
            state, n27360, \neopxl_color[9] , \neopxl_color[8] , \neopxl_color[5] , 
            \neopxl_color[4] , timer, LED_c, VCC_net, n32028, n59083, 
            \bit_ctr[4] , n31915, t0, n31914, n31913, n31912, n31911, 
            n31910, n31909, n31908, n31907, n31906, NEOPXL_c, n31708, 
            \neopxl_color[14] , \neopxl_color[15] , \neopxl_color[12] , 
            \neopxl_color[13] , n71658, \neopxl_color[20] , \neopxl_color[22] , 
            \neopxl_color[21] , \neopxl_color[23] , \neopxl_color[17] , 
            \neopxl_color[19] , \neopxl_color[16] , \neopxl_color[18] , 
            n3178, \neopxl_color[6] , \neopxl_color[7] , \neopxl_color[10] , 
            \neopxl_color[11] ) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output n67418;
    input GND_net;
    output [4:0]bit_ctr;
    output n40859;
    output n54840;
    output \color_bit_N_502[1] ;
    output n30217;
    output [1:0]state;
    output n27360;
    input \neopxl_color[9] ;
    input \neopxl_color[8] ;
    input \neopxl_color[5] ;
    input \neopxl_color[4] ;
    output [10:0]timer;
    input LED_c;
    input VCC_net;
    input n32028;
    input n59083;
    output \bit_ctr[4] ;
    input n31915;
    output [10:0]t0;
    input n31914;
    input n31913;
    input n31912;
    input n31911;
    input n31910;
    input n31909;
    input n31908;
    input n31907;
    input n31906;
    output NEOPXL_c;
    input n31708;
    input \neopxl_color[14] ;
    input \neopxl_color[15] ;
    input \neopxl_color[12] ;
    input \neopxl_color[13] ;
    input n71658;
    input \neopxl_color[20] ;
    input \neopxl_color[22] ;
    input \neopxl_color[21] ;
    input \neopxl_color[23] ;
    input \neopxl_color[17] ;
    input \neopxl_color[19] ;
    input \neopxl_color[16] ;
    input \neopxl_color[18] ;
    output n3178;
    input \neopxl_color[6] ;
    input \neopxl_color[7] ;
    input \neopxl_color[10] ;
    input \neopxl_color[11] ;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n62573, \neo_pixel_transmitter.done , 
        start_N_507, n59349, start, n54873;
    wire [5:0]color_bit_N_502;
    
    wire n41254, n8, n81, n31647, n40798, n30029, n71619, n71622, 
        n71613, n71616, n30211;
    wire [10:0]n49;
    
    wire n53516, n53515, n53514, n53513, n53512, n53511, n53510, 
        n53509, n53508, n53507, n31129;
    wire [31:0]n149;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    
    wire n27859, n25041, n23410;
    wire [10:0]n1;
    
    wire n52994, n52993, n52992;
    wire [1:0]state_1__N_451;
    
    wire n31128, n52991, one_wire_N_499, n44, n62727, n52990, n52989, 
        n52988, n52987, n52986, n52985, n64395, n15, n27910, n27912, 
        n61151, n15_adj_5730, n62285, n61120, n32, n27907, n67416, 
        n61046, n62600, n22, n25, n7206, n67805, n68, n53_adj_5731, 
        n60093, n64825, n64824, n71262, n64826, n64780, n64779, 
        n64781, n64614, n64615, n64888, n64887, n40761, n61020, 
        n6_adj_5732, n67797, n67795, n71259, n6_adj_5733, n63023;
    
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n62573), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n59349), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i47923_2_lut (.I0(n54873), .I1(color_bit_N_502[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67418));
    defparam i47923_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[3]), .I1(n40859), .I2(GND_net), .I3(GND_net), 
            .O(n54840));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1174_4_lut (.I0(\color_bit_N_502[1] ), .I1(n41254), .I2(n8), 
            .I3(color_bit_N_502[2]), .O(n81));   // verilog/neopixel.v(24[26:38])
    defparam i1174_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i13456_2_lut (.I0(n30217), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n31647));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13456_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_4_lut (.I0(n27360), .I1(state[1]), .I2(n40798), .I3(state[0]), 
            .O(n30029));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hee2e;
    SB_LUT4 n71619_bdd_4_lut (.I0(n71619), .I1(\neopxl_color[9] ), .I2(\neopxl_color[8] ), 
            .I3(\color_bit_N_502[1] ), .O(n71622));
    defparam n71619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n71613_bdd_4_lut (.I0(n71613), .I1(\neopxl_color[5] ), .I2(\neopxl_color[4] ), 
            .I3(\color_bit_N_502[1] ), .O(n71616));
    defparam n71613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut (.I0(n27360), .I1(state[1]), .I2(n30211), .I3(GND_net), 
            .O(n30217));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2201_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));   // verilog/neopixel.v(65[23:32])
    defparam i2201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 timer_2039_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n53516), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2039_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n53515), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_11 (.CI(n53515), .I0(GND_net), .I1(timer[9]), 
            .CO(n53516));
    SB_LUT4 timer_2039_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n53514), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n30211));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_CARRY timer_2039_add_4_10 (.CI(n53514), .I0(GND_net), .I1(timer[8]), 
            .CO(n53515));
    SB_LUT4 timer_2039_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n53513), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_9 (.CI(n53513), .I0(GND_net), .I1(timer[7]), 
            .CO(n53514));
    SB_LUT4 timer_2039_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n53512), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_8 (.CI(n53512), .I0(GND_net), .I1(timer[6]), 
            .CO(n53513));
    SB_LUT4 timer_2039_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n53511), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_7 (.CI(n53511), .I0(GND_net), .I1(timer[5]), 
            .CO(n53512));
    SB_LUT4 timer_2039_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n53510), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_6 (.CI(n53510), .I0(GND_net), .I1(timer[4]), 
            .CO(n53511));
    SB_LUT4 timer_2039_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n53509), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_5 (.CI(n53509), .I0(GND_net), .I1(timer[3]), 
            .CO(n53510));
    SB_LUT4 timer_2039_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n53508), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_4 (.CI(n53508), .I0(GND_net), .I1(timer[2]), 
            .CO(n53509));
    SB_LUT4 timer_2039_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n53507), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_3 (.CI(n53507), .I0(GND_net), .I1(timer[1]), 
            .CO(n53508));
    SB_LUT4 timer_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n53507));
    SB_DFFE bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(VCC_net), .D(n32028));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i12938_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n31129));   // verilog/neopixel.v(35[4] 112[11])
    defparam i12938_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n59083));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2039__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n30217), 
            .D(n149[2]), .R(n31647));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr[3]), .C(clk16MHz), .E(n30217), .D(n149[3]), 
            .R(n31647));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n30217), 
            .D(n149[4]), .R(n31647));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n31915));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n31914));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n31913));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n31912));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n31911));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n31910));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n31909));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n31908));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n31907));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n31906));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i5573_3_lut_4_lut (.I0(start), .I1(n27859), .I2(n25041), .I3(bit_ctr[0]), 
            .O(n23410));
    defparam i5573_3_lut_4_lut.LUT_INIT = 16'hfb04;
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n52994), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n52993), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n52993), .I0(timer[9]), .I1(n1[9]), 
            .CO(n52994));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n52992), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n30211), .D(n23410), 
            .R(n31129));   // verilog/neopixel.v(34[12] 113[6])
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n52992), .I0(timer[8]), .I1(n1[8]), 
            .CO(n52993));
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n30029), .D(state_1__N_451[0]), 
            .S(n31128));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n52991), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n44), .D(one_wire_N_499), 
            .R(n62727));   // verilog/neopixel.v(34[12] 113[6])
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n52991), .I0(timer[7]), .I1(n1[7]), 
            .CO(n52992));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n52990), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1782 (.I0(start), .I1(n27859), .I2(n25041), 
            .I3(GND_net), .O(n27360));
    defparam i1_2_lut_3_lut_adj_1782.LUT_INIT = 16'h0404;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n52990), .I0(timer[6]), .I1(n1[6]), 
            .CO(n52991));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n52989), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n52989), .I0(timer[5]), .I1(n1[5]), 
            .CO(n52990));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n52988), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n52988), .I0(timer[4]), .I1(n1[4]), 
            .CO(n52989));
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n52987), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n52987), .I0(timer[3]), .I1(n1[3]), 
            .CO(n52988));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n52986), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n52986), .I0(timer[2]), .I1(n1[2]), 
            .CO(n52987));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n52985), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n52985), .I0(timer[1]), .I1(n1[1]), 
            .CO(n52986));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n52985));
    SB_LUT4 i1_2_lut_3_lut_adj_1783 (.I0(bit_ctr[3]), .I1(n40859), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n54873));
    defparam i1_2_lut_3_lut_adj_1783.LUT_INIT = 16'h7878;
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_LUT4 i23157_2_lut_3_lut (.I0(bit_ctr[3]), .I1(n40859), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n41254));
    defparam i23157_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_LUT4 i3_3_lut_4_lut (.I0(t1[0]), .I1(t1[4]), .I2(t1[2]), .I3(n64395), 
            .O(n15));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut (.I0(t1[0]), .I1(t1[4]), .I2(t1[3]), .I3(t1[1]), 
            .O(n27910));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1784 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n27912), .I3(state[1]), .O(n62727));
    defparam i2_3_lut_4_lut_adj_1784.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1785 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n61151), .I3(n15_adj_5730), .O(n62285));
    defparam i2_3_lut_4_lut_adj_1785.LUT_INIT = 16'hfffe;
    SB_LUT4 i41672_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n27912), .I3(GND_net), .O(n61120));
    defparam i41672_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n31708));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2039__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 i1_2_lut_3_lut_adj_1786 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1786.LUT_INIT = 16'h1e1e;
    SB_LUT4 i22767_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n40859));
    defparam i22767_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_4_lut_adj_1787 (.I0(n15), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(n15_adj_5730), .O(n32));
    defparam i1_4_lut_4_lut_adj_1787.LUT_INIT = 16'h14d7;
    SB_LUT4 i3_3_lut_4_lut_adj_1788 (.I0(t1[9]), .I1(t1[6]), .I2(t1[7]), 
            .I3(t1[5]), .O(n27907));   // verilog/neopixel.v(100[14:42])
    defparam i3_3_lut_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i6917_3_lut_4_lut (.I0(n15), .I1(t1[2]), .I2(n27910), .I3(state[0]), 
            .O(n25041));   // verilog/neopixel.v(35[4] 112[11])
    defparam i6917_3_lut_4_lut.LUT_INIT = 16'hf3aa;
    SB_LUT4 i2208_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2208_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i47921_2_lut_3_lut (.I0(n54873), .I1(bit_ctr[3]), .I2(n40859), 
            .I3(GND_net), .O(n67416));   // verilog/neopixel.v(24[26:38])
    defparam i47921_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i41600_2_lut_3_lut (.I0(n27912), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n61046));
    defparam i41600_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1789 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(t1[2]), .I3(n27910), .O(n62600));
    defparam i2_3_lut_4_lut_adj_1789.LUT_INIT = 16'h0080;
    SB_LUT4 i47_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n22));
    defparam i47_3_lut_4_lut_3_lut.LUT_INIT = 16'h8181;
    SB_LUT4 i46_3_lut_4_lut_3_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25));
    defparam i46_3_lut_4_lut_3_lut.LUT_INIT = 16'h1818;
    SB_LUT4 i2215_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(bit_ctr[3]), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2215_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i2222_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n7206), .I2(bit_ctr[3]), 
            .I3(\bit_ctr[4] ), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2222_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49300_3_lut (.I0(n27912), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n67805));
    defparam i49300_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i72_4_lut (.I0(n62285), .I1(n67805), .I2(state[1]), .I3(start), 
            .O(n68));
    defparam i72_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i51688_4_lut (.I0(n61151), .I1(n68), .I2(n62600), .I3(n53_adj_5731), 
            .O(n44));
    defparam i51688_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22706_2_lut (.I0(n27912), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n40798));
    defparam i22706_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(start), .I1(n61046), .I2(state[1]), .I3(n60093), 
            .O(n31128));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i45330_3_lut (.I0(\neopxl_color[14] ), .I1(\neopxl_color[15] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64825));
    defparam i45330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45329_3_lut (.I0(\neopxl_color[12] ), .I1(\neopxl_color[13] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n64824));
    defparam i45329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45331_4_lut (.I0(n64825), .I1(n71262), .I2(n54873), .I3(n54840), 
            .O(n64826));
    defparam i45331_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45285_4_lut (.I0(n64826), .I1(n64824), .I2(n54873), .I3(\color_bit_N_502[1] ), 
            .O(n64780));
    defparam i45285_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i45284_3_lut (.I0(n71658), .I1(n71616), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n64779));
    defparam i45284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45286_3_lut (.I0(n64780), .I1(n71622), .I2(n67418), .I3(GND_net), 
            .O(n64781));
    defparam i45286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22607_4_lut (.I0(n64781), .I1(n81), .I2(n64779), .I3(n67416), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i22607_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i45119_3_lut_4_lut (.I0(\neopxl_color[20] ), .I1(\neopxl_color[22] ), 
            .I2(bit_ctr[1]), .I3(bit_ctr[0]), .O(n64614));
    defparam i45119_3_lut_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i45120_3_lut_4_lut (.I0(\neopxl_color[21] ), .I1(\neopxl_color[23] ), 
            .I2(bit_ctr[1]), .I3(bit_ctr[0]), .O(n64615));
    defparam i45120_3_lut_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i45393_3_lut_4_lut (.I0(\neopxl_color[17] ), .I1(\neopxl_color[19] ), 
            .I2(bit_ctr[1]), .I3(bit_ctr[0]), .O(n64888));
    defparam i45393_3_lut_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i45392_3_lut_4_lut (.I0(\neopxl_color[16] ), .I1(\neopxl_color[18] ), 
            .I2(bit_ctr[1]), .I3(bit_ctr[0]), .O(n64887));
    defparam i45392_3_lut_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i22669_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n40761));
    defparam i22669_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41574_2_lut (.I0(t1[10]), .I1(t1[9]), .I2(GND_net), .I3(GND_net), 
            .O(n61020));
    defparam i41574_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i41703_4_lut (.I0(t1[8]), .I1(n61020), .I2(n6_adj_5732), .I3(t1[5]), 
            .O(n61151));
    defparam i41703_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49080_4_lut (.I0(n22), .I1(n25), .I2(n40761), .I3(state[0]), 
            .O(n67797));
    defparam i49080_4_lut.LUT_INIT = 16'h0c0a;
    SB_LUT4 i49728_4_lut (.I0(n67797), .I1(t1[4]), .I2(t1[2]), .I3(n61151), 
            .O(n67795));
    defparam i49728_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i45_3_lut (.I0(n67795), .I1(state[1]), .I2(start), .I3(GND_net), 
            .O(n3178));
    defparam i45_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2203_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n7206));   // verilog/neopixel.v(65[23:32])
    defparam i2203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 bit_ctr_0__bdd_4_lut_52048_4_lut (.I0(bit_ctr[0]), .I1(\neopxl_color[6] ), 
            .I2(\neopxl_color[7] ), .I3(bit_ctr[1]), .O(n71613));
    defparam bit_ctr_0__bdd_4_lut_52048_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(\neopxl_color[10] ), 
            .I2(\neopxl_color[11] ), .I3(bit_ctr[1]), .O(n71619));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_52043 (.I0(bit_ctr[0]), .I1(n64614), .I2(n64615), 
            .I3(color_bit_N_502[2]), .O(n71259));
    defparam bit_ctr_0__bdd_4_lut_52043.LUT_INIT = 16'he4aa;
    SB_LUT4 n71259_bdd_4_lut (.I0(n71259), .I1(n64888), .I2(n64887), .I3(color_bit_N_502[2]), 
            .O(n71262));
    defparam n71259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_4_lut_adj_1790 (.I0(bit_ctr[3]), .I1(n40859), .I2(n54873), 
            .I3(bit_ctr[0]), .O(n8));
    defparam i3_3_lut_4_lut_adj_1790.LUT_INIT = 16'hff9f;
    SB_LUT4 i3_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n27907), .I2(t1[10]), 
            .I3(t1[8]), .O(n27859));
    defparam i3_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_1791 (.I0(n25041), .I1(n27859), .I2(GND_net), 
            .I3(GND_net), .O(n60093));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_adj_1791.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1792 (.I0(n27907), .I1(t1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5733));   // verilog/neopixel.v(100[14:42])
    defparam i1_2_lut_adj_1792.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(t1[10]), .I1(n27910), .I2(t1[2]), .I3(n6_adj_5733), 
            .O(n27912));   // verilog/neopixel.v(100[14:42])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i22_4_lut (.I0(n60093), .I1(n61120), .I2(state[1]), .I3(start), 
            .O(n59349));
    defparam i22_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i51612_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i51612_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(t1[6]), .I1(t1[7]), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5732));   // verilog/neopixel.v(100[14:42])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i44909_2_lut (.I0(t1[1]), .I1(t1[3]), .I2(GND_net), .I3(GND_net), 
            .O(n64395));
    defparam i44909_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1793 (.I0(t1[2]), .I1(n27910), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5730));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1793.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n15), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n53_adj_5731));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i3_4_lut_adj_1794 (.I0(n27907), .I1(n32), .I2(t1[10]), .I3(t1[8]), 
            .O(n63023));
    defparam i3_4_lut_adj_1794.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut (.I0(state[1]), .I1(n63023), .I2(start), .I3(GND_net), 
            .O(n62573));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_1__I_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1800, ENCODER0_A_N_keep, 
            n1757, GND_net, n1759, n1761, n1763, n1765, n1767, 
            n1769, n1771, n1773, \encoder0_position[22] , \encoder0_position[21] , 
            \encoder0_position[20] , \encoder0_position[19] , \encoder0_position[18] , 
            \encoder0_position[17] , \encoder0_position[16] , \encoder0_position[15] , 
            \encoder0_position[14] , \encoder0_position[13] , \encoder0_position[12] , 
            \encoder0_position[11] , \encoder0_position[10] , \encoder0_position[9] , 
            \encoder0_position[8] , \encoder0_position[7] , \encoder0_position[6] , 
            \encoder0_position[5] , \encoder0_position[4] , \encoder0_position[3] , 
            \encoder0_position[2] , \encoder0_position[1] , \encoder0_position[0] , 
            VCC_net, \a_new[1] , \b_new[1] , n31820, n1755, n31819, 
            a_prev, n31817, b_prev, position_31__N_3836, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1800;
    input ENCODER0_A_N_keep;
    output n1757;
    input GND_net;
    output n1759;
    output n1761;
    output n1763;
    output n1765;
    output n1767;
    output n1769;
    output n1771;
    output n1773;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    output \a_new[1] ;
    output \b_new[1] ;
    input n31820;
    output n1755;
    input n31819;
    output a_prev;
    input n31817;
    output b_prev;
    output position_31__N_3836;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n53672, n53671, n53670, n53669, n53668, 
        n53667, n53666, n53665, n53664, n53663, n53662, n53661, 
        n53660, n53659, n53658, n53657, n53656, n53655, n53654, 
        n53653, n53652, n53651, n53650, n53649, n53648, n53647, 
        n53646, n53645, n53644, n53643, n53642;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1800), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1800), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1757), .I3(n53672), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1759), .I3(n53671), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n53671), .I0(direction_N_3840), 
            .I1(n1759), .CO(n53672));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1761), .I3(n53670), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n53670), .I0(direction_N_3840), 
            .I1(n1761), .CO(n53671));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1763), .I3(n53669), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n53669), .I0(direction_N_3840), 
            .I1(n1763), .CO(n53670));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1765), .I3(n53668), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n53668), .I0(direction_N_3840), 
            .I1(n1765), .CO(n53669));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1767), .I3(n53667), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n53667), .I0(direction_N_3840), 
            .I1(n1767), .CO(n53668));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1769), .I3(n53666), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n53666), .I0(direction_N_3840), 
            .I1(n1769), .CO(n53667));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1771), .I3(n53665), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n53665), .I0(direction_N_3840), 
            .I1(n1771), .CO(n53666));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1773), .I3(n53664), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n53664), .I0(direction_N_3840), 
            .I1(n1773), .CO(n53665));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n53663), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n53663), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n53664));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n53662), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n53662), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n53663));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n53661), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n53661), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n53662));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n53660), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n53660), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n53661));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n53659), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n53659), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n53660));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n53658), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n53658), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n53659));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n53657), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n53657), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n53658));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n53656), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n53656), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n53657));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n53655), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n53655), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n53656));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n53654), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n53654), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n53655));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n53653), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n53653), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n53654));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n53652), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n53652), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n53653));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n53651), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n53651), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n53652));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n53650), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n53650), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n53651));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n53649), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n53649), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n53650));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n53648), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n53648), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n53649));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n53647), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n53647), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n53648));
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n53646), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n53646), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n53647));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n53645), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_6 (.CI(n53645), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n53646));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n53644), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n53644), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n53645));
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n53643), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n53643), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n53644));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n53642), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n53642), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n53643));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n53642));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1800), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1800), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1755), .C(n1800), .D(n31820));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1800), .D(n31819));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1800), .D(n31817));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i0 (.Q(\encoder0_position[0] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(\encoder0_position[1] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(\encoder0_position[2] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(\encoder0_position[3] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(\encoder0_position[4] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(\encoder0_position[5] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(\encoder0_position[6] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(\encoder0_position[7] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(\encoder0_position[8] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(\encoder0_position[9] ), .C(n1800), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(\encoder0_position[10] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(\encoder0_position[11] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(\encoder0_position[12] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(\encoder0_position[13] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(\encoder0_position[14] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(\encoder0_position[15] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(\encoder0_position[16] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(\encoder0_position[17] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(\encoder0_position[18] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(\encoder0_position[19] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(\encoder0_position[20] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(\encoder0_position[21] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(\encoder0_position[22] ), .C(n1800), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(n1773), .C(n1800), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(n1771), .C(n1800), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(n1769), .C(n1800), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(n1767), .C(n1800), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(n1765), .C(n1800), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(n1763), .C(n1800), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(n1761), .C(n1800), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(n1759), .C(n1800), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i31 (.Q(n1757), .C(n1800), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (clk16MHz, GND_net, VCC_net, n30062, \current[15] , 
            n31866, \current[1] , n31865, \current[2] , n31864, \current[3] , 
            n31863, \current[4] , n31862, \current[5] , n31861, \current[6] , 
            n31860, \current[7] , n31859, \current[8] , n31858, \current[9] , 
            n31857, \current[10] , n31856, \current[11] , \data[15] , 
            \data[12] , CS_c, CS_CLK_c, n32677, n32676, n32675, 
            \data[11] , n32674, \data[10] , n32673, \data[9] , n32672, 
            \data[8] , n32671, \data[7] , n32670, \data[6] , n32669, 
            \data[5] , n32668, \data[4] , n32667, \data[3] , n32666, 
            \data[2] , n32665, \data[1] , n32299, \data[0] , n31699, 
            \current[0] , n27916, n27891, n11, n27938, n5, n5_adj_25, 
            n40832, n27925, n5_adj_26, state_7__N_4319) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    input GND_net;
    input VCC_net;
    output n30062;
    output \current[15] ;
    input n31866;
    output \current[1] ;
    input n31865;
    output \current[2] ;
    input n31864;
    output \current[3] ;
    input n31863;
    output \current[4] ;
    input n31862;
    output \current[5] ;
    input n31861;
    output \current[6] ;
    input n31860;
    output \current[7] ;
    input n31859;
    output \current[8] ;
    input n31858;
    output \current[9] ;
    input n31857;
    output \current[10] ;
    input n31856;
    output \current[11] ;
    output \data[15] ;
    output \data[12] ;
    output CS_c;
    output CS_CLK_c;
    input n32677;
    input n32676;
    input n32675;
    output \data[11] ;
    input n32674;
    output \data[10] ;
    input n32673;
    output \data[9] ;
    input n32672;
    output \data[8] ;
    input n32671;
    output \data[7] ;
    input n32670;
    output \data[6] ;
    input n32669;
    output \data[5] ;
    input n32668;
    output \data[4] ;
    input n32667;
    output \data[3] ;
    input n32666;
    output \data[2] ;
    input n32665;
    output \data[1] ;
    input n32299;
    output \data[0] ;
    input n31699;
    output \current[0] ;
    output n27916;
    output n27891;
    output n11;
    output n27938;
    output n5;
    output n5_adj_25;
    output n40832;
    output n27925;
    output n5_adj_26;
    output state_7__N_4319;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire clk_slow_N_4232;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n53634, n53633;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n53632, n53631, n53630, n53629, n53628, n53627, n53626, 
        n53625, n53624, n53623, n53622;
    wire [7:0]n37;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n53608, n53607, n53606, n53605, n67653, n53604, n2, n67659, 
        n53603, n67660, n53602, n67654;
    wire [13:0]n241;
    
    wire n30197, n31660, n24999, delay_counter_15__N_4314, clk_slow_N_4233;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n41177, n30129, n31165, clk_out, n9, n10548, n25003, 
        n31701, n25005, n25007, n15, n6, n6_adj_5728, n62544, 
        n8, n7;
    
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 counter_2050_2051_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n53634), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2050_2051_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n53633), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_3 (.CI(n53633), .I0(GND_net), .I1(counter[1]), 
            .CO(n53634));
    SB_LUT4 counter_2050_2051_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n53633));
    SB_LUT4 delay_counter_2048_2049_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n53632), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2048_2049_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n53631), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_12 (.CI(n53631), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n53632));
    SB_LUT4 delay_counter_2048_2049_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n53630), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_11 (.CI(n53630), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n53631));
    SB_LUT4 delay_counter_2048_2049_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n53629), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_10 (.CI(n53629), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n53630));
    SB_LUT4 delay_counter_2048_2049_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n53628), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_9 (.CI(n53628), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n53629));
    SB_LUT4 delay_counter_2048_2049_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n53627), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_8 (.CI(n53627), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n53628));
    SB_LUT4 delay_counter_2048_2049_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n53626), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_7 (.CI(n53626), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n53627));
    SB_LUT4 delay_counter_2048_2049_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n53625), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_6 (.CI(n53625), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n53626));
    SB_LUT4 delay_counter_2048_2049_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n53624), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_5 (.CI(n53624), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n53625));
    SB_LUT4 delay_counter_2048_2049_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n53623), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_4 (.CI(n53623), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n53624));
    SB_LUT4 delay_counter_2048_2049_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n53622), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_3 (.CI(n53622), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n53623));
    SB_LUT4 delay_counter_2048_2049_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n53622));
    SB_LUT4 bit_counter_2044_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n53608), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2044_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n53607), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_8 (.CI(n53607), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n53608));
    SB_LUT4 bit_counter_2044_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n53606), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_7 (.CI(n53606), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n53607));
    SB_LUT4 bit_counter_2044_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n53605), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_6 (.CI(n53605), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n53606));
    SB_LUT4 bit_counter_2044_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n53604), .O(n67653)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_5 (.CI(n53604), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n53605));
    SB_LUT4 bit_counter_2044_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n53603), .O(n67659)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_4 (.CI(n53603), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n53604));
    SB_LUT4 bit_counter_2044_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n53602), .O(n67660)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_3 (.CI(n53602), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n53603));
    SB_LUT4 bit_counter_2044_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n67654)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n53602));
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n30062), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_2044__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n30197), 
            .D(n37[7]), .R(n31660));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n30197), 
            .D(n37[6]), .R(n31660));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n30197), 
            .D(n37[5]), .R(n31660));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n30197), 
            .D(n37[4]), .R(n31660));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n31866));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n31865));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n31864));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n31863));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n31862));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n31861));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n31860));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n31859));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n31858));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n31857));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n31856));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n30197), 
            .D(n24999));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i51468_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n30062));
    defparam i51468_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2243_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2243_1_lut.LUT_INIT = 16'h5555;
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n30129), .D(n41177), 
            .S(n31165));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2521_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2521_1_lut.LUT_INIT = 16'h5555;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n32677));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n32676));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n32675));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n32674));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n32673));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n32672));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n32671));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n32670));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n32669));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n32668));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n32667));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n32666));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n32665));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n32299));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n30129), .D(n10548), 
            .R(n31165));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n30197), 
            .D(n25003));   // verilog/tli4970.v(55[24:39])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n31701));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n31699));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n30197), 
            .D(n25005));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n30197), 
            .D(n25007));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i2179_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2179_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7072_3_lut (.I0(state[0]), .I1(n67653), .I2(state[1]), .I3(GND_net), 
            .O(n25007));   // verilog/tli4970.v(55[24:39])
    defparam i7072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7070_3_lut (.I0(state[0]), .I1(n67659), .I2(state[1]), .I3(GND_net), 
            .O(n25005));   // verilog/tli4970.v(55[24:39])
    defparam i7070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7068_3_lut (.I0(state[0]), .I1(n67660), .I2(state[1]), .I3(GND_net), 
            .O(n25003));   // verilog/tli4970.v(55[24:39])
    defparam i7068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2153_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n10548));
    defparam mux_2153_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13469_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31660));   // verilog/tli4970.v(55[24:39])
    defparam i13469_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(bit_counter[3]), 
            .I3(bit_counter[2]), .O(n27916));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1777 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n27891));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1777.LUT_INIT = 16'hffbf;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1778 (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n27938));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1778.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_25));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n30129));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i12974_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n31165));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12974_2_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 i22740_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n40832));
    defparam i22740_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n27925));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_330_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_26));   // verilog/tli4970.v(54[9:26])
    defparam equal_330_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51503_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n41177));
    defparam i51503_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1779 (.I0(delay_counter[2]), .I1(delay_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5728));
    defparam i1_2_lut_adj_1779.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1780 (.I0(delay_counter[3]), .I1(delay_counter[1]), 
            .I2(delay_counter[0]), .I3(n6_adj_5728), .O(n62544));
    defparam i4_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n62544), .I1(delay_counter[10]), .I2(delay_counter[6]), 
            .I3(delay_counter[5]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i1_2_lut_adj_1781 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(delay_counter[9]), .I1(n7), .I2(delay_counter[8]), 
            .I3(n8), .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7065_3_lut (.I0(state[0]), .I1(n67654), .I2(state[1]), .I3(GND_net), 
            .O(n24999));   // verilog/tli4970.v(55[24:39])
    defparam i7065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12084_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n30197));
    defparam i12084_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13510_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n31701));
    defparam i13510_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i51681_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9));
    defparam i51681_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1800, ENCODER1_A_N_keep, 
            \a_new[1] , encoder1_position, GND_net, \b_new[1] , b_prev, 
            VCC_net, n31821, a_prev, position_31__N_3836, n31707, 
            n31706, n1805, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1800;
    input ENCODER1_A_N_keep;
    output \a_new[1] ;
    output [31:0]encoder1_position;
    input GND_net;
    output \b_new[1] ;
    output b_prev;
    input VCC_net;
    input n31821;
    output a_prev;
    output position_31__N_3836;
    input n31707;
    input n31706;
    output n1805;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n53570, n53569, n53568, n53567, n53566, 
        n53565, n53564, n53563, n53562, n53561, n53560, n53559, 
        n53558, n53557, n53556, n53555, n53554, n53553, n53552, 
        n53551, n53550, n53549, n53548, n53547, n53546, n53545, 
        n53544, n53543, n53542, n53541, n53540;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1800), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1800), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1800), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2041_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[31]), .I3(n53570), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2041_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[30]), .I3(n53569), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_32 (.CI(n53569), .I0(direction_N_3840), 
            .I1(encoder1_position[30]), .CO(n53570));
    SB_LUT4 position_2041_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[29]), .I3(n53568), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_31 (.CI(n53568), .I0(direction_N_3840), 
            .I1(encoder1_position[29]), .CO(n53569));
    SB_LUT4 position_2041_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[28]), .I3(n53567), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_30 (.CI(n53567), .I0(direction_N_3840), 
            .I1(encoder1_position[28]), .CO(n53568));
    SB_LUT4 position_2041_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[27]), .I3(n53566), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_29 (.CI(n53566), .I0(direction_N_3840), 
            .I1(encoder1_position[27]), .CO(n53567));
    SB_LUT4 position_2041_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[26]), .I3(n53565), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_28 (.CI(n53565), .I0(direction_N_3840), 
            .I1(encoder1_position[26]), .CO(n53566));
    SB_LUT4 position_2041_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[25]), .I3(n53564), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_27 (.CI(n53564), .I0(direction_N_3840), 
            .I1(encoder1_position[25]), .CO(n53565));
    SB_LUT4 position_2041_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[24]), .I3(n53563), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_26 (.CI(n53563), .I0(direction_N_3840), 
            .I1(encoder1_position[24]), .CO(n53564));
    SB_LUT4 position_2041_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[23]), .I3(n53562), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1800), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_CARRY position_2041_add_4_25 (.CI(n53562), .I0(direction_N_3840), 
            .I1(encoder1_position[23]), .CO(n53563));
    SB_LUT4 position_2041_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[22]), .I3(n53561), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_24 (.CI(n53561), .I0(direction_N_3840), 
            .I1(encoder1_position[22]), .CO(n53562));
    SB_LUT4 position_2041_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[21]), .I3(n53560), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_23 (.CI(n53560), .I0(direction_N_3840), 
            .I1(encoder1_position[21]), .CO(n53561));
    SB_LUT4 position_2041_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[20]), .I3(n53559), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_22 (.CI(n53559), .I0(direction_N_3840), 
            .I1(encoder1_position[20]), .CO(n53560));
    SB_LUT4 position_2041_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[19]), .I3(n53558), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_21 (.CI(n53558), .I0(direction_N_3840), 
            .I1(encoder1_position[19]), .CO(n53559));
    SB_LUT4 position_2041_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[18]), .I3(n53557), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_20 (.CI(n53557), .I0(direction_N_3840), 
            .I1(encoder1_position[18]), .CO(n53558));
    SB_LUT4 position_2041_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[17]), .I3(n53556), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_19 (.CI(n53556), .I0(direction_N_3840), 
            .I1(encoder1_position[17]), .CO(n53557));
    SB_LUT4 position_2041_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[16]), .I3(n53555), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_18 (.CI(n53555), .I0(direction_N_3840), 
            .I1(encoder1_position[16]), .CO(n53556));
    SB_LUT4 position_2041_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[15]), .I3(n53554), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_17 (.CI(n53554), .I0(direction_N_3840), 
            .I1(encoder1_position[15]), .CO(n53555));
    SB_LUT4 position_2041_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[14]), .I3(n53553), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_16 (.CI(n53553), .I0(direction_N_3840), 
            .I1(encoder1_position[14]), .CO(n53554));
    SB_LUT4 position_2041_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[13]), .I3(n53552), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_15 (.CI(n53552), .I0(direction_N_3840), 
            .I1(encoder1_position[13]), .CO(n53553));
    SB_LUT4 position_2041_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[12]), .I3(n53551), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY position_2041_add_4_14 (.CI(n53551), .I0(direction_N_3840), 
            .I1(encoder1_position[12]), .CO(n53552));
    SB_LUT4 position_2041_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[11]), .I3(n53550), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_13 (.CI(n53550), .I0(direction_N_3840), 
            .I1(encoder1_position[11]), .CO(n53551));
    SB_LUT4 position_2041_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[10]), .I3(n53549), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_12 (.CI(n53549), .I0(direction_N_3840), 
            .I1(encoder1_position[10]), .CO(n53550));
    SB_LUT4 position_2041_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[9]), .I3(n53548), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_11 (.CI(n53548), .I0(direction_N_3840), 
            .I1(encoder1_position[9]), .CO(n53549));
    SB_LUT4 position_2041_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[8]), .I3(n53547), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_10 (.CI(n53547), .I0(direction_N_3840), 
            .I1(encoder1_position[8]), .CO(n53548));
    SB_LUT4 position_2041_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[7]), .I3(n53546), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_9 (.CI(n53546), .I0(direction_N_3840), 
            .I1(encoder1_position[7]), .CO(n53547));
    SB_LUT4 position_2041_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[6]), .I3(n53545), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_8 (.CI(n53545), .I0(direction_N_3840), 
            .I1(encoder1_position[6]), .CO(n53546));
    SB_LUT4 position_2041_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[5]), .I3(n53544), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_7 (.CI(n53544), .I0(direction_N_3840), 
            .I1(encoder1_position[5]), .CO(n53545));
    SB_LUT4 position_2041_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[4]), .I3(n53543), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_6 (.CI(n53543), .I0(direction_N_3840), 
            .I1(encoder1_position[4]), .CO(n53544));
    SB_LUT4 position_2041_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[3]), .I3(n53542), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_5 (.CI(n53542), .I0(direction_N_3840), 
            .I1(encoder1_position[3]), .CO(n53543));
    SB_LUT4 position_2041_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[2]), .I3(n53541), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_4 (.CI(n53541), .I0(direction_N_3840), 
            .I1(encoder1_position[2]), .CO(n53542));
    SB_LUT4 position_2041_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[1]), .I3(n53540), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_3 (.CI(n53540), .I0(direction_N_3840), 
            .I1(encoder1_position[1]), .CO(n53541));
    SB_LUT4 position_2041_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n53540));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1800), .D(n31821));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i0 (.Q(encoder1_position[0]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1800), .D(n31707));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1805), .C(n1800), .D(n31706));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i1 (.Q(encoder1_position[1]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i2 (.Q(encoder1_position[2]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i3 (.Q(encoder1_position[3]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i4 (.Q(encoder1_position[4]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i5 (.Q(encoder1_position[5]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i6 (.Q(encoder1_position[6]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i7 (.Q(encoder1_position[7]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i8 (.Q(encoder1_position[8]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i9 (.Q(encoder1_position[9]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i10 (.Q(encoder1_position[10]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i11 (.Q(encoder1_position[11]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i12 (.Q(encoder1_position[12]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i13 (.Q(encoder1_position[13]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i14 (.Q(encoder1_position[14]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i15 (.Q(encoder1_position[15]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i16 (.Q(encoder1_position[16]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i17 (.Q(encoder1_position[17]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i18 (.Q(encoder1_position[18]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i19 (.Q(encoder1_position[19]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i20 (.Q(encoder1_position[20]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i21 (.Q(encoder1_position[21]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i22 (.Q(encoder1_position[22]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i23 (.Q(encoder1_position[23]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i24 (.Q(encoder1_position[24]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i25 (.Q(encoder1_position[25]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i26 (.Q(encoder1_position[26]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i27 (.Q(encoder1_position[27]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i28 (.Q(encoder1_position[28]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i29 (.Q(encoder1_position[29]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i30 (.Q(encoder1_position[30]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i31 (.Q(encoder1_position[31]), .C(n1800), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (reset, rx_data, \data_in_frame[6] , n2887, \data_out_frame[18] , 
            clk16MHz, n59931, n59925, n59095, VCC_net, \data_in_frame[16] , 
            n59924, n32202, n59923, n59922, n59921, n59933, n59920, 
            \data_out_frame[19] , n59919, n59918, n59917, n59916, 
            \data_in_frame[4] , n59915, n59914, n59913, n59912, \data_out_frame[20] , 
            n59911, \data_out_frame[0][2] , n59934, n32199, \data_out_frame[0][3] , 
            n60050, n59473, \data_out_frame[0][4] , n60049, \data_out_frame[1][0] , 
            n60048, \data_out_frame[1][1] , n60047, n59910, \data_out_frame[1][3] , 
            n60046, \data_out_frame[1][5] , n59932, \data_out_frame[6] , 
            \data_out_frame[7] , byte_transmit_counter, GND_net, \data_out_frame[4] , 
            \data_out_frame[5] , \data_out_frame[1][6] , n60045, n59909, 
            n59908, n59907, n59906, n59905, n59904, \data_out_frame[21] , 
            n59903, n59902, n59901, n59900, n59899, n31492, n59898, 
            \data_out_frame[1][7] , n60044, n31490, \data_out_frame[22] , 
            n59897, n59896, \data_out_frame[3][1] , n60043, \data_out_frame[13] , 
            n67793, \data_out_frame[3][3] , n60042, \data_in_frame[2] , 
            deadband, \data_in_frame[13] , IntegralLimit, \data_in_frame[3] , 
            \Kp[0] , \data_in_frame[5] , \Ki[0] , \data_in_frame[10] , 
            PWMLimit, \data_out_frame[3][4] , n60041, \data_out_frame[3][6] , 
            n60040, \data_out_frame[3][7] , n60039, n60038, n60037, 
            n59936, n60036, n60035, n60034, n32171, \data_in_frame[14] , 
            n60033, n32168, n60032, n32165, n60031, n59895, n59894, 
            n59893, n31484, n59892, n59891, \data_out_frame[23] , 
            n59890, n59889, n32162, n60030, n31793, n60029, n32158, 
            n59888, n59887, n59886, n60028, n59885, n31475, n31474, 
            \data_out_frame[24] , n59884, n59883, n31471, n31470, 
            n32155, n59882, n59881, n31467, n59880, \data_out_frame[25] , 
            n59879, n59878, n60027, n59873, \data_in_frame[9] , \data_out_frame[9] , 
            n59877, \data_out_frame[10] , \data_out_frame[11] , n31461, 
            n60134, n32152, n31460, \data_out_frame[14] , \data_out_frame[15] , 
            \data_out_frame[12] , n59876, n59875, \FRAME_MATCHER.state[3] , 
            n60514, \data_out_frame[26] , n60082, \data_out_frame[16] , 
            \data_out_frame[17] , n32149, n60026, LED_c, n60081, \Ki[15] , 
            \FRAME_MATCHER.i_31__N_2513 , n35072, n31455, \Ki[14] , 
            \Ki[13] , setpoint, \Ki[12] , n32146, n60080, n60076, 
            \Ki[11] , n60077, \Ki[10] , n31451, \Ki[9] , n64802, 
            \Ki[8] , \Ki[7] , n60075, n60025, \data_out_frame[27] , 
            n60072, \Ki[6] , n60073, \FRAME_MATCHER.i_31__N_2509 , \encoder0_position_scaled[21] , 
            n31447, n32143, n60078, n60079, n32140, \Ki[5] , \Ki[4] , 
            \Ki[3] , \Ki[2] , n60071, n55748, \Ki[1] , \Kp[15] , 
            n60024, n55746, \encoder0_position_scaled[20] , \Kp[14] , 
            n31443, n60074, n60414, n55760, n60523, \Kp[13] , \encoder0_position_scaled[19] , 
            \Kp[12] , \Kp[11] , n55781, n32137, \Kp[10] , n32134, 
            n60150, n31796, n60023, n32130, n32127, n32124, n55267, 
            n55737, \Kp[9] , n60022, \Kp[8] , n60021, \Kp[7] , \Kp[6] , 
            n71628, \data_out_frame[8][2] , \FRAME_MATCHER.i[2] , \FRAME_MATCHER.i[1] , 
            \data_in_frame[3][5] , \Kp[5] , \data_in_frame[21][7] , \data_in_frame[17] , 
            \data_in_frame[20] , \data_in_frame[18] , \data_in_frame[21][1] , 
            \data_in_frame[21][2] , \data_in_frame[21][4] , \data_in_frame[21][0] , 
            \data_in_frame[18][7] , \Kp[4] , \FRAME_MATCHER.i[0] , \data_in_frame[21][3] , 
            n31802, \data_in_frame[3][3] , \Kp[3] , \Kp[2] , \Kp[1] , 
            n60020, \data_in_frame[18][1] , \data_in_frame[18][3] , n60019, 
            n32068, n32065, n32062, n60018, n71574, control_mode, 
            n62692, n30673, n32059, n32056, n32053, n32050, n32047, 
            n32044, n32041, n32038, n31806, \control_mode[6] , \control_mode[7] , 
            n31811, n31853, n31916, n31919, n31922, n31925, n32018, 
            n32015, n60609, n32012, n32009, n32005, n60017, \data_in_frame[6][6] , 
            \data_in_frame[17][6] , \data_in_frame[18][0] , DE_c, n60016, 
            n60015, n60014, n60013, n60012, n60011, n60010, n60009, 
            n60008, \data_out_frame[8][1] , n60007, n60006, \data_out_frame[8][3] , 
            n60005, \data_out_frame[8][4] , n60004, \data_out_frame[8][5] , 
            n60003, \data_out_frame[8][6] , n60002, \data_out_frame[8][7] , 
            n60001, n60000, n59999, n59998, n59997, n59996, n59995, 
            n59994, n59993, n59992, n59991, n59990, n59989, n59988, 
            n59987, n59986, n59985, n59984, n59983, n59982, n59981, 
            n59980, n59979, n59978, n59977, n59976, n59975, n59974, 
            n59973, n59972, n60051, n59971, n59970, n59935, n59969, 
            n59968, n59967, n59966, n59965, n59964, n59963, n59962, 
            n59961, n59960, n59959, n59958, n59957, n59956, n59955, 
            n59954, n59953, n59952, n59951, n59950, n59949, n59948, 
            n59947, n59946, n59874, n59945, n59944, n59943, n59942, 
            n59941, n59940, n31818, \FRAME_MATCHER.rx_data_ready_prev , 
            n59939, n59938, n59937, n59930, displacement, n59929, 
            \data_in_frame[1] , n59928, \data_in_frame[22] , \data_in_frame[22][3] , 
            \data_in_frame[22][7] , Kp_23__N_715, n60538, Kp_23__N_869, 
            n3489, n59927, \encoder0_position_scaled[18] , \encoder0_position_scaled[17] , 
            n59203, n39602, n61124, n76, n59201, n59197, n59193, 
            n59189, n59315, n32704, n59313, n59185, n59181, n59177, 
            n32290, n32300, \data_in_frame[18][5] , n59173, n32306, 
            n32632, n32363, n59263, n59265, n59255, n59309, \data_in_frame[21][5] , 
            n32387, n32390, n32393, n32396, n32403, \data_in_frame[22][5] , 
            n32406, n32409, n31736, n31739, n31742, n32489, neopxl_color, 
            n32488, n32487, n32484, n32483, n32482, n32481, n32480, 
            n32479, n32478, n32477, n32475, n32474, n32472, n32471, 
            n32470, n32469, n32468, n32467, \control_mode[1] , n31745, 
            n32462, n32461, n32460, n32459, n32458, current_limit, 
            n32457, n37917, n32455, n30619, n59926, n32454, n32452, 
            n32451, n32450, n32449, n32448, n32447, n32446, n32445, 
            n32444, n31748, n31751, n31754, n31757, n67702, n59777, 
            n31766, n31772, n31695, \control_mode[0] , n31693, n31784, 
            n31787, \encoder0_position_scaled[16] , ID, n55567, \encoder0_position_scaled[22] , 
            n71580, n55802, n30671, n25151, pwm_setpoint, n25082, 
            n8, rx_data_ready, n65, n30627, n59773, n67698, n89, 
            n30669, tx_active, control_update, n30039, n30709, n30708, 
            n15, n30702, n15_adj_6, n15_adj_7, \current[15] , n7, 
            n64811, n64809, n30700, n59779, n28460, encoder1_position_scaled, 
            n41236, \encoder0_position_scaled[7] , \encoder0_position_scaled[6] , 
            \encoder0_position_scaled[5] , \encoder0_position_scaled[4] , 
            \encoder0_position_scaled[3] , \encoder0_position_scaled[2] , 
            \encoder0_position_scaled[1] , n6, \encoder0_position_scaled[15] , 
            \encoder0_position_scaled[14] , n8_adj_8, n30621, \encoder0_position_scaled[13] , 
            \encoder0_position_scaled[12] , \encoder0_position_scaled[11] , 
            \encoder0_position_scaled[10] , \encoder0_position_scaled[9] , 
            \encoder0_position_scaled[8] , \encoder0_position_scaled[23] , 
            n39603, \current[7] , \current[6] , \current[5] , n30623, 
            \current[4] , \current[3] , \current[2] , n59772, n30323, 
            \current[1] , n30278, n64817, n64815, \current[0] , \current[11] , 
            \current[10] , \current[9] , \current[8] , n64584, n64585, 
            n64582, n64581, n1, tx_o, \tx_data[0] , r_SM_Main, \r_Bit_Index[0] , 
            n59789, n63279, n27, \r_SM_Main_2__N_3536[1] , r_Clock_Count, 
            n32272, n71737, n30087, n31705, n5233, \o_Rx_DV_N_3488[12] , 
            \o_Rx_DV_N_3488[24] , n29, n23, n61776, n6_adj_9, n60925, 
            n63255, tx_enable, baudrate, n27889, r_SM_Main_adj_23, 
            r_Rx_Data, RX_N_2, r_Clock_Count_adj_24, \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \r_Bit_Index[0]_adj_21 , n59798, n63269, 
            \r_SM_Main_2__N_3446[1] , \o_Rx_DV_N_3488[0] , n5230, n32278, 
            n55993, n30084, n32606, n32605, n32604, n32603, n32600, 
            n32599, n32598, n32286, n60086, n4, n6_adj_22, n30080, 
            n60927, n63257, n63621, n63605, n63549, n63515, n63551, 
            n63641, n63587, n63623) /* synthesis syn_module_defined=1 */ ;
    input reset;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[6] ;
    input n2887;
    output [7:0]\data_out_frame[18] ;
    input clk16MHz;
    input n59931;
    input n59925;
    input n59095;
    input VCC_net;
    output [7:0]\data_in_frame[16] ;
    input n59924;
    input n32202;
    input n59923;
    input n59922;
    input n59921;
    input n59933;
    input n59920;
    output [7:0]\data_out_frame[19] ;
    input n59919;
    input n59918;
    input n59917;
    input n59916;
    output [7:0]\data_in_frame[4] ;
    input n59915;
    input n59914;
    input n59913;
    input n59912;
    output [7:0]\data_out_frame[20] ;
    input n59911;
    output \data_out_frame[0][2] ;
    input n59934;
    input n32199;
    output \data_out_frame[0][3] ;
    input n60050;
    input n59473;
    output \data_out_frame[0][4] ;
    input n60049;
    output \data_out_frame[1][0] ;
    input n60048;
    output \data_out_frame[1][1] ;
    input n60047;
    input n59910;
    output \data_out_frame[1][3] ;
    input n60046;
    output \data_out_frame[1][5] ;
    input n59932;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]byte_transmit_counter;
    input GND_net;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output \data_out_frame[1][6] ;
    input n60045;
    input n59909;
    input n59908;
    input n59907;
    input n59906;
    input n59905;
    input n59904;
    output [7:0]\data_out_frame[21] ;
    input n59903;
    input n59902;
    input n59901;
    input n59900;
    input n59899;
    input n31492;
    input n59898;
    output \data_out_frame[1][7] ;
    input n60044;
    input n31490;
    output [7:0]\data_out_frame[22] ;
    input n59897;
    input n59896;
    output \data_out_frame[3][1] ;
    input n60043;
    output [7:0]\data_out_frame[13] ;
    input n67793;
    output \data_out_frame[3][3] ;
    input n60042;
    output [7:0]\data_in_frame[2] ;
    output [23:0]deadband;
    output [7:0]\data_in_frame[13] ;
    output [23:0]IntegralLimit;
    output [7:0]\data_in_frame[3] ;
    output \Kp[0] ;
    output [7:0]\data_in_frame[5] ;
    output \Ki[0] ;
    output [7:0]\data_in_frame[10] ;
    output [23:0]PWMLimit;
    output \data_out_frame[3][4] ;
    input n60041;
    output \data_out_frame[3][6] ;
    input n60040;
    output \data_out_frame[3][7] ;
    input n60039;
    input n60038;
    input n60037;
    input n59936;
    input n60036;
    input n60035;
    input n60034;
    input n32171;
    output [7:0]\data_in_frame[14] ;
    input n60033;
    input n32168;
    input n60032;
    input n32165;
    input n60031;
    input n59895;
    input n59894;
    input n59893;
    input n31484;
    input n59892;
    input n59891;
    output [7:0]\data_out_frame[23] ;
    input n59890;
    input n59889;
    input n32162;
    input n60030;
    input n31793;
    input n60029;
    input n32158;
    input n59888;
    input n59887;
    input n59886;
    input n60028;
    input n59885;
    input n31475;
    input n31474;
    output [7:0]\data_out_frame[24] ;
    input n59884;
    input n59883;
    input n31471;
    input n31470;
    input n32155;
    input n59882;
    input n59881;
    input n31467;
    input n59880;
    output [7:0]\data_out_frame[25] ;
    input n59879;
    input n59878;
    input n60027;
    input n59873;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_out_frame[9] ;
    input n59877;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    input n31461;
    output n60134;
    input n32152;
    input n31460;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    input n59876;
    input n59875;
    output \FRAME_MATCHER.state[3] ;
    input n60514;
    output [7:0]\data_out_frame[26] ;
    input n60082;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    input n32149;
    input n60026;
    output LED_c;
    input n60081;
    output \Ki[15] ;
    output \FRAME_MATCHER.i_31__N_2513 ;
    output n35072;
    input n31455;
    output \Ki[14] ;
    output \Ki[13] ;
    output [23:0]setpoint;
    output \Ki[12] ;
    input n32146;
    input n60080;
    input n60076;
    output \Ki[11] ;
    input n60077;
    output \Ki[10] ;
    input n31451;
    output \Ki[9] ;
    output n64802;
    output \Ki[8] ;
    output \Ki[7] ;
    input n60075;
    input n60025;
    output [7:0]\data_out_frame[27] ;
    input n60072;
    output \Ki[6] ;
    input n60073;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input \encoder0_position_scaled[21] ;
    input n31447;
    input n32143;
    input n60078;
    input n60079;
    input n32140;
    output \Ki[5] ;
    output \Ki[4] ;
    output \Ki[3] ;
    output \Ki[2] ;
    input n60071;
    output n55748;
    output \Ki[1] ;
    output \Kp[15] ;
    input n60024;
    input n55746;
    input \encoder0_position_scaled[20] ;
    output \Kp[14] ;
    input n31443;
    input n60074;
    output n60414;
    output n55760;
    output n60523;
    output \Kp[13] ;
    input \encoder0_position_scaled[19] ;
    output \Kp[12] ;
    output \Kp[11] ;
    input n55781;
    input n32137;
    output \Kp[10] ;
    input n32134;
    output n60150;
    input n31796;
    input n60023;
    input n32130;
    input n32127;
    input n32124;
    output n55267;
    input n55737;
    output \Kp[9] ;
    input n60022;
    output \Kp[8] ;
    input n60021;
    output \Kp[7] ;
    output \Kp[6] ;
    output n71628;
    output \data_out_frame[8][2] ;
    output \FRAME_MATCHER.i[2] ;
    output \FRAME_MATCHER.i[1] ;
    output \data_in_frame[3][5] ;
    output \Kp[5] ;
    output \data_in_frame[21][7] ;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[20] ;
    output [7:0]\data_in_frame[18] ;
    output \data_in_frame[21][1] ;
    output \data_in_frame[21][2] ;
    output \data_in_frame[21][4] ;
    output \data_in_frame[21][0] ;
    output \data_in_frame[18][7] ;
    output \Kp[4] ;
    output \FRAME_MATCHER.i[0] ;
    output \data_in_frame[21][3] ;
    input n31802;
    output \data_in_frame[3][3] ;
    output \Kp[3] ;
    output \Kp[2] ;
    output \Kp[1] ;
    input n60020;
    output \data_in_frame[18][1] ;
    output \data_in_frame[18][3] ;
    input n60019;
    input n32068;
    input n32065;
    input n32062;
    input n60018;
    output n71574;
    output [7:0]control_mode;
    output n62692;
    output n30673;
    input n32059;
    input n32056;
    input n32053;
    input n32050;
    input n32047;
    input n32044;
    input n32041;
    input n32038;
    input n31806;
    output \control_mode[6] ;
    output \control_mode[7] ;
    input n31811;
    input n31853;
    input n31916;
    input n31919;
    input n31922;
    input n31925;
    input n32018;
    input n32015;
    input n60609;
    input n32012;
    input n32009;
    input n32005;
    input n60017;
    output \data_in_frame[6][6] ;
    output \data_in_frame[17][6] ;
    output \data_in_frame[18][0] ;
    output DE_c;
    input n60016;
    input n60015;
    input n60014;
    input n60013;
    input n60012;
    input n60011;
    input n60010;
    input n60009;
    input n60008;
    output \data_out_frame[8][1] ;
    input n60007;
    input n60006;
    output \data_out_frame[8][3] ;
    input n60005;
    output \data_out_frame[8][4] ;
    input n60004;
    output \data_out_frame[8][5] ;
    input n60003;
    output \data_out_frame[8][6] ;
    input n60002;
    output \data_out_frame[8][7] ;
    input n60001;
    input n60000;
    input n59999;
    input n59998;
    input n59997;
    input n59996;
    input n59995;
    input n59994;
    input n59993;
    input n59992;
    input n59991;
    input n59990;
    input n59989;
    input n59988;
    input n59987;
    input n59986;
    input n59985;
    input n59984;
    input n59983;
    input n59982;
    input n59981;
    input n59980;
    input n59979;
    input n59978;
    input n59977;
    input n59976;
    input n59975;
    input n59974;
    input n59973;
    input n59972;
    input n60051;
    input n59971;
    input n59970;
    input n59935;
    input n59969;
    input n59968;
    input n59967;
    input n59966;
    input n59965;
    input n59964;
    input n59963;
    input n59962;
    input n59961;
    input n59960;
    input n59959;
    input n59958;
    input n59957;
    input n59956;
    input n59955;
    input n59954;
    input n59953;
    input n59952;
    input n59951;
    input n59950;
    input n59949;
    input n59948;
    input n59947;
    input n59946;
    input n59874;
    input n59945;
    input n59944;
    input n59943;
    input n59942;
    input n59941;
    input n59940;
    input n31818;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n59939;
    input n59938;
    input n59937;
    input n59930;
    input [23:0]displacement;
    input n59929;
    output [7:0]\data_in_frame[1] ;
    input n59928;
    output [7:0]\data_in_frame[22] ;
    output \data_in_frame[22][3] ;
    output \data_in_frame[22][7] ;
    output Kp_23__N_715;
    input n60538;
    output Kp_23__N_869;
    output n3489;
    input n59927;
    input \encoder0_position_scaled[18] ;
    input \encoder0_position_scaled[17] ;
    input n59203;
    output n39602;
    output n61124;
    output n76;
    input n59201;
    input n59197;
    input n59193;
    input n59189;
    input n59315;
    input n32704;
    input n59313;
    input n59185;
    input n59181;
    input n59177;
    input n32290;
    input n32300;
    output \data_in_frame[18][5] ;
    input n59173;
    input n32306;
    input n32632;
    input n32363;
    input n59263;
    input n59265;
    input n59255;
    input n59309;
    output \data_in_frame[21][5] ;
    input n32387;
    input n32390;
    input n32393;
    input n32396;
    input n32403;
    output \data_in_frame[22][5] ;
    input n32406;
    input n32409;
    input n31736;
    input n31739;
    input n31742;
    input n32489;
    output [23:0]neopxl_color;
    input n32488;
    input n32487;
    input n32484;
    input n32483;
    input n32482;
    input n32481;
    input n32480;
    input n32479;
    input n32478;
    input n32477;
    input n32475;
    input n32474;
    input n32472;
    input n32471;
    input n32470;
    input n32469;
    input n32468;
    input n32467;
    output \control_mode[1] ;
    input n31745;
    input n32462;
    input n32461;
    input n32460;
    input n32459;
    input n32458;
    output [15:0]current_limit;
    input n32457;
    input n37917;
    input n32455;
    output n30619;
    input n59926;
    input n32454;
    input n32452;
    input n32451;
    input n32450;
    input n32449;
    input n32448;
    input n32447;
    input n32446;
    input n32445;
    input n32444;
    input n31748;
    input n31751;
    input n31754;
    input n31757;
    output n67702;
    output n59777;
    input n31766;
    input n31772;
    input n31695;
    output \control_mode[0] ;
    input n31693;
    input n31784;
    input n31787;
    input \encoder0_position_scaled[16] ;
    input [7:0]ID;
    output n55567;
    input \encoder0_position_scaled[22] ;
    input n71580;
    output n55802;
    output n30671;
    output n25151;
    input [23:0]pwm_setpoint;
    input n25082;
    output n8;
    output rx_data_ready;
    output n65;
    output n30627;
    output n59773;
    output n67698;
    output n89;
    output n30669;
    output tx_active;
    input control_update;
    output n30039;
    output n30709;
    input n30708;
    output n15;
    output n30702;
    output n15_adj_6;
    output n15_adj_7;
    input \current[15] ;
    output n7;
    input n64811;
    input n64809;
    input n30700;
    output n59779;
    output n28460;
    input [23:0]encoder1_position_scaled;
    input n41236;
    input \encoder0_position_scaled[7] ;
    input \encoder0_position_scaled[6] ;
    input \encoder0_position_scaled[5] ;
    input \encoder0_position_scaled[4] ;
    input \encoder0_position_scaled[3] ;
    input \encoder0_position_scaled[2] ;
    input \encoder0_position_scaled[1] ;
    output n6;
    input \encoder0_position_scaled[15] ;
    input \encoder0_position_scaled[14] ;
    output n8_adj_8;
    input n30621;
    input \encoder0_position_scaled[13] ;
    input \encoder0_position_scaled[12] ;
    input \encoder0_position_scaled[11] ;
    input \encoder0_position_scaled[10] ;
    input \encoder0_position_scaled[9] ;
    input \encoder0_position_scaled[8] ;
    input \encoder0_position_scaled[23] ;
    input n39603;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    output n30623;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    output n59772;
    output n30323;
    input \current[1] ;
    output n30278;
    input n64817;
    input n64815;
    input \current[0] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input n64584;
    input n64585;
    input n64582;
    input n64581;
    output n1;
    output tx_o;
    input \tx_data[0] ;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output n59789;
    input n63279;
    output n27;
    input \r_SM_Main_2__N_3536[1] ;
    output [8:0]r_Clock_Count;
    input n32272;
    input n71737;
    output n30087;
    input n31705;
    input n5233;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    input n61776;
    output n6_adj_9;
    output n60925;
    output n63255;
    output tx_enable;
    input [31:0]baudrate;
    output n27889;
    output [2:0]r_SM_Main_adj_23;
    output r_Rx_Data;
    input RX_N_2;
    output [7:0]r_Clock_Count_adj_24;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0]_adj_21 ;
    output n59798;
    input n63269;
    input \r_SM_Main_2__N_3446[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n5230;
    input n32278;
    input n55993;
    output n30084;
    input n32606;
    input n32605;
    input n32604;
    input n32603;
    input n32600;
    input n32599;
    input n32598;
    input n32286;
    input n60086;
    output n4;
    output n6_adj_22;
    output n30080;
    output n60927;
    output n63257;
    input n63621;
    output n63605;
    input n63549;
    output n63515;
    output n63551;
    output n63641;
    output n63587;
    output n63623;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n30637, n31949, n2, n2_adj_5316, n2_adj_5317, n2_adj_5318, 
        n2_adj_5319, n2_adj_5320, n2_adj_5321, n8_c, n59771;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    
    wire n32121, n2_adj_5322, n2_adj_5323, n2_adj_5324, n2_adj_5325, 
        n2_adj_5326, n54798, Kp_23__N_878, n60217, Kp_23__N_993, n2_adj_5327, 
        n2_adj_5328, n2_adj_5329, n2_adj_5330, n2_adj_5331, n2_adj_5332, 
        n2_adj_5333, n2_adj_5334, n32195;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5335, n2_adj_5336, n2_adj_5337, n2_adj_5338, n32192, 
        n2_adj_5339, n5, n4_c, n2_adj_5340, n2_adj_5341, n2_adj_5342, 
        n2_adj_5343, n2_adj_5344, n2_adj_5345, n2_adj_5346, n2_adj_5347, 
        n2_adj_5348, n2_adj_5349, n2_adj_5350, n2_adj_5351, n2_adj_5352, 
        n2_adj_5353, n2_adj_5354, n32189, n26, n2_adj_5355, n69720, 
        n67736, n71691, n71244, n7_c;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n2_adj_5356, n2_adj_5357, n29047, n54796, n27445, n54834, 
        n71196, n71685, n2_adj_5358, n26984, Kp_23__N_767;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n28555, n71322, n7_adj_5359, n28947;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n60753, n71202, n67748, n71679, Kp_23__N_1748, n41, n31689, 
        n31690, n71292, n71646, n31691, n31692, n31696;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    
    wire n32421, n2_adj_5360, n31928, n32186, n2_adj_5361, n2_adj_5362, 
        n2_adj_5363, n32183, n2_adj_5364, n2_adj_5365, n32180, n2_adj_5366, 
        n32177, n2_adj_5367, n32174, n2_adj_5368, n2_adj_5369, n32422, 
        n2_adj_5370, n32423, n71208, n67740, n71673, n2_adj_5371, 
        n2_adj_5372, n2_adj_5373, n2_adj_5374, n2_adj_5375, n2_adj_5376, 
        n2_adj_5377, n2_adj_5378, n2_adj_5379, n2_adj_5380, n71280, 
        n71640, n2_adj_5381, n2_adj_5382, n2_adj_5383, n2_adj_5384, 
        n2_adj_5385, n2_adj_5386, n2_adj_5387, n2_adj_5388, n2_adj_5389, 
        n2_adj_5390, n2_adj_5391, n2_adj_5392, n2_adj_5393, n32424, 
        n32425, n2_adj_5394, n2_adj_5395, n2_adj_5396, n2_adj_5397, 
        n32426, n32427, n2_adj_5398, n32428, n2_adj_5399, n71214, 
        n67792, n71667, n2_adj_5400, n32429, n32430, n71238, n7_adj_5401, 
        n67666, n2_adj_5402, n32431, n9, n32432, n2_adj_5403, n31814, 
        n32433, n32434, n32435, n55740, n60685, n2_adj_5404, n12, 
        n11, n2_adj_5405, n32436, n2_adj_5406, n55956, n3, n3_adj_5407, 
        n32437, n60052, n64843, n64844, n32438, n32439, n64842, 
        n32440, n32441, n2_adj_5408, n5_adj_5409, n31324, n32442, 
        n32443, n3_adj_5410, n32494, n30094, n3_adj_5411, n32495, 
        n2081, n32496, n59365;
    wire [23:0]n4945;
    
    wire n32497, n3_adj_5412, n32498, n3_adj_5413, n71649;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n10, n14, n32499, n62849, n3_adj_5414, n32500, n30, n34, 
        n32, n33, n31, n27873, n71562, n67791, n71538, n71346, 
        n70058, n4452, \FRAME_MATCHER.i_31__N_2514 , n71643, n32501, 
        n32502, n3_adj_5415, n2_adj_5416, n3_adj_5417, n32503, n3_adj_5418;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5419, n3_adj_5420, n3_adj_5421, n3_adj_5422, n32504, 
        n32505, n32506, n60265, n60667, n10_adj_5423, n55796, n62192, 
        n32507, n55788, n60570, n55879, n60283, n3_adj_5424, n60499, 
        n12_adj_5425, n32508, n67668, n67667, n54970, n8_adj_5426, 
        n60480, n32509, n60691, n55291, n2_adj_5427, n4_adj_5428, 
        n60912, n4_adj_5429, n5_adj_5430, n71637, n60605, n2_adj_5431, 
        n32510, n3_adj_5432, n55830, n62437, n6_c, n60291, n3_adj_5433, 
        n54792, n10_adj_5434, n60417, n67669, n1_c, n60342, n59359, 
        n1_adj_5435, n60064, n1_adj_5436, n60063, n1_adj_5437, n60062, 
        n1_adj_5438, n60061, n1_adj_5439;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n60065, n60298, n55783, n60520, n60778, n6_adj_5440, n60815, 
        n55464, n26026, n60900, n28433, n60482, n54876, n61784, 
        n60427, n60596, n28441, n55273, n32511, n60918, n28170, 
        n2_adj_5441, n60153, n28070, n60154, n62880, n60441, n26_adj_5442, 
        n32512, n60876, n60374, n24, n59385, n32513, n25, n23_c, 
        n55514, n71631, n60445, n29117, n60812, n28907, n12_adj_5443, 
        n54742, n32514, n2_adj_5444, n28961, n60836, n60646, n60517, 
        n55462, n55734, n28483, n55907, n18, n60854, n20, n15_c, 
        n32515, n1522, n60485, n1513, n20_adj_5445, n62099, n55856, 
        n19, n28456, n1510, n28873, n21, n2_adj_5446;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(99[12:25])
    
    wire n32516, n2_adj_5447, n32118, n62023, n32115, n71634, n6_adj_5448, 
        n61794, n55577, n60599;
    wire [7:0]\data_in_frame[3]_c ;   // verilog/coms.v(99[12:25])
    
    wire n32517, n60335, n6_adj_5449, n30407, n30616, n53601, n67553, 
        n30405, n53600, n67554, n30403, n53599, n67555, n30401, 
        n53598, n67556, n55838, n54865, n1_adj_5450, n60060, n30399, 
        n53597, n67557, n30397, n53596, n67563, n30395, n53595, 
        n67564, n30393, n53594, n67568, n32518, n30391, n53593, 
        n67571, n1_adj_5451, n60066, n30389, n53592, n67573, n30387, 
        n53591, n67576, n30385, n53590, n67577, n30383, n53589, 
        n67578, n30381, n53588, n67579, n28056, n6_adj_5452, n30379, 
        n53587, n67609, n30377, n53586, n67610, n55744, n31799, 
        n30375, n53585, n67611, n30373, n53584, n67612, n62212, 
        n60764, n28, n54974, n32_adj_5453, n30371, n53583, n67613, 
        n30_adj_5454, n60762, n31_adj_5455, n30369, n53582, n67614, 
        n30367, n53581, n67615, n30365, n53580, n67642, n30363, 
        n53579, n67643, n29_c, n30361, n53578, n67644, n30359, 
        n53577, n67647, n30357, n53576, n67648, n10_adj_5456, n30355, 
        n53575, n67649, n30353, n53574, n67651, n60682, n8_adj_5457, 
        n30351, n53573, n67670, n71625, n71607, n71610, n71601, 
        n71604, n71595, n71598, n71589, n71592, n71583, n62281, 
        n61840, n12_adj_5458, n30349, n53572, n67693, n30347, n53571, 
        n67694, n32519;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    
    wire n26256, n20_adj_5459, n60156, n60802, Kp_23__N_1518, n30_adj_5460;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    
    wire n34_adj_5461, n60147, n54869, n32_adj_5462, n62188, n60511, 
        n60621, n33_adj_5463, n60897, n54931, n54794, n31_adj_5464, 
        n28352, n62882, n60688, n62194, n60574, n60851, n60805, 
        n27587, n29130, n60676, n6_adj_5465, n54882, n61920, n60731, 
        n60394;
    wire [7:0]\data_in_frame[18]_c ;   // verilog/coms.v(99[12:25])
    
    wire n64231, n60873, n60391, n55757, n60320, n54824, n55428, 
        n60385, n55952, n54912, n10_adj_5466, n32520;
    wire [31:0]n133;
    
    wire n161, n60162, n71586, n55932, n55903, n64159, n28548, 
        n60747, n60274, n60885, n60775, n60252, n62616, n32110, 
        n32104;
    wire [7:0]\data_in_frame[17]_c ;   // verilog/coms.v(99[12:25])
    
    wire n61788, n60535, n60784, n60587, n28505, n29167, n62765, 
        n60810, n54800, n4_adj_5467, n32521, n60245, n55864, n55754, 
        n28836, n60200, n29204, n60833, \FRAME_MATCHER.i_31__N_2507 , 
        n32101, n32098, n32095, n64131, n60302, n64135, n60624, 
        n55895, n60174, n64141, n64171, n60888, Kp_23__N_1389, n64177, 
        n32522, n60827, n60584, n64147, n32092;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    
    wire n32089, n28130, n60864, n64183, n64151, n64155, n32523, 
        n29007, n60191, n29193, n60232, n10_adj_5468, n60652, n61964, 
        n60906, n60411, n28761, n28249, n32086, n32083, n32080, 
        n32077, n55300, n32074, n32071, n60894, n28392, n64103, 
        n60673, n20_adj_5469, n26207, n55319, n19_adj_5470, n60420, 
        n21_adj_5471, n60280, n28332, Kp_23__N_974, n6_adj_5472, n32524, 
        n60591, n60462, n60756, n62109, n8_adj_5473, n71571, n11_adj_5474, 
        n55777, n28224, n13;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(246[14:26])
    
    wire n71565, n16, n60721, n60435, n17, n71250, n39176, n38177, 
        n32525, n71559, n32526, n32527, n28809, n60891, n60491, 
        n30_adj_5475, n60221, n60649, n34_adj_5476, n60882, n60528, 
        n32_adj_5477, n60368, n60277, Kp_23__N_875, n33_adj_5478, 
        n60549, n60323, n55074, n31_adj_5479, n62168, n60171, n60630, 
        n12_adj_5480, n71718, n28677, n60718, n29417, \FRAME_MATCHER.i_31__N_2508 , 
        n2061, n2062, n32002, n31999, n60694, n31996, n32528, 
        n23519, \FRAME_MATCHER.i_31__N_2511 , n58999, \FRAME_MATCHER.i_31__N_2512 , 
        n2073, n29420, n31993, n31990, n31987, n2_adj_5481, n31984, 
        n32529, n31980, n31976, n31973, n59373;
    wire [7:0]\data_in_frame[6]_c ;   // verilog/coms.v(99[12:25])
    
    wire n32530, n31969, n31966, n32531, n59379, n31962, n31959, 
        n31946, n12_adj_5482, n60773, n28122, n31955, n31952, n14_adj_5483, 
        n71274, n67738, n71553, n32532, n29303, n31283, n67624, 
        n71286, n71556, n9_adj_5484, n28299, n32533, n1_adj_5485;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n31268, n32534, n28342, n28067, Kp_23__N_1085, n32535, 
        n32536, n52833, n60058, n52832, n60314, n60561, n28228, 
        n60381, n20_adj_5486, n32537, n32538, n52831, n60432, n60796, 
        n19_adj_5487, n21_adj_5488, n52830, n52829, n52828, n52827, 
        n60059, tx_transmit_N_3416, n2_adj_5489, n2_adj_5490, n2_adj_5491, 
        n2_adj_5492, n2_adj_5493, n2_adj_5494, n2_adj_5495, n2_adj_5496, 
        n2_adj_5497, n2_adj_5498, n2_adj_5499, n2_adj_5500, n2_adj_5501, 
        n2_adj_5502, n2_adj_5503, n2_adj_5504, n2_adj_5505, n2_adj_5506, 
        n2_adj_5507, n2_adj_5508, n2_adj_5509, n2_adj_5510, n2_adj_5511, 
        n2_adj_5512, n2_adj_5513, n2_adj_5514, n2_adj_5515, n2_adj_5516, 
        n2_adj_5517, n2_adj_5518, n2_adj_5519, n2_adj_5520, n2_adj_5521, 
        n2_adj_5522, n2_adj_5523, n2_adj_5524, n2_adj_5525, n2_adj_5526, 
        n2_adj_5527, n2_adj_5528, n2_adj_5529, n2_adj_5530, n2_adj_5531, 
        n2_adj_5532, n2_adj_5533, n2_adj_5534, n2_adj_5535, n2_adj_5536, 
        n2_adj_5537, n2_adj_5538, n2_adj_5539, n2_adj_5540, n2_adj_5541, 
        n2_adj_5542, n2_adj_5543, n2_adj_5544, n2_adj_5545, n2_adj_5546, 
        n2_adj_5547, n2_adj_5548, n2_adj_5549, n2_adj_5550, n2_adj_5551, 
        n2_adj_5552, n2_adj_5553, n2_adj_5554, n2_adj_5555, n2_adj_5556, 
        n2_adj_5557, n2_adj_5558, n2_adj_5559, n31852;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n31851, n31850, n31849, n2_adj_5560, n31848, n31847, n31846, 
        n2_adj_5561, n31845;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n31844, n31843, n2_adj_5562, n31842, n31841, n31840, n2_adj_5563, 
        n31839, n31838, n31837;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n2_adj_5564, n31836, n31835, n31834, n2_adj_5565, n31833, 
        n31832, n31831, n2_adj_5566, n31830, n31829;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n31828, n31827, n31826, n31825, n2_adj_5567, n31824, n31823, 
        n31822, n2_adj_5568, n2_adj_5569, n2_adj_5570, n32539, n2_adj_5571, 
        n2_adj_5572, n55176, n60787, n32540, n32541, n32542, n62101, 
        n60361, n32543, n29250, n13_adj_5573, n30308, n11_adj_5574, 
        n60488, n62398, n55809, n32544, n60477, n29078, n60697, 
        n60271, n64121, n60670, n60311, n64095, n28812, n28337, 
        n6_adj_5575, n2_adj_5576, n32545, n32546, n32547, n60238, 
        n32548, n60184, n60203, n29044, n28742, n55607, n60377, 
        n60848, n10_adj_5577, n32549, n32550, n60473, n12_adj_5578, 
        n71535, n60767, n28213, n60494, n1_adj_5579, n32551, n32552, 
        n36, n60807, n34_adj_5580, n26_adj_5581, n40, n60262, n38, 
        n32553, n39, n37, n55793, n32554, n60921, n60602, n60759, 
        n10_adj_5582, n6_adj_5583, n27478, n10_adj_5584, n6_adj_5585, 
        n32555, n2_adj_5586, n60679, n8_adj_5587, n7_adj_5588, n60339, 
        n8_adj_5589, n32_adj_5590, n64455, n62756, n61937, n6_adj_5591, 
        n62141, n64195, n12_adj_5592;
    wire [7:0]\data_in_frame[22]_c ;   // verilog/coms.v(99[12:25])
    
    wire n64197;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n62426, n62467, n4_adj_5593, n32556, n62881, n62732, n64203, 
        n61933, n62114, n6_adj_5594, n64209, n62116, n64211, n14_adj_5595, 
        n64213, n28517, n13_adj_5596, n64217, n32557, n32558, n32559, 
        n28702, n28266, n4_adj_5597, n28782, n32560, n60308, n29010, 
        n54762, n60324, n55742, n37239, n6_adj_5598, n60459, n60227, 
        n60456, n12_adj_5599, Kp_23__N_758, n60700, Kp_23__N_872, 
        n7_adj_5600, n60845, n28690, n28157, n60332, Kp_23__N_772, 
        n60326, n28715, n60305, n12_adj_5601, n60658, n60241, n32561, 
        n60224, n32562, n32563, n60772, n32564, n32565, n60640, 
        n60197, n2_adj_5602, n62503, n6_adj_5603, n32566;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    
    wire n60821, n32567, n32568, n32569, n31683, n31686, n32222, 
        n59223, n59247, n59251, n59237, n59233, n32259, n32262, 
        n59105, n32690, n32687, n32684, n32681, n32678, n32293, 
        n59161, n32310, n32313, n59117, n32320, n32323, n32326, 
        n32329, n32332, n32335, n32338, n32341, n32344, n32347, 
        n31709, n32350, n32353, n31712, n59243, n59297, n59305, 
        n32624, n32413, n32416, n59395, n31718, n31721, n32491, 
        n59159, n31724, n31727, n31730, n24_adj_5604, n32486, n32485, 
        n32476, n32473, n32466, n32465, n32463, n2_adj_5605, n32453, 
        n59453, n79, n60259, n4_adj_5606, Kp_23__N_748, n31703, 
        n60130, n41173, n59415, n60248, n59457, n31694, n31775, 
        n31778, n59465, n28106, n64245, n64247, n64253, n64257, 
        n64261, n64269, n64267, n64085, n6_adj_5607, n6_adj_5608, 
        n5_adj_5609, n5_adj_5610, n10_adj_5611, n15_adj_5612, n14_adj_5613, 
        n22, n21_adj_5614, n23_adj_5615, n6_adj_5616, n28357, n31_adj_5617, 
        n60119, n35084, n62343, n60744, n60909, n14_adj_5618, n60531, 
        n13_adj_5619, n60739, n60405, n60452, n60879, n8_adj_5620, 
        n60858, n60643, n28968, n60830, n10_adj_5621, n60388, n28427, 
        n1699, n29148, n60709, n6_adj_5622, n60349, n60861, n60235, 
        n13_adj_5623, n55800, n12_adj_5624, n1563, n1312, n60736, 
        n60188, n60544, n71343, n10_adj_5625, n60168, n55852, n60655, 
        n60555, n60317, n60345, n29177, n46, n54859, n60818, n8_adj_5626, 
        n60209, n60712, n44, n60706, n60255, n45, n43, n60397, 
        n1130, n42, n52, n47, n41_adj_5627, n28031, n10_adj_5628, 
        n62234, n64617, n64618, n64837, n64836, n64608, n64609, 
        n64612, n60867, n60839, n64611, n64587, n64588, n64591, 
        n64590, n28024, n40_adj_5629, n14_adj_5630, n10_adj_5631, 
        n60715, n60355, n15_adj_5632, n14_adj_5633, n64899, n64900, 
        n64897, n64896, n64596, n64597, n64894, n28446, n28888, 
        n64893, n64623, n64624, n64849, n60286, n64848, n67742, 
        n64884, n64885, n64867, n64866, n64620, n64621, n28453, 
        n64861, n64828, n64862, n64827, n64797, n64798, n64630, 
        n64629, n60546, n7_adj_5634, n64860, n64792, n10_adj_5635, 
        n60567, n55840, n28745, n55769, n55750, n64791, n64793, 
        n9_adj_5636, n8_adj_5637, n60558, n62457, n29259, n10_adj_5638, 
        n60842, n28615, n40_adj_5639, n38_adj_5640, n55985, n39_adj_5641, 
        n60206, n37_adj_5642, n42_adj_5643, n46_adj_5644, n29017, 
        n41_adj_5645, n10_adj_5646, n71331, n16_adj_5647, n12_adj_5648, 
        n55732, n8_adj_5649, n60552, n7_adj_5650, n60824, n60903, 
        n60352, n60703, n62217, n14_adj_5651, n54842, n15_adj_5652, 
        n60633, n12_adj_5653, n28020, n1191, n1168, n60329, n14_adj_5654, 
        n60627, n15_adj_5655, n28697, n60268, n1964, n61999, n23514, 
        n60498, n12_adj_5656, n60915, n25071, n4_adj_5657, n14_adj_5658, 
        n9_adj_5659, n60365, n60724, n60727, n3303, n10_adj_5660, 
        n60799, n8_adj_5661, n12_adj_5662, n10_adj_5663, n60618, n10_adj_5664, 
        n1519, n1967, n1970, n64282, n1655, n60214, n62119, n60793, 
        n55179, n54978, n8_adj_5665, n6_adj_5666, n6_adj_5667, n60466, 
        n1968, n27855, n60159, n8_adj_5668, n12_adj_5669, n28824, 
        n771, n10_adj_5670, n27746, n61010, n55362, n5_adj_5672, 
        n29976, n62594, n27864, n40721, n4_adj_5673, n4_adj_5674, 
        n41206, n10_adj_5675, n14_adj_5676, n27904, n20_adj_5677, 
        n27759, n19_adj_5678, n64453, n28014, n18_adj_5679, n27913, 
        n20_adj_5680, n15_adj_5682, n10_adj_5683, n6_adj_5684, n60295, 
        n10_adj_5685, n14_adj_5686, n15_adj_5687, n16_adj_5688, n17_adj_5691, 
        n64823, n64821, n64865, n64863, n35070, n62063, n6_adj_5693, 
        n40778, n60118, n30635, n7_adj_5694, n4_adj_5695, n64822, 
        n71334, n71319, n30330, n64864, n30655, n70932, n71289, 
        n71283, n71277, n22_adj_5698, n71271, n20_adj_5699, n28_adj_5700, 
        n26_adj_5701, n25_adj_5702, n29_adj_5703, n31_adj_5704, n9_adj_5705, 
        n71247, n71241, n71235, n60135, n71211, n71205, n71199, 
        n71193;
    
    SB_LUT4 i13758_3_lut_4_lut (.I0(n30637), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n31949));
    defparam i13758_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2), .S(n59931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5316), .S(n59925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n59095));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5317), .S(n59924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32202));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5318), .S(n59923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5319), .S(n59922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5320), .S(n59921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5321), .S(n59933));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13930_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n32121));
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5322), .S(n59920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5323), .S(n59919));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5324), .S(n59918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5325), .S(n59917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5326), .S(n59916));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[4] [4]), .I1(n54798), .I2(Kp_23__N_878), 
            .I3(n60217), .O(Kp_23__N_993));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5327), .S(n59915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5328), .S(n59914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5329), .S(n59913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5330), .S(n59912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5331), .S(n59911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5332), .S(n59934));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32199));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5333), .S(n60050));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n59473));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5334), .S(n60049));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32195));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5335), .S(n60048));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5336), .S(n60047));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5337), .S(n59910));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5338), .S(n60046));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32192));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5339), .S(n59932));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_c));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5340), .S(n60045));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5341), .S(n59909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5342), .S(n59908));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5343), .S(n59907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5344), .S(n59906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5345), .S(n59905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5346), .S(n59904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5347), .S(n59903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5348), .S(n59902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5349), .S(n59901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5350), .S(n59900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5351), .S(n59899));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5352), .S(n31492));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5353), .S(n59898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5354), .S(n60044));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32189));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2887), .D(n26), .S(n31490));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5355), .S(n59897));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n69720), .I2(n67736), .I3(byte_transmit_counter[4]), .O(n71691));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71691_bdd_4_lut (.I0(n71691), .I1(n71244), .I2(n7_c), .I3(byte_transmit_counter[4]), 
            .O(tx_data[7]));
    defparam n71691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5356), .S(n59896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5357), .S(n60043));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1085 (.I0(n29047), .I1(n54796), .I2(\data_out_frame[13] [5]), 
            .I3(n27445), .O(n54834));
    defparam i2_3_lut_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52107 (.I0(byte_transmit_counter[3]), 
            .I1(n71196), .I2(n67793), .I3(byte_transmit_counter[4]), .O(n71685));
    defparam byte_transmit_counter_3__bdd_4_lut_52107.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5358), .S(n60042));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1086 (.I0(n26984), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_767), .I3(\data_in_frame[0] [7]), .O(n28555));
    defparam i2_3_lut_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 n71685_bdd_4_lut (.I0(n71685), .I1(n71322), .I2(n7_adj_5359), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n71685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1087 (.I0(n26984), .I1(\data_in_frame[2] [7]), 
            .I2(n28947), .I3(\data_in_frame[7] [4]), .O(n60753));
    defparam i2_3_lut_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52102 (.I0(byte_transmit_counter[3]), 
            .I1(n71202), .I2(n67748), .I3(byte_transmit_counter[4]), .O(n71679));
    defparam byte_transmit_counter_3__bdd_4_lut_52102.LUT_INIT = 16'he4aa;
    SB_LUT4 i13498_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n31689));   // verilog/coms.v(148[4] 304[11])
    defparam i13498_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13499_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n31690));   // verilog/coms.v(148[4] 304[11])
    defparam i13499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71679_bdd_4_lut (.I0(n71679), .I1(n71292), .I2(n71646), .I3(byte_transmit_counter[4]), 
            .O(tx_data[4]));
    defparam n71679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13500_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n31691));   // verilog/coms.v(148[4] 304[11])
    defparam i13500_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13501_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n31692));   // verilog/coms.v(148[4] 304[11])
    defparam i13501_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13505_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n31696));   // verilog/coms.v(148[4] 304[11])
    defparam i13505_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14230_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n32421));   // verilog/coms.v(148[4] 304[11])
    defparam i14230_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5360), .S(n60041));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13737_3_lut_4_lut (.I0(n30637), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n31928));
    defparam i13737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32186));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5361), .S(n60040));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5362), .S(n60039));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5363), .S(n60038));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32183));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5364), .S(n60037));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5365), .S(n59936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32180));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5366), .S(n60036));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32177));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5367), .S(n60035));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32174));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5368), .S(n60034));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32171));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5369), .S(n60033));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32168));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14231_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n32422));   // verilog/coms.v(148[4] 304[11])
    defparam i14231_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5370), .S(n60032));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32165));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14232_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n32423));   // verilog/coms.v(148[4] 304[11])
    defparam i14232_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52097 (.I0(byte_transmit_counter[3]), 
            .I1(n71208), .I2(n67740), .I3(byte_transmit_counter[4]), .O(n71673));
    defparam byte_transmit_counter_3__bdd_4_lut_52097.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5371), .S(n60031));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5372), .S(n59895));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5373), .S(n59894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5374), .S(n59893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5375), .S(n31484));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5376), .S(n59892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5377), .S(n59891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5378), .S(n59890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5379), .S(n59889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32162));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5380), .S(n60030));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n31793));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71673_bdd_4_lut (.I0(n71673), .I1(n71280), .I2(n71640), .I3(byte_transmit_counter[4]), 
            .O(tx_data[3]));
    defparam n71673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5381), .S(n60029));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32158));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5382), .S(n59888));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5383), .S(n59887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5384), .S(n59886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5385), .S(n60028));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5386), .S(n59885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5387), .S(n31475));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5388), .S(n31474));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5389), .S(n59884));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5390), .S(n59883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5391), .S(n31471));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5392), .S(n31470));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32155));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5393), .S(n59882));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14233_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n32424));   // verilog/coms.v(148[4] 304[11])
    defparam i14233_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14234_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n32425));   // verilog/coms.v(148[4] 304[11])
    defparam i14234_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5394), .S(n59881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5395), .S(n31467));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5396), .S(n59880));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5397), .S(n59879));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14235_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n32426));   // verilog/coms.v(148[4] 304[11])
    defparam i14235_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14236_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n32427));   // verilog/coms.v(148[4] 304[11])
    defparam i14236_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5398), .S(n59878));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14237_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n32428));   // verilog/coms.v(148[4] 304[11])
    defparam i14237_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5399), .S(n60027));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52092 (.I0(byte_transmit_counter[3]), 
            .I1(n71214), .I2(n67792), .I3(byte_transmit_counter[4]), .O(n71667));
    defparam byte_transmit_counter_3__bdd_4_lut_52092.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5400), .S(n59873));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14238_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n32429));   // verilog/coms.v(148[4] 304[11])
    defparam i14238_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14239_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n32430));   // verilog/coms.v(148[4] 304[11])
    defparam i14239_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71667_bdd_4_lut (.I0(n71667), .I1(n71238), .I2(n7_adj_5401), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n71667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48671_2_lut (.I0(\data_out_frame[9] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67666));
    defparam i48671_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5402), .S(n59877));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14240_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n32431));   // verilog/coms.v(148[4] 304[11])
    defparam i14240_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i9_3_lut (.I0(\data_out_frame[10] [0]), 
            .I1(\data_out_frame[11] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14241_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n32432));   // verilog/coms.v(148[4] 304[11])
    defparam i14241_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5403), .S(n31461));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13623_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n60134), 
            .I3(GND_net), .O(n31814));   // verilog/coms.v(130[12] 305[6])
    defparam i13623_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32152));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14242_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n32433));   // verilog/coms.v(148[4] 304[11])
    defparam i14242_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14243_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n32434));   // verilog/coms.v(148[4] 304[11])
    defparam i14243_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14244_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n32435));   // verilog/coms.v(148[4] 304[11])
    defparam i14244_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[24] [5]), .I1(n55740), .I2(GND_net), 
            .I3(GND_net), .O(n60685));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5404), .S(n31460));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i12_3_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\data_out_frame[15] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i11_3_lut (.I0(\data_out_frame[12] [0]), 
            .I1(\data_out_frame[13] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5405), .S(n59876));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14245_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n32436));   // verilog/coms.v(148[4] 304[11])
    defparam i14245_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5406), .S(n59875));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_212_i3_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n60514), .I3(n55956), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_212_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5407), .S(n60082));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14246_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n32437));   // verilog/coms.v(148[4] 304[11])
    defparam i14246_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1088 (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n60052));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h2222;
    SB_LUT4 i45348_3_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64843));
    defparam i45348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45349_4_lut (.I0(n64843), .I1(n60052), .I2(byte_transmit_counter[4]), 
            .I3(\data_out_frame[1][5] ), .O(n64844));
    defparam i45349_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i14247_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n32438));   // verilog/coms.v(148[4] 304[11])
    defparam i14247_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14248_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n32439));   // verilog/coms.v(148[4] 304[11])
    defparam i14248_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i45347_3_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[17] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64842));
    defparam i45347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14249_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n32440));   // verilog/coms.v(148[4] 304[11])
    defparam i14249_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32149));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14250_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n32441));   // verilog/coms.v(148[4] 304[11])
    defparam i14250_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5408), .S(n60026));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2887), .D(n5_adj_5409), 
            .S(n31324));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14251_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n32442));   // verilog/coms.v(148[4] 304[11])
    defparam i14251_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14252_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n32443));   // verilog/coms.v(148[4] 304[11])
    defparam i14252_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5410), .S(n60081));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19184_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n32494));   // verilog/coms.v(148[4] 304[11])
    defparam i19184_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16890_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(n35072), .I3(n41), .O(n30094));   // verilog/coms.v(18[27:29])
    defparam i16890_4_lut.LUT_INIT = 16'he420;
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5411), .S(n31455));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14304_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n32495));   // verilog/coms.v(148[4] 304[11])
    defparam i14304_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2081), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i14305_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n32496));   // verilog/coms.v(148[4] 304[11])
    defparam i14305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_4_lut_4_lut (.I0(n30637), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n59365));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n30094), 
            .D(n4945[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14306_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n32497));   // verilog/coms.v(148[4] 304[11])
    defparam i14306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32146));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5412), .S(n60080));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2887), .D(n3), .S(n60076));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14307_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n32498));   // verilog/coms.v(148[4] 304[11])
    defparam i14307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5413), .S(n60077));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n11), .I2(n12), .I3(byte_transmit_counter[2]), .O(n71649));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [8]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i [19]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [25]), .O(n14));   // verilog/coms.v(157[7:23])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14308_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n32499));   // verilog/coms.v(148[4] 304[11])
    defparam i14308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n14), .I2(n10), 
            .I3(\FRAME_MATCHER.i [26]), .O(n62849));   // verilog/coms.v(157[7:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5414), .S(n31451));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14309_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n32500));   // verilog/coms.v(148[4] 304[11])
    defparam i14309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_4_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [29]), .O(n30));   // verilog/coms.v(157[7:23])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n30), .I2(\FRAME_MATCHER.i [13]), 
            .I3(n62849), .O(n34));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 n71649_bdd_4_lut (.I0(n71649), .I1(n9), .I2(n67666), .I3(byte_transmit_counter[2]), 
            .O(n64802));
    defparam n71649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13_4_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [9]), .O(n32));   // verilog/coms.v(157[7:23])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i [16]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [20]), .O(n33));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [21]), .O(n31));   // verilog/coms.v(157[7:23])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n27873));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49269_2_lut (.I0(n71562), .I1(byte_transmit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n67791));
    defparam i49269_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50563_3_lut (.I0(n71538), .I1(n71346), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n70058));
    defparam i50563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22820_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27873), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i22820_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2081));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52073 (.I0(byte_transmit_counter[1]), 
            .I1(n4_c), .I2(n5), .I3(byte_transmit_counter[2]), .O(n71643));
    defparam byte_transmit_counter_1__bdd_4_lut_52073.LUT_INIT = 16'he4aa;
    SB_LUT4 i14310_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n32501));   // verilog/coms.v(148[4] 304[11])
    defparam i14310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14311_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n32502));   // verilog/coms.v(148[4] 304[11])
    defparam i14311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5415), .S(n60075));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5416), .S(n60025));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5417), .S(n60072));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14312_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n32503));   // verilog/coms.v(148[4] 304[11])
    defparam i14312_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5418), .S(n60073));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5420), .S(n31447));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32143));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5421), .S(n60078));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5422), .S(n60079));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32140));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14313_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n32504));   // verilog/coms.v(148[4] 304[11])
    defparam i14313_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14314_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n32505));   // verilog/coms.v(148[4] 304[11])
    defparam i14314_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14315_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n32506));   // verilog/coms.v(148[4] 304[11])
    defparam i14315_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut (.I0(n60265), .I1(\data_out_frame[24] [0]), .I2(\data_out_frame[24] [1]), 
            .I3(n60667), .O(n10_adj_5423));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_210_i3_4_lut (.I0(n55796), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5423), .I3(n62192), .O(n3_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i19071_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n32507));   // verilog/coms.v(148[4] 304[11])
    defparam i19071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[24] [0]), .I1(n55788), .I2(\data_out_frame[25] [7]), 
            .I3(GND_net), .O(n60570));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1089 (.I0(\data_out_frame[22] [4]), .I1(n60570), 
            .I2(n55879), .I3(GND_net), .O(n60283));
    defparam i2_3_lut_adj_1089.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5424), .S(n60071));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[19] [0]), 
            .I2(n60499), .I3(n55748), .O(n12_adj_5425));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14317_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n32508));   // verilog/coms.v(148[4] 304[11])
    defparam i14317_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n71643_bdd_4_lut (.I0(n71643), .I1(n67668), .I2(n67667), .I3(byte_transmit_counter[2]), 
            .O(n71646));
    defparam n71643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[23] [3]), .I1(n54970), .I2(n12_adj_5425), 
            .I3(n8_adj_5426), .O(n60480));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14318_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n32509));   // verilog/coms.v(148[4] 304[11])
    defparam i14318_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1090 (.I0(\data_out_frame[22] [3]), .I1(n60691), 
            .I2(\data_out_frame[22] [4]), .I3(GND_net), .O(n55291));
    defparam i2_3_lut_adj_1090.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5427), .S(n60024));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n55746), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5428));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[22] [7]), 
            .I2(\data_out_frame[20] [6]), .I3(n4_adj_5428), .O(n60912));   // verilog/coms.v(81[16:27])
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52068 (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5429), .I2(n5_adj_5430), .I3(byte_transmit_counter[2]), 
            .O(n71637));
    defparam byte_transmit_counter_1__bdd_4_lut_52068.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[21] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60605));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14319_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n32510));   // verilog/coms.v(148[4] 304[11])
    defparam i14319_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5432), .S(n31443));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1093 (.I0(\data_out_frame[20] [0]), .I1(n55830), 
            .I2(n62437), .I3(n6_c), .O(n60291));
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(\data_out_frame[21] [5]), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[21] [6]), .I3(GND_net), .O(n60667));
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2887), .D(n3_adj_5433), .S(n60074));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1095 (.I0(n54792), .I1(\data_out_frame[22] [1]), 
            .I2(\data_out_frame[21] [7]), .I3(n60291), .O(n10_adj_5434));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n60417), .I1(n10_adj_5434), .I2(n55879), .I3(GND_net), 
            .O(n60414));
    defparam i5_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 n71637_bdd_4_lut (.I0(n71637), .I1(n67669), .I2(n1_c), .I3(byte_transmit_counter[2]), 
            .O(n71640));
    defparam n71637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60342));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_4_lut_adj_1097 (.I0(n30637), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n59359));
    defparam i11_4_lut_4_lut_adj_1097.LUT_INIT = 16'hfe10;
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5435), .S(n60064));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5436), .S(n60063));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5437), .S(n60062));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5438), .S(n60061));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2887), .D(n1_adj_5439), .S(n60065));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1098 (.I0(n55760), .I1(n60298), .I2(\data_out_frame[19] [7]), 
            .I3(GND_net), .O(n60691));
    defparam i2_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_out_frame[16] [0]), .I1(n55783), 
            .I2(GND_net), .I3(GND_net), .O(n60520));
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1100 (.I0(n27445), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n60778));
    defparam i2_3_lut_adj_1100.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5440));
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1102 (.I0(n60778), .I1(n60520), .I2(n60815), 
            .I3(n6_adj_5440), .O(n60523));
    defparam i4_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(n55464), .I1(n60523), .I2(GND_net), 
            .I3(GND_net), .O(n26026));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1104 (.I0(\data_out_frame[16] [4]), .I1(n60900), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n28433));
    defparam i2_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1105 (.I0(n28433), .I1(n60482), .I2(n54876), 
            .I3(GND_net), .O(n61784));
    defparam i2_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1106 (.I0(n60427), .I1(n60596), .I2(n28441), 
            .I3(GND_net), .O(n55273));
    defparam i2_3_lut_adj_1106.LUT_INIT = 16'h9696;
    SB_LUT4 i14320_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n32511));   // verilog/coms.v(148[4] 304[11])
    defparam i14320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1107 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n60918));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28170));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1109 (.I0(n60153), .I1(\data_out_frame[18] [0]), 
            .I2(n55830), .I3(GND_net), .O(n60298));
    defparam i2_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(n28070), .I1(\data_out_frame[17] [5]), .I2(\data_out_frame[17] [7]), 
            .I3(n60154), .O(n62880));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1110 (.I0(n28170), .I1(n60918), .I2(\data_out_frame[14] [3]), 
            .I3(n60441), .O(n26_adj_5442));
    defparam i11_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i14321_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n32512));   // verilog/coms.v(148[4] 304[11])
    defparam i14321_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9_4_lut (.I0(n60876), .I1(\data_out_frame[19] [4]), .I2(n62880), 
            .I3(n60374), .O(n24));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_4_lut_adj_1111 (.I0(n30637), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n59385));
    defparam i11_4_lut_4_lut_adj_1111.LUT_INIT = 16'hfe10;
    SB_LUT4 i14322_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n32513));   // verilog/coms.v(148[4] 304[11])
    defparam i14322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[17] [3]), .I3(\data_out_frame[18] [5]), 
            .O(n25));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1112 (.I0(n23_c), .I1(n25), .I2(n24), .I3(n26_adj_5442), 
            .O(n55514));
    defparam i14_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n71631));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1113 (.I0(n55514), .I1(n60445), .I2(n29117), 
            .I3(GND_net), .O(n60812));
    defparam i2_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1114 (.I0(\data_out_frame[19] [5]), .I1(n60427), 
            .I2(n28907), .I3(n60812), .O(n12_adj_5443));
    defparam i5_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1115 (.I0(n55781), .I1(n12_adj_5443), .I2(n60900), 
            .I3(\data_out_frame[17] [0]), .O(n54742));
    defparam i6_4_lut_adj_1115.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32137));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14323_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n32514));   // verilog/coms.v(148[4] 304[11])
    defparam i14323_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32134));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_out_frame[18] [4]), .I1(n55273), 
            .I2(GND_net), .I3(GND_net), .O(n60150));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n31796));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5444), .S(n60023));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32130));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32127));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1117 (.I0(n28961), .I1(n60417), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n54876));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1118 (.I0(n62437), .I1(n60836), .I2(n60646), 
            .I3(n60517), .O(n55462));
    defparam i3_4_lut_adj_1118.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(n55462), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55734));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32124));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1120 (.I0(n28483), .I1(n54876), .I2(n55267), 
            .I3(n55907), .O(n18));
    defparam i7_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1121 (.I0(n54792), .I1(n18), .I2(n26026), .I3(n60854), 
            .O(n20));
    defparam i9_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1122 (.I0(n15_c), .I1(n20), .I2(n55737), .I3(\data_out_frame[22] [1]), 
            .O(n55956));
    defparam i10_4_lut_adj_1122.LUT_INIT = 16'h9669;
    SB_LUT4 i14324_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n32515));   // verilog/coms.v(148[4] 304[11])
    defparam i14324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8_4_lut (.I0(n1522), .I1(n60485), .I2(n1513), .I3(n54796), 
            .O(n20_adj_5445));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1123 (.I0(\data_out_frame[12] [0]), .I1(n62099), 
            .I2(\data_out_frame[14] [1]), .I3(n55856), .O(n19));
    defparam i7_4_lut_adj_1123.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1124 (.I0(n28456), .I1(\data_out_frame[13] [7]), 
            .I2(n1510), .I3(n28873), .O(n21));
    defparam i9_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5446), .S(n60022));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32121));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14325_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2]_c [0]), 
            .I3(\Kp[8] ), .O(n32516));   // verilog/coms.v(148[4] 304[11])
    defparam i14325_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5447), .S(n60021));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32118));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19), .I2(n20_adj_5445), .I3(GND_net), 
            .O(n62023));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32115));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71631_bdd_4_lut (.I0(n71631), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n71634));
    defparam n71631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1125 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(n62023), .I3(n6_adj_5448), .O(n61794));
    defparam i4_4_lut_adj_1125.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[15] [6]), .I1(n55577), 
            .I2(GND_net), .I3(GND_net), .O(n60599));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i14326_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [7]), 
            .I3(\Kp[7] ), .O(n32517));   // verilog/coms.v(148[4] 304[11])
    defparam i14326_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1127 (.I0(\data_out_frame[18] [2]), .I1(n60335), 
            .I2(n60599), .I3(n6_adj_5449), .O(n55464));
    defparam i4_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_33_lut  (.I0(n67553), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n53601), .O(n30407)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_32_lut  (.I0(n67554), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n53600), .O(n30405)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_32  (.CI(n53600), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n53601));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_31_lut  (.I0(n67555), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n53599), .O(n30403)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_31  (.CI(n53599), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n53600));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_30_lut  (.I0(n67556), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n53598), .O(n30401)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_30  (.CI(n53598), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n53599));
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[18] [3]), .I1(n61794), 
            .I2(GND_net), .I3(GND_net), .O(n55838));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_out_frame[20] [4]), .I1(n28483), 
            .I2(GND_net), .I3(GND_net), .O(n54865));
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2887), .D(n1_adj_5450), .S(n60060));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_29_lut  (.I0(n67557), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n53597), .O(n30399)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_29  (.CI(n53597), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n53598));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_28_lut  (.I0(n67563), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n53596), .O(n30397)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_28  (.CI(n53596), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n53597));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_27_lut  (.I0(n67564), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n53595), .O(n30395)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_27  (.CI(n53595), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n53596));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_26_lut  (.I0(n67568), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n53594), .O(n30393)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i19420_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [6]), 
            .I3(\Kp[6] ), .O(n32518));   // verilog/coms.v(148[4] 304[11])
    defparam i19420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_26  (.CI(n53594), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n53595));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_25_lut  (.I0(n67571), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n53593), .O(n30391)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_25  (.CI(n53593), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n53594));
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2887), .D(n1_adj_5451), .S(n60066));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_24_lut  (.I0(n67573), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n53592), .O(n30389)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_24  (.CI(n53592), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n53593));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_23_lut  (.I0(n67576), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n53591), .O(n30387)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_23  (.CI(n53591), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n53592));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_22_lut  (.I0(n67577), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n53590), .O(n30385)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_22  (.CI(n53590), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n53591));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_21_lut  (.I0(n67578), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n53589), .O(n30383)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_21  (.CI(n53589), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n53590));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_20_lut  (.I0(n67579), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n53588), .O(n30381)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(n28056), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5452));
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_20  (.CI(n53588), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n53589));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_19_lut  (.I0(n67609), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n53587), .O(n30379)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_19  (.CI(n53587), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n53588));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_18_lut  (.I0(n67610), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n53586), .O(n30377)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(\data_out_frame[17] [4]), .I1(n55744), 
            .I2(\data_out_frame[15] [3]), .I3(n6_adj_5452), .O(n62437));
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n31799));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_18  (.CI(n53586), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n53587));
    SB_LUT4 i3_4_lut_adj_1132 (.I0(n62437), .I1(\data_out_frame[22] [0]), 
            .I2(\data_out_frame[19] [6]), .I3(n60154), .O(n60854));
    defparam i3_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_17_lut  (.I0(n67611), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n53585), .O(n30375)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_17  (.CI(n53585), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n53586));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_16_lut  (.I0(n67612), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n53584), .O(n30373)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_16  (.CI(n53584), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n53585));
    SB_LUT4 i3_4_lut_adj_1133 (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[24] [3]), 
            .I2(\data_out_frame[23] [1]), .I3(n54865), .O(n62212));
    defparam i3_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1134 (.I0(\data_out_frame[20] [1]), .I1(n62212), 
            .I2(n60764), .I3(\data_out_frame[24] [4]), .O(n28));
    defparam i10_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(n60854), .I1(n28), .I2(n54974), .I3(GND_net), 
            .O(n32_adj_5453));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_15_lut  (.I0(n67613), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n53583), .O(n30371)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i12_4_lut_adj_1135 (.I0(n60342), .I1(\data_out_frame[23] [0]), 
            .I2(n60414), .I3(n60667), .O(n30_adj_5454));
    defparam i12_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_15  (.CI(n53583), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n53584));
    SB_LUT4 i13_4_lut_adj_1136 (.I0(n60605), .I1(n60912), .I2(n60762), 
            .I3(\data_out_frame[24] [6]), .O(n31_adj_5455));
    defparam i13_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_14_lut  (.I0(n67614), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n53582), .O(n30369)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_14  (.CI(n53582), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n53583));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_13_lut  (.I0(n67615), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n53581), .O(n30367)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_13  (.CI(n53581), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n53582));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_12_lut  (.I0(n67642), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n53580), .O(n30365)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_12  (.CI(n53580), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n53581));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_11_lut  (.I0(n67643), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n53579), .O(n30363)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_11  (.CI(n53579), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n53580));
    SB_LUT4 i11_4_lut_adj_1137 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[23] [7]), 
            .I2(n55291), .I3(n60480), .O(n29_c));
    defparam i11_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_10_lut  (.I0(n67644), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n53578), .O(n30361)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_10  (.CI(n53578), .I0(n30616), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n53579));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_9_lut  (.I0(n67647), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n53577), .O(n30359)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_9  (.CI(n53577), .I0(n30616), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n53578));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_8_lut  (.I0(n67648), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n53576), .O(n30357)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i17_4_lut (.I0(n29_c), .I1(n31_adj_5455), .I2(n30_adj_5454), 
            .I3(n32_adj_5453), .O(n55788));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1138 (.I0(n55956), .I1(n60265), .I2(n55734), 
            .I3(\data_out_frame[23] [7]), .O(n10_adj_5456));
    defparam i4_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_8  (.CI(n53576), .I0(n30616), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n53577));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_7_lut  (.I0(n67649), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n53575), .O(n30355)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_7  (.CI(n53575), .I0(n30616), .I1(\FRAME_MATCHER.i [5]), 
            .CO(n53576));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_6_lut  (.I0(n67651), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n53574), .O(n30353)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_6  (.CI(n53574), .I0(n30616), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n53575));
    SB_LUT4 i1_2_lut_adj_1139 (.I0(n60682), .I1(n55788), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5457));
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_5_lut  (.I0(n67670), .I1(n30616), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n53573), .O(n30351)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_5  (.CI(n53573), .I0(n30616), .I1(\FRAME_MATCHER.i [3]), 
            .CO(n53574));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52058 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n71625));
    defparam byte_transmit_counter_0__bdd_4_lut_52058.LUT_INIT = 16'he4aa;
    SB_LUT4 n71625_bdd_4_lut (.I0(n71625), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n71628));
    defparam n71625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52053 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71607));
    defparam byte_transmit_counter_0__bdd_4_lut_52053.LUT_INIT = 16'he4aa;
    SB_LUT4 n71607_bdd_4_lut (.I0(n71607), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71610));
    defparam n71607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52038 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n71601));
    defparam byte_transmit_counter_0__bdd_4_lut_52038.LUT_INIT = 16'he4aa;
    SB_LUT4 n71601_bdd_4_lut (.I0(n71601), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n71604));
    defparam n71601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52033 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n71595));
    defparam byte_transmit_counter_0__bdd_4_lut_52033.LUT_INIT = 16'he4aa;
    SB_LUT4 n71595_bdd_4_lut (.I0(n71595), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71598));
    defparam n71595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52028 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n71589));
    defparam byte_transmit_counter_0__bdd_4_lut_52028.LUT_INIT = 16'he4aa;
    SB_LUT4 n71589_bdd_4_lut (.I0(n71589), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8][2] ), .I3(byte_transmit_counter[1]), 
            .O(n71592));
    defparam n71589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52023 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n71583));
    defparam byte_transmit_counter_0__bdd_4_lut_52023.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_4_lut_adj_1140 (.I0(n62281), .I1(n60283), .I2(n61840), 
            .I3(n60762), .O(n12_adj_5458));
    defparam i5_4_lut_adj_1140.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_209_i3_4_lut (.I0(n55740), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5458), .I3(n8_adj_5457), .O(n3_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_4_lut  (.I0(n67693), .I1(n30616), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n53572), .O(n30349)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_4  (.CI(n53572), .I0(n30616), .I1(\FRAME_MATCHER.i[2] ), 
            .CO(n53573));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_3_lut  (.I0(n67694), .I1(n30616), 
            .I2(\FRAME_MATCHER.i[1] ), .I3(n53571), .O(n30347)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_3  (.CI(n53571), .I0(n30616), .I1(\FRAME_MATCHER.i[1] ), 
            .CO(n53572));
    SB_LUT4 i14328_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3][5] ), 
            .I3(\Kp[5] ), .O(n32519));   // verilog/coms.v(148[4] 304[11])
    defparam i14328_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[21] [6]), .I1(n26256), .I2(\data_in_frame[21][7] ), 
            .I3(GND_net), .O(n20_adj_5459));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1141 (.I0(n60156), .I1(\data_in_frame[17] [7]), 
            .I2(n60802), .I3(Kp_23__N_1518), .O(n30_adj_5460));
    defparam i11_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1142 (.I0(\data_in_frame[19] [7]), .I1(n30_adj_5460), 
            .I2(n20_adj_5459), .I3(\data_in_frame[20] [0]), .O(n34_adj_5461));
    defparam i15_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1143 (.I0(\data_in_frame[16] [3]), .I1(n60147), 
            .I2(\data_in_frame[18] [6]), .I3(n54869), .O(n32_adj_5462));
    defparam i13_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1144 (.I0(n62188), .I1(n60511), .I2(\data_in_frame[20] [1]), 
            .I3(n60621), .O(n33_adj_5463));
    defparam i14_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1145 (.I0(n60897), .I1(\data_in_frame[20] [7]), 
            .I2(n54931), .I3(n54794), .O(n31_adj_5464));
    defparam i12_4_lut_adj_1145.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1146 (.I0(\data_in_frame[21][1] ), .I1(\data_in_frame[21][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n28352));
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h6666;
    SB_LUT4 i18_4_lut_adj_1147 (.I0(n31_adj_5464), .I1(n33_adj_5463), .I2(n32_adj_5462), 
            .I3(n34_adj_5461), .O(n62882));
    defparam i18_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1148 (.I0(n62882), .I1(n28352), .I2(n26256), 
            .I3(n60688), .O(n62194));
    defparam i3_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1149 (.I0(n60574), .I1(\data_in_frame[21][4] ), 
            .I2(n62194), .I3(n60851), .O(n60805));
    defparam i2_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1150 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[20] [6]), 
            .I2(n27587), .I3(n29130), .O(n60156));
    defparam i3_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1151 (.I0(\data_in_frame[21][0] ), .I1(n60156), 
            .I2(n60676), .I3(n6_adj_5465), .O(n54882));
    defparam i4_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_in_frame[18] [2]), .I1(n61920), 
            .I2(GND_net), .I3(GND_net), .O(n60731));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(n27587), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60394));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1154 (.I0(n60394), .I1(\data_in_frame[18]_c [4]), 
            .I2(\data_in_frame[18][7] ), .I3(\data_in_frame[20] [7]), .O(n64231));
    defparam i1_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1155 (.I0(n60873), .I1(n60731), .I2(n60391), 
            .I3(n64231), .O(n55757));
    defparam i1_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(\data_in_frame[14] [6]), .I1(n60320), 
            .I2(n54824), .I3(n55428), .O(n29130));
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(n60385), .I1(\data_in_frame[19] [0]), 
            .I2(n29130), .I3(GND_net), .O(n60391));
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(n55952), .I1(n54912), .I2(GND_net), 
            .I3(GND_net), .O(n60574));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1159 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[18][7] ), 
            .I2(\data_in_frame[19] [1]), .I3(\data_in_frame[16] [6]), .O(n10_adj_5466));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i14329_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [4]), 
            .I3(\Kp[4] ), .O(n32520));   // verilog/coms.v(148[4] 304[11])
    defparam i14329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1160 (.I0(n60162), .I1(\data_in_frame[21][3] ), 
            .I2(n54869), .I3(GND_net), .O(n54912));
    defparam i2_3_lut_adj_1160.LUT_INIT = 16'h9696;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n53571));
    SB_LUT4 n71583_bdd_4_lut (.I0(n71583), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n71586));
    defparam n71583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1161 (.I0(n55932), .I1(Kp_23__N_1518), .I2(n55903), 
            .I3(n64159), .O(n60873));
    defparam i1_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1162 (.I0(n28548), .I1(n60873), .I2(n60747), 
            .I3(GND_net), .O(n60274));
    defparam i1_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1163 (.I0(\data_in_frame[13] [1]), .I1(n60885), 
            .I2(n60775), .I3(n60252), .O(n55932));
    defparam i3_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1164 (.I0(n55932), .I1(n62188), .I2(n55903), 
            .I3(\data_in_frame[17] [5]), .O(n62616));
    defparam i1_4_lut_adj_1164.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n31802));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32110));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32104));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1165 (.I0(\data_in_frame[17]_c [1]), .I1(n61788), 
            .I2(n60535), .I3(n60784), .O(n60587));
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(n62616), .I1(n28505), .I2(GND_net), 
            .I3(GND_net), .O(n29167));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(n62765), .I1(n60587), .I2(GND_net), 
            .I3(GND_net), .O(n60810));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1168 (.I0(\data_in_frame[16] [7]), .I1(n54800), 
            .I2(\data_in_frame[12] [4]), .I3(n4_adj_5467), .O(n60320));
    defparam i1_4_lut_adj_1168.LUT_INIT = 16'h9669;
    SB_LUT4 i14330_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3][3] ), 
            .I3(\Kp[3] ), .O(n32521));   // verilog/coms.v(148[4] 304[11])
    defparam i14330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1169 (.I0(n60245), .I1(n60320), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n55428));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(n55428), .I1(\data_in_frame[17]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n55864));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60784));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_in_frame[15] [5]), .I1(n55754), 
            .I2(GND_net), .I3(GND_net), .O(n60511));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1173 (.I0(n28836), .I1(n60200), .I2(n29204), 
            .I3(\data_in_frame[12] [4]), .O(n54824));
    defparam i3_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(n54824), .I1(n28548), .I2(GND_net), 
            .I3(GND_net), .O(n60833));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i48708_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67694));   // verilog/coms.v(158[12:15])
    defparam i48708_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32101));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32098));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32095));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i49178_2_lut (.I0(\FRAME_MATCHER.i[2] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67693));   // verilog/coms.v(158[12:15])
    defparam i49178_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60200));
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1176 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n64131));
    defparam i1_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1177 (.I0(n64131), .I1(n60302), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[15] [4]), .O(n64135));
    defparam i1_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1178 (.I0(n60624), .I1(n55895), .I2(n60174), 
            .I3(n64135), .O(n64141));
    defparam i1_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1179 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[15] [7]), .O(n64171));
    defparam i1_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1180 (.I0(n60888), .I1(n60784), .I2(Kp_23__N_1389), 
            .I3(n64171), .O(n64177));
    defparam i1_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i14331_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [2]), 
            .I3(\Kp[2] ), .O(n32522));   // verilog/coms.v(148[4] 304[11])
    defparam i14331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1181 (.I0(n60827), .I1(n60245), .I2(n60584), 
            .I3(n64141), .O(n64147));
    defparam i1_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i48697_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67670));   // verilog/coms.v(158[12:15])
    defparam i48697_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32092));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32089));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1182 (.I0(n28130), .I1(n60833), .I2(n60864), 
            .I3(n64177), .O(n64183));
    defparam i1_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1183 (.I0(n27587), .I1(n64151), .I2(n55864), 
            .I3(n64147), .O(n64155));
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1184 (.I0(n60810), .I1(n64155), .I2(n64183), 
            .I3(n29167), .O(Kp_23__N_1518));
    defparam i1_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i48628_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67651));   // verilog/coms.v(158[12:15])
    defparam i48628_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14332_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [1]), 
            .I3(\Kp[1] ), .O(n32523));   // verilog/coms.v(148[4] 304[11])
    defparam i14332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5441), .S(n60020));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[18][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n29007));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1186 (.I0(n60191), .I1(n29193), .I2(\data_in_frame[14] [3]), 
            .I3(n60232), .O(n10_adj_5468));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1187 (.I0(n60652), .I1(n10_adj_5468), .I2(n61964), 
            .I3(GND_net), .O(n60906));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_adj_1187.LUT_INIT = 16'h6969;
    SB_LUT4 i48626_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67649));   // verilog/coms.v(158[12:15])
    defparam i48626_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5431), .S(n60019));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1188 (.I0(\data_in_frame[9] [7]), .I1(n60411), 
            .I2(n28761), .I3(n28249), .O(n29204));
    defparam i3_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32086));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1189 (.I0(n29204), .I1(n60906), .I2(\data_in_frame[12] [2]), 
            .I3(GND_net), .O(n28548));
    defparam i2_3_lut_adj_1189.LUT_INIT = 16'h9696;
    SB_LUT4 i48625_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67648));   // verilog/coms.v(158[12:15])
    defparam i48625_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[12] [2]), .I1(n54800), 
            .I2(GND_net), .I3(GND_net), .O(n60584));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i48623_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67647));   // verilog/coms.v(158[12:15])
    defparam i48623_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32083));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32080));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48621_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67644));   // verilog/coms.v(158[12:15])
    defparam i48621_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48620_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67643));   // verilog/coms.v(158[12:15])
    defparam i48620_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32077));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1191 (.I0(n55300), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60775));
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32074));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32071));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1192 (.I0(n60894), .I1(n60775), .I2(n28392), 
            .I3(n64103), .O(n62188));
    defparam i1_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1193 (.I0(n60673), .I1(n60676), .I2(n60747), 
            .I3(n60385), .O(n20_adj_5469));
    defparam i8_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i48414_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67642));   // verilog/coms.v(158[12:15])
    defparam i48414_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1194 (.I0(n26207), .I1(n55319), .I2(\data_in_frame[20] [1]), 
            .I3(n29007), .O(n19_adj_5470));
    defparam i7_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1195 (.I0(n27587), .I1(n61920), .I2(Kp_23__N_1518), 
            .I3(n60420), .O(n21_adj_5471));
    defparam i9_4_lut_adj_1195.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32068));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i11_3_lut_adj_1196 (.I0(n21_adj_5471), .I1(n19_adj_5470), .I2(n20_adj_5469), 
            .I3(GND_net), .O(n60280));
    defparam i11_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_LUT4 i48603_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67615));   // verilog/coms.v(158[12:15])
    defparam i48603_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48602_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67614));   // verilog/coms.v(158[12:15])
    defparam i48602_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n28332), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60864));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1198 (.I0(\data_in_frame[11] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[8] [6]), .I3(n6_adj_5472), .O(n60894));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i48601_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67613));   // verilog/coms.v(158[12:15])
    defparam i48601_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32065));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14333_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n32524));   // verilog/coms.v(148[4] 304[11])
    defparam i14333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[15] [1]), .I1(n28392), 
            .I2(GND_net), .I3(GND_net), .O(n60591));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32062));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48600_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67612));   // verilog/coms.v(158[12:15])
    defparam i48600_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(n60462), .I1(n60756), .I2(\data_in_frame[14] [7]), 
            .I3(GND_net), .O(n62109));
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[17]_c [2]), 
            .I2(n62109), .I3(GND_net), .O(n8_adj_5473));
    defparam i3_3_lut.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5419), .S(n60018));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48599_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67611));   // verilog/coms.v(158[12:15])
    defparam i48599_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52013 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[0]), .O(n71571));
    defparam byte_transmit_counter_1__bdd_4_lut_52013.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1201 (.I0(n60756), .I1(\data_in_frame[14] [6]), 
            .I2(n8_adj_5473), .I3(n60885), .O(n11_adj_5474));
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1202 (.I0(\data_in_frame[12] [6]), .I1(n60591), 
            .I2(n55777), .I3(n28224), .O(n13));
    defparam i5_4_lut_adj_1202.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1203 (.I0(n13), .I1(n11_adj_5474), .I2(\data_in_frame[15] [0]), 
            .I3(\data_in_frame[14] [7]), .O(n62765));
    defparam i7_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 n71571_bdd_4_lut (.I0(n71571), .I1(\data_out_frame[26] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[0]), 
            .O(n71574));
    defparam n71571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1204 (.I0(control_mode[4]), .I1(control_mode[5]), 
            .I2(control_mode_c[3]), .I3(control_mode_c[2]), .O(n62692));
    defparam i1_4_lut_adj_1204.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52087 (.I0(byte_transmit_counter[3]), 
            .I1(n70058), .I2(n67791), .I3(byte_transmit_counter[2]), .O(n71565));
    defparam byte_transmit_counter_3__bdd_4_lut_52087.LUT_INIT = 16'he4aa;
    SB_LUT4 i13608_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n30673), 
            .I3(GND_net), .O(n31799));   // verilog/coms.v(130[12] 305[6])
    defparam i13608_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48598_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67610));   // verilog/coms.v(158[12:15])
    defparam i48598_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1205 (.I0(n55895), .I1(\data_in_frame[17]_c [3]), 
            .I2(n60864), .I3(n60591), .O(n16));
    defparam i6_4_lut_adj_1205.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32059));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32056));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1206 (.I0(n55754), .I1(n60721), .I2(n60894), 
            .I3(n60435), .O(n17));
    defparam i7_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32053));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32050));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48356_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67609));   // verilog/coms.v(158[12:15])
    defparam i48356_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32047));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32044));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n32041));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32038));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n31806));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71565_bdd_4_lut (.I0(n71565), .I1(n71250), .I2(n39176), .I3(byte_transmit_counter[2]), 
            .O(tx_data[5]));
    defparam n71565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_1207 (.I0(\control_mode[6] ), .I1(n62692), .I2(\control_mode[7] ), 
            .I3(GND_net), .O(n38177));
    defparam i1_3_lut_adj_1207.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut_adj_1208 (.I0(n17), .I1(n55300), .I2(n16), .I3(n62109), 
            .O(n28505));
    defparam i9_4_lut_adj_1208.LUT_INIT = 16'h9669;
    SB_LUT4 i14334_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n32525));   // verilog/coms.v(148[4] 304[11])
    defparam i14334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n31811));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n31814));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n31853));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n31916));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n31919));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n31922));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n31925));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
           .D(n31928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n30094), 
            .D(n4945[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_52018 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n71559));
    defparam byte_transmit_counter_0__bdd_4_lut_52018.LUT_INIT = 16'he4aa;
    SB_LUT4 i14335_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n32526));   // verilog/coms.v(148[4] 304[11])
    defparam i14335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n30094), 
            .D(n4945[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n30094), 
            .D(n4945[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n30094), 
            .D(n4945[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n30094), 
            .D(n4945[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n30094), 
            .D(n4945[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14336_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n32527));   // verilog/coms.v(148[4] 304[11])
    defparam i14336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n30094), 
            .D(n4945[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n30094), 
            .D(n4945[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n30094), 
            .D(n4945[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n30094), 
            .D(n4945[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n30094), 
            .D(n4945[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n30094), 
            .D(n4945[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n30094), 
            .D(n4945[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n30094), 
            .D(n4945[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n30094), 
            .D(n4945[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n30094), 
            .D(n4945[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n30094), 
            .D(n4945[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n30094), 
            .D(n4945[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n30094), 
            .D(n4945[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n30094), 
            .D(n4945[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n30094), 
            .D(n4945[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n30094), 
            .D(n4945[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n30094), 
            .D(n4945[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32018));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1209 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n60652));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(n28809), .I1(\data_in_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60624));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1211 (.I0(n60891), .I1(\data_in_frame[9] [0]), 
            .I2(n60491), .I3(n60753), .O(n30_adj_5475));
    defparam i11_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32015));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15_4_lut_adj_1212 (.I0(\data_in_frame[5] [1]), .I1(n30_adj_5475), 
            .I2(n60221), .I3(n60649), .O(n34_adj_5476));
    defparam i15_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1213 (.I0(n60882), .I1(n60609), .I2(n60652), 
            .I3(n60528), .O(n32_adj_5477));
    defparam i13_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 n71559_bdd_4_lut (.I0(n71559), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71562));
    defparam n71559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32012));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32009));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48497_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67579));   // verilog/coms.v(158[12:15])
    defparam i48497_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14_4_lut_adj_1214 (.I0(n60368), .I1(\data_in_frame[8] [6]), 
            .I2(n60277), .I3(Kp_23__N_875), .O(n33_adj_5478));
    defparam i14_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1215 (.I0(n60549), .I1(\data_in_frame[6] [3]), 
            .I2(n60323), .I3(n55074), .O(n31_adj_5479));
    defparam i12_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n59365));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i18_4_lut_adj_1216 (.I0(n31_adj_5479), .I1(n33_adj_5478), .I2(n32_adj_5477), 
            .I3(n34_adj_5476), .O(n62168));
    defparam i18_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1217 (.I0(n60171), .I1(n60630), .I2(\data_in_frame[13] [3]), 
            .I3(\data_in_frame[13] [1]), .O(n12_adj_5480));
    defparam i5_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n32005));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n71718), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i6_4_lut_adj_1218 (.I0(n28677), .I1(n12_adj_5480), .I2(n60718), 
            .I3(\data_in_frame[16] [0]), .O(n26207));
    defparam i6_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n29417), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2061), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2062), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n32002));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31999));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1219 (.I0(\data_in_frame[14] [2]), .I1(n62168), 
            .I2(n28677), .I3(GND_net), .O(n60694));
    defparam i2_3_lut_adj_1219.LUT_INIT = 16'h6969;
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31996));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14337_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n32528));   // verilog/coms.v(148[4] 304[11])
    defparam i14337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n23519), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n58999), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2073), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n29420), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31993));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31990));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5481), .S(n60017));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31984));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n59359));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14338_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n32529));   // verilog/coms.v(148[4] 304[11])
    defparam i14338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31980));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n59385));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n31973));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60302));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6]_c [4]), .C(clk16MHz), 
           .D(n59373));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14339_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n32530));   // verilog/coms.v(148[4] 304[11])
    defparam i14339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n31969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n31966));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48496_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67578));   // verilog/coms.v(158[12:15])
    defparam i48496_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14340_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n32531));   // verilog/coms.v(148[4] 304[11])
    defparam i14340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6]_c [5]), .C(clk16MHz), 
           .D(n59379));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48495_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67577));   // verilog/coms.v(158[12:15])
    defparam i48495_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n31962));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n31959));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48486_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67576));   // verilog/coms.v(158[12:15])
    defparam i48486_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6][6] ), .C(clk16MHz), 
           .D(n31946));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60252));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1222 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[15] [6]), .I3(n28332), .O(n12_adj_5482));   // verilog/coms.v(78[16:43])
    defparam i5_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1223 (.I0(n60773), .I1(n12_adj_5482), .I2(n28122), 
            .I3(\data_in_frame[13] [5]), .O(n60171));   // verilog/coms.v(78[16:43])
    defparam i6_4_lut_adj_1223.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n31955));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17][6] ), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1224 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[18][0] ), 
            .I2(n60171), .I3(\data_in_frame[13] [4]), .O(n60897));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n31952));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1225 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(n60252), .I3(\data_in_frame[13] [3]), .O(n14_adj_5483));
    defparam i6_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_52003 (.I0(byte_transmit_counter[3]), 
            .I1(n71274), .I2(n67738), .I3(byte_transmit_counter[1]), .O(n71553));
    defparam byte_transmit_counter_3__bdd_4_lut_52003.LUT_INIT = 16'he4aa;
    SB_LUT4 i14341_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n32532));   // verilog/coms.v(148[4] 304[11])
    defparam i14341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2887), .D(n29303), 
            .S(n31283));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n71553_bdd_4_lut (.I0(n71553), .I1(n67624), .I2(n71286), .I3(byte_transmit_counter[1]), 
            .O(n71556));
    defparam n71553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1226 (.I0(n9_adj_5484), .I1(n14_adj_5483), .I2(n60773), 
            .I3(n28299), .O(n55903));
    defparam i7_4_lut_adj_1226.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n31949));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14342_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n32533));   // verilog/coms.v(148[4] 304[11])
    defparam i14342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5485), .S(n31268));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14343_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n32534));   // verilog/coms.v(148[4] 304[11])
    defparam i14343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1227 (.I0(n28342), .I1(n28067), .I2(n60232), 
            .I3(Kp_23__N_1085), .O(n60277));
    defparam i1_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i14344_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n32535));   // verilog/coms.v(148[4] 304[11])
    defparam i14344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14345_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n32536));   // verilog/coms.v(148[4] 304[11])
    defparam i14345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(n60277), .I1(\data_in_frame[11] [7]), 
            .I2(n61964), .I3(GND_net), .O(n60191));
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h6969;
    SB_LUT4 add_1194_9_lut (.I0(n60058), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n52833), .O(n60066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1194_8_lut (.I0(n60058), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n52832), .O(n60060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1229 (.I0(n60314), .I1(n60561), .I2(n28228), 
            .I3(n60381), .O(n20_adj_5486));
    defparam i8_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_CARRY add_1194_8 (.CI(n52832), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n52833));
    SB_LUT4 i14346_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n32537));   // verilog/coms.v(148[4] 304[11])
    defparam i14346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14347_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n32538));   // verilog/coms.v(148[4] 304[11])
    defparam i14347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_1194_7_lut (.I0(n60058), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n52831), .O(n60065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_7 (.CI(n52831), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n52832));
    SB_LUT4 i7_4_lut_adj_1230 (.I0(\data_in_frame[8] [3]), .I1(n60432), 
            .I2(\data_in_frame[9] [6]), .I3(n60796), .O(n19_adj_5487));
    defparam i7_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1231 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[8] [0]), .I3(n60191), .O(n21_adj_5488));
    defparam i9_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 add_1194_6_lut (.I0(n60058), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n52830), .O(n60061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_6 (.CI(n52830), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n52831));
    SB_LUT4 add_1194_5_lut (.I0(n60058), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n52829), .O(n60062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_5 (.CI(n52829), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n52830));
    SB_LUT4 i11_3_lut_adj_1232 (.I0(n21_adj_5488), .I1(n19_adj_5487), .I2(n20_adj_5486), 
            .I3(GND_net), .O(n60368));
    defparam i11_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 add_1194_4_lut (.I0(n60058), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n52828), .O(n60063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_4 (.CI(n52828), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n52829));
    SB_LUT4 add_1194_3_lut (.I0(n60058), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n52827), .O(n60064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_3 (.CI(n52827), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n52828));
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\data_in_frame[12] [5]), .I1(n28392), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5467));
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 add_1194_2_lut (.I0(n60058), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n60059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n52827));
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5489), .S(n60016));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5490), .S(n60015));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5491), .S(n60014));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5492), .S(n60013));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5493), .S(n60012));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5494), .S(n60011));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5495), .S(n60010));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5496), .S(n60009));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5497), .S(n60008));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8][1] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5498), .S(n60007));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8][2] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5499), .S(n60006));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8][3] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5500), .S(n60005));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8][4] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5501), .S(n60004));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8][5] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5502), .S(n60003));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8][6] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5503), .S(n60002));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8][7] ), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5504), .S(n60001));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5505), .S(n60000));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5506), .S(n59999));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5507), .S(n59998));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5508), .S(n59997));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5509), .S(n59996));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5510), .S(n59995));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5511), .S(n59994));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5512), .S(n59993));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5513), .S(n59992));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5514), .S(n59991));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5515), .S(n59990));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5516), .S(n59989));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5517), .S(n59988));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5518), .S(n59987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5519), .S(n59986));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5520), .S(n59985));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5521), .S(n59984));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5522), .S(n59983));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5523), .S(n59982));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5524), .S(n59981));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5525), .S(n59980));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5526), .S(n59979));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5527), .S(n59978));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5528), .S(n59977));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5529), .S(n59976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5530), .S(n59975));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5531), .S(n59974));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5532), .S(n59973));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5533), .S(n59972));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5534), .S(n60051));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5535), .S(n59971));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5536), .S(n59970));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5537), .S(n59935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5538), .S(n59969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5539), .S(n59968));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5540), .S(n59967));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5541), .S(n59966));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5542), .S(n59965));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5543), .S(n59964));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5544), .S(n59963));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5545), .S(n59962));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5546), .S(n59961));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5547), .S(n59960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5548), .S(n59959));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5549), .S(n59958));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5550), .S(n59957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5551), .S(n59956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5552), .S(n59955));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5553), .S(n59954));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5554), .S(n59953));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5555), .S(n59952));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5556), .S(n59951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5557), .S(n59950));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5558), .S(n59949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5559), .S(n59948));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n31852));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n31851));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n31850));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n31849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5560), .S(n59947));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n31848));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n31847));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n31846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5561), .S(n59946));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n31845));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n31844));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n31843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5562), .S(n59874));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n31842));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n31841));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n31840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5563), .S(n59945));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n31839));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n31838));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n31837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5564), .S(n59944));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n31836));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n31835));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n31834));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5565), .S(n59943));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n31833));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n31832));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n31831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5566), .S(n59942));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n31830));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n31829));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n31828));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n31827));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n31826));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n31825));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5567), .S(n59941));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n31824));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n31823));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n31822));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5568), .S(n59940));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n31818));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5569), .S(n59939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5570), .S(n59938));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14348_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n32539));   // verilog/coms.v(148[4] 304[11])
    defparam i14348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5571), .S(n59937));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5572), .S(n59930));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1234 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60549));
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1235 (.I0(n55176), .I1(n60787), .I2(n60549), 
            .I3(Kp_23__N_993), .O(n55895));
    defparam i3_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14349_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n32540));   // verilog/coms.v(148[4] 304[11])
    defparam i14349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14350_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n32541));   // verilog/coms.v(148[4] 304[11])
    defparam i14350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14351_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n32542));   // verilog/coms.v(148[4] 304[11])
    defparam i14351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1236 (.I0(n62101), .I1(n55895), .I2(\data_in_frame[13] [7]), 
            .I3(GND_net), .O(n60718));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1237 (.I0(n60718), .I1(\data_in_frame[16] [1]), 
            .I2(n60361), .I3(GND_net), .O(n60630));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1237.LUT_INIT = 16'h9696;
    SB_LUT4 i14352_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n32543));   // verilog/coms.v(148[4] 304[11])
    defparam i14352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1238 (.I0(\data_in_frame[14] [1]), .I1(n60368), 
            .I2(\data_in_frame[13] [7]), .I3(n29250), .O(n13_adj_5573));
    defparam i5_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 select_1745_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \FRAME_MATCHER.i_2043__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n30308), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i7_4_lut_adj_1239 (.I0(n13_adj_5573), .I1(n11_adj_5574), .I2(n60488), 
            .I3(n28122), .O(n62398));
    defparam i7_4_lut_adj_1239.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(n60721), .I1(n60827), .I2(GND_net), 
            .I3(GND_net), .O(n55809));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i14353_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n32544));   // verilog/coms.v(148[4] 304[11])
    defparam i14353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48482_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67573));   // verilog/coms.v(158[12:15])
    defparam i48482_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(GND_net), .I3(GND_net), .O(n60477));
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1242 (.I0(n29078), .I1(n60697), .I2(n60477), 
            .I3(n28299), .O(n61964));
    defparam i1_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1243 (.I0(n29250), .I1(n60271), .I2(n64121), 
            .I3(n60670), .O(n60697));
    defparam i1_4_lut_adj_1243.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1244 (.I0(n60697), .I1(n61964), .I2(n60311), 
            .I3(n64095), .O(n55300));
    defparam i1_4_lut_adj_1244.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28067));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(n28812), .I1(n28337), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5575));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(n28332), .I1(\data_in_frame[11] [6]), 
            .I2(n28067), .I3(n6_adj_5575), .O(n28809));
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5576), .S(n59929));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14354_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n32545));   // verilog/coms.v(148[4] 304[11])
    defparam i14354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[12] [5]), .I1(n28224), 
            .I2(GND_net), .I3(GND_net), .O(n60535));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_LUT4 i14355_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n32546));   // verilog/coms.v(148[4] 304[11])
    defparam i14355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1249 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n60882));
    defparam i2_3_lut_adj_1249.LUT_INIT = 16'h9696;
    SB_LUT4 i14356_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n32547));   // verilog/coms.v(148[4] 304[11])
    defparam i14356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1250 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n60238));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1085));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48396_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67571));   // verilog/coms.v(158[12:15])
    defparam i48396_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(n60773), .I1(n28812), .I2(GND_net), 
            .I3(GND_net), .O(n29078));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h9999;
    SB_LUT4 i14357_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [6]), 
            .I3(deadband[22]), .O(n32548));   // verilog/coms.v(148[4] 304[11])
    defparam i14357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[1] [5]), .I1(n60184), 
            .I2(GND_net), .I3(GND_net), .O(n28228));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1253 (.I0(\data_in_frame[8] [0]), .I1(n60203), 
            .I2(n29044), .I3(n28742), .O(n28249));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[8] [1]), .I1(n28249), 
            .I2(GND_net), .I3(GND_net), .O(n60670));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1255 (.I0(n55607), .I1(n60377), .I2(\data_in_frame[10] [2]), 
            .I3(n60848), .O(n10_adj_5577));
    defparam i4_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i14358_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n32549));   // verilog/coms.v(148[4] 304[11])
    defparam i14358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48467_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67568));   // verilog/coms.v(158[12:15])
    defparam i48467_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14359_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n32550));   // verilog/coms.v(148[4] 304[11])
    defparam i14359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1256 (.I0(n60314), .I1(n60473), .I2(\data_in_frame[10] [3]), 
            .I3(n60203), .O(n12_adj_5578));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51998 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [5]), .I2(\data_out_frame[7] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71535));
    defparam byte_transmit_counter_0__bdd_4_lut_51998.LUT_INIT = 16'he4aa;
    SB_LUT4 i48430_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67564));   // verilog/coms.v(158[12:15])
    defparam i48430_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1257 (.I0(\data_in_frame[6] [1]), .I1(n12_adj_5578), 
            .I2(n60767), .I3(\data_in_frame[4] [0]), .O(n28836));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[10] [0]), .I1(n60561), 
            .I2(GND_net), .I3(GND_net), .O(n55074));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1259 (.I0(\data_in_frame[12] [6]), .I1(n28213), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n60494));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2887), .D(n1_adj_5579), .S(n60059));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1260 (.I0(n28836), .I1(n54800), .I2(GND_net), 
            .I3(GND_net), .O(n55777));
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1261 (.I0(\data_in_frame[10] [7]), .I1(n29078), 
            .I2(\data_in_frame[11] [1]), .I3(Kp_23__N_974), .O(n60311));
    defparam i3_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(n28342), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60411));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i14360_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n32551));   // verilog/coms.v(148[4] 304[11])
    defparam i14360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14361_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n32552));   // verilog/coms.v(148[4] 304[11])
    defparam i14361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14_4_lut_adj_1263 (.I0(n60238), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[10] [6]), .I3(n60882), .O(n36));
    defparam i14_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1264 (.I0(n60311), .I1(n55777), .I2(n60807), 
            .I3(n60494), .O(n34_adj_5580));
    defparam i12_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1265 (.I0(n60488), .I1(n36), .I2(n26_adj_5581), 
            .I3(\data_in_frame[12] [0]), .O(n40));
    defparam i18_4_lut_adj_1265.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut (.I0(n60262), .I1(\data_in_frame[10] [4]), .I2(\data_in_frame[3][5] ), 
            .I3(\data_in_frame[8] [1]), .O(n38));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n71535_bdd_4_lut (.I0(n71535), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[4] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71538));
    defparam n71535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14362_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n32553));   // verilog/coms.v(148[4] 304[11])
    defparam i14362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48420_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67563));   // verilog/coms.v(158[12:15])
    defparam i48420_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48381_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67557));   // verilog/coms.v(158[12:15])
    defparam i48381_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i17_3_lut (.I0(\data_in_frame[11] [4]), .I1(n34_adj_5580), .I2(\data_in_frame[12] [1]), 
            .I3(GND_net), .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1266 (.I0(n60787), .I1(n60473), .I2(n60535), 
            .I3(n60377), .O(n37));
    defparam i15_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n55793));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14363_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n32554));   // verilog/coms.v(148[4] 304[11])
    defparam i14363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[13] [2]), .I1(n55793), 
            .I2(GND_net), .I3(GND_net), .O(n60921));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(n55300), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60602));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1269 (.I0(n60888), .I1(n28809), .I2(n62101), 
            .I3(n60759), .O(n10_adj_5582));
    defparam i4_4_lut_adj_1269.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1270 (.I0(\data_in_frame[13] [6]), .I1(n60602), 
            .I2(n10_adj_5582), .I3(n60921), .O(n6_adj_5583));
    defparam i1_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1271 (.I0(n28809), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[15] [5]), .I3(n6_adj_5583), .O(n27478));
    defparam i4_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1272 (.I0(\data_in_frame[9] [3]), .I1(n29193), 
            .I2(\data_in_frame[9] [4]), .I3(n60462), .O(n10_adj_5584));
    defparam i4_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(\data_in_frame[16] [2]), .I1(n60759), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5585));
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1274 (.I0(n55809), .I1(n62398), .I2(n60630), 
            .I3(n6_adj_5585), .O(n55319));
    defparam i4_4_lut_adj_1274.LUT_INIT = 16'h9669;
    SB_LUT4 i14364_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n32555));   // verilog/coms.v(148[4] 304[11])
    defparam i14364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5586), .S(n59928));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1275 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[20] [4]), 
            .I2(n27478), .I3(\data_in_frame[20] [3]), .O(n54931));
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1276 (.I0(\data_in_frame[22] [1]), .I1(n60679), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5587));
    defparam i2_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1277 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[21][7] ), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n7_adj_5588));
    defparam i1_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1278 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[18] [2]), 
            .I2(n60339), .I3(GND_net), .O(n8_adj_5589));
    defparam i3_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 i44969_4_lut (.I0(n26207), .I1(n32_adj_5590), .I2(n8_adj_5589), 
            .I3(\data_in_frame[22] [4]), .O(n64455));
    defparam i44969_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i3_4_lut_adj_1279 (.I0(\data_in_frame[20] [4]), .I1(n60147), 
            .I2(n54794), .I3(\data_in_frame[22] [6]), .O(n62756));
    defparam i3_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1280 (.I0(n29167), .I1(n7_adj_5588), .I2(\data_in_frame[19] [5]), 
            .I3(n8_adj_5587), .O(n61937));
    defparam i5_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1281 (.I0(n60621), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[21][7] ), .I3(GND_net), .O(n6_adj_5591));
    defparam i2_3_lut_adj_1281.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1282 (.I0(n61937), .I1(n62141), .I2(n62756), 
            .I3(n64455), .O(n64195));
    defparam i1_4_lut_adj_1282.LUT_INIT = 16'h0040;
    SB_LUT4 i5_4_lut_adj_1283 (.I0(\data_in_frame[22] [2]), .I1(n60280), 
            .I2(\data_in_frame[19] [6]), .I3(n62188), .O(n12_adj_5592));
    defparam i5_4_lut_adj_1283.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1284 (.I0(\data_in_frame[22]_c [0]), .I1(n64195), 
            .I2(n6_adj_5591), .I3(n62616), .O(n64197));
    defparam i1_4_lut_adj_1284.LUT_INIT = 16'h4884;
    SB_LUT4 i3_4_lut_adj_1285 (.I0(\data_in_frame[23] [7]), .I1(n60851), 
            .I2(n60688), .I3(\data_in_frame[21] [6]), .O(n62426));
    defparam i3_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1286 (.I0(\data_in_frame[21][4] ), .I1(n26256), 
            .I2(n54912), .I3(\data_in_frame[23] [5]), .O(n62467));
    defparam i3_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(n60339), .I1(\data_in_frame[22][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5593));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i14365_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n32556));   // verilog/coms.v(148[4] 304[11])
    defparam i14365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48374_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67556));   // verilog/coms.v(158[12:15])
    defparam i48374_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_1288 (.I0(n26256), .I1(\data_in_frame[21][4] ), 
            .I2(\data_in_frame[23] [6]), .I3(n60851), .O(n62881));
    defparam i2_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1289 (.I0(n62732), .I1(n62467), .I2(n62426), 
            .I3(n64197), .O(n64203));
    defparam i1_4_lut_adj_1289.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut_adj_1290 (.I0(n27478), .I1(n12_adj_5592), .I2(n60679), 
            .I3(\data_in_frame[20] [0]), .O(n61933));
    defparam i6_4_lut_adj_1290.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1291 (.I0(n60280), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[18][1] ), .I3(n4_adj_5593), .O(n62114));
    defparam i2_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1292 (.I0(\data_in_frame[21][1] ), .I1(n55757), 
            .I2(\data_in_frame[21][2] ), .I3(GND_net), .O(n6_adj_5594));
    defparam i2_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1293 (.I0(n62114), .I1(n61933), .I2(n64203), 
            .I3(n62881), .O(n64209));
    defparam i1_4_lut_adj_1293.LUT_INIT = 16'h0080;
    SB_LUT4 i2_3_lut_adj_1294 (.I0(\data_in_frame[21][1] ), .I1(\data_in_frame[23] [2]), 
            .I2(n54882), .I3(GND_net), .O(n62116));
    defparam i2_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1295 (.I0(\data_in_frame[23] [3]), .I1(n64209), 
            .I2(n6_adj_5594), .I3(n55952), .O(n64211));
    defparam i1_4_lut_adj_1295.LUT_INIT = 16'h8448;
    SB_LUT4 i6_4_lut_adj_1296 (.I0(n60805), .I1(\data_in_frame[20] [6]), 
            .I2(n60394), .I3(n54882), .O(n14_adj_5595));
    defparam i6_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1297 (.I0(n62116), .I1(\data_in_frame[23] [0]), 
            .I2(n54882), .I3(n60805), .O(n64213));
    defparam i1_4_lut_adj_1297.LUT_INIT = 16'h2882;
    SB_LUT4 i5_4_lut_adj_1298 (.I0(\data_in_frame[22][7] ), .I1(n60802), 
            .I2(n28517), .I3(\data_in_frame[20] [5]), .O(n13_adj_5596));
    defparam i5_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1299 (.I0(n13_adj_5596), .I1(n64213), .I2(n14_adj_5595), 
            .I3(n64211), .O(n64217));
    defparam i1_4_lut_adj_1299.LUT_INIT = 16'h8400;
    SB_LUT4 i1_4_lut_adj_1300 (.I0(n64217), .I1(n60805), .I2(n55757), 
            .I3(\data_in_frame[23] [1]), .O(n41));
    defparam i1_4_lut_adj_1300.LUT_INIT = 16'h2882;
    SB_LUT4 i14366_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n32557));   // verilog/coms.v(148[4] 304[11])
    defparam i14366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14367_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n32558));   // verilog/coms.v(148[4] 304[11])
    defparam i14367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14368_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n32559));   // verilog/coms.v(148[4] 304[11])
    defparam i14368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[3]_c [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29044));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1302 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[5] [5]), 
            .I2(n28702), .I3(n28266), .O(n60184));
    defparam i3_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1303 (.I0(\data_in_frame[8] [2]), .I1(Kp_23__N_715), 
            .I2(\data_in_frame[6] [1]), .I3(n28761), .O(n4_adj_5597));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_in_frame[8] [3]), .I1(n60538), 
            .I2(GND_net), .I3(GND_net), .O(n28782));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 i48376_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67555));   // verilog/coms.v(158[12:15])
    defparam i48376_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14369_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n32560));   // verilog/coms.v(148[4] 304[11])
    defparam i14369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1305 (.I0(n60184), .I1(n60488), .I2(GND_net), 
            .I3(GND_net), .O(n55607));
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1306 (.I0(\data_in_frame[8] [5]), .I1(n60308), 
            .I2(Kp_23__N_875), .I3(GND_net), .O(n28213));   // verilog/coms.v(239[9:81])
    defparam i2_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1307 (.I0(\data_in_frame[6] [7]), .I1(n29010), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[5] [0]), .O(n60221));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_in_frame[3]_c [1]), .I1(\data_in_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60323));
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i48375_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67554));   // verilog/coms.v(158[12:15])
    defparam i48375_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1309 (.I0(\data_in_frame[2] [6]), .I1(n60221), 
            .I2(n54762), .I3(GND_net), .O(n55176));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1309.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(n28702), .I1(n60323), .I2(GND_net), 
            .I3(GND_net), .O(n60324));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1311 (.I0(n28555), .I1(\data_in_frame[5] [4]), 
            .I2(n60324), .I3(\data_in_frame[7] [5]), .O(n28342));
    defparam i2_4_lut_adj_1311.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_in_frame[7] [1]), .I1(n55176), 
            .I2(GND_net), .I3(GND_net), .O(n55742));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1313 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n37239));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\data_in_frame[3]_c [2]), .I1(n60753), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5598));
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(n37239), .I1(\data_in_frame[5] [2]), 
            .I2(n60459), .I3(n6_adj_5598), .O(n28337));
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60432));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(\data_in_frame[7] [3]), .I1(n28555), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[2] [6]), .O(n60649));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1318 (.I0(n60227), .I1(n60649), .I2(n29010), 
            .I3(GND_net), .O(n29193));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1318.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1319 (.I0(\data_in_frame[2] [4]), .I1(n60456), 
            .I2(\data_in_frame[7] [2]), .I3(\data_in_frame[5] [1]), .O(n12_adj_5599));
    defparam i5_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1320 (.I0(Kp_23__N_758), .I1(n12_adj_5599), .I2(n60700), 
            .I3(n28947), .O(n28812));
    defparam i6_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i48427_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n67553));   // verilog/coms.v(158[12:15])
    defparam i48427_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1321 (.I0(\data_in_frame[6] [2]), .I1(n60432), 
            .I2(Kp_23__N_869), .I3(Kp_23__N_872), .O(n28299));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1322 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5600));
    defparam i2_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_in_frame[3]_c [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60845));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\data_in_frame[3][5] ), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28742));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1325 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(n28690), .I3(GND_net), .O(n60491));
    defparam i2_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1326 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n28157));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60381));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1328 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(n60332), .I3(n60381), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1329 (.I0(Kp_23__N_772), .I1(n60326), .I2(n28715), 
            .I3(\data_in_frame[2]_c [0]), .O(Kp_23__N_875));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60305));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1331 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[1] [4]), .O(n12_adj_5601));   // verilog/coms.v(99[12:25])
    defparam i5_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1332 (.I0(\data_in_frame[3]_c [6]), .I1(n12_adj_5601), 
            .I2(n60305), .I3(\data_in_frame[1] [7]), .O(Kp_23__N_869));   // verilog/coms.v(99[12:25])
    defparam i6_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1333 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60658));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1333.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1334 (.I0(n28742), .I1(n60845), .I2(n60658), 
            .I3(n60241), .O(Kp_23__N_715));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i14370_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n32561));   // verilog/coms.v(148[4] 304[11])
    defparam i14370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(Kp_23__N_875), .I1(Kp_23__N_878), .I2(GND_net), 
            .I3(GND_net), .O(n60224));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 i14371_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n32562));   // verilog/coms.v(148[4] 304[11])
    defparam i14371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12426_1_lut (.I0(n3489), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30616));   // verilog/coms.v(148[4] 304[11])
    defparam i12426_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14372_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n32563));   // verilog/coms.v(148[4] 304[11])
    defparam i14372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1336 (.I0(n28157), .I1(n60772), .I2(n60491), 
            .I3(\data_in_frame[6][6] ), .O(n60773));
    defparam i3_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i14373_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n32564));   // verilog/coms.v(148[4] 304[11])
    defparam i14373_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60796));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h6666;
    SB_LUT4 i14374_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n32565));   // verilog/coms.v(148[4] 304[11])
    defparam i14374_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1338 (.I0(\data_in_frame[0] [0]), .I1(n60796), 
            .I2(n60640), .I3(n60197), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5602), .S(n59927));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48612_4_lut (.I0(\data_out_frame[12] [2]), .I1(byte_transmit_counter[4]), 
            .I2(\data_out_frame[13] [2]), .I3(byte_transmit_counter[0]), 
            .O(n67624));
    defparam i48612_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(n62503), .I1(n60217), .I2(GND_net), 
            .I3(GND_net), .O(n60891));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1340 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5603), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n29303));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1340.LUT_INIT = 16'haaa8;
    SB_LUT4 select_787_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48563_4_lut (.I0(\data_out_frame[14] [2]), .I1(byte_transmit_counter[4]), 
            .I2(\data_out_frame[15] [2]), .I3(byte_transmit_counter[0]), 
            .O(n67738));
    defparam i48563_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i14375_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n32566));   // verilog/coms.v(148[4] 304[11])
    defparam i14375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[3]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60473));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\data_in_frame[6][6] ), .I1(\data_in_frame[6]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60821));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1343 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n28715));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n59203));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i41676_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(n39602), .O(n61124));   // verilog/coms.v(157[7:23])
    defparam i41676_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i[0] ), .O(n76));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i14376_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n32567));   // verilog/coms.v(148[4] 304[11])
    defparam i14376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14377_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n32568));   // verilog/coms.v(148[4] 304[11])
    defparam i14377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14378_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n32569));   // verilog/coms.v(148[4] 304[11])
    defparam i14378_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(n28690), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60332));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_LUT4 equal_309_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_c));   // verilog/coms.v(157[7:23])
    defparam equal_309_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n59201));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n59197));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n59193));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n31683));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n31686));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n32222));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n59189));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17]_c [0]), .C(clk16MHz), 
           .D(n59223));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17]_c [1]), .C(clk16MHz), 
           .D(n59247));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17]_c [2]), .C(clk16MHz), 
           .D(n59251));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17]_c [3]), .C(clk16MHz), 
           .D(n59237));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17]_c [4]), .C(clk16MHz), 
           .D(n59233));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n59315));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17][6] ), .C(clk16MHz), 
           .D(n32704));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n59313));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n32259));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n32262));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n59105));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18][0] ), .C(clk16MHz), 
           .D(n59185));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18][1] ), .C(clk16MHz), 
           .D(n59181));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n59177));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18][3] ), .C(clk16MHz), 
           .D(n32290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n32690));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n32687));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n32684));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n32681));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n32678));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n32293));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18]_c [4]), .C(clk16MHz), 
           .D(n59161));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18][5] ), .C(clk16MHz), 
           .D(n32300));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n59173));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18][7] ), .C(clk16MHz), 
           .D(n32306));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n32310));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n32313));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n59117));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n32320));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n32323));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n32326));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n32329));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n32332));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n32335));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n32338));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n32341));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n32344));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n32347));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1]_c [0]), .C(clk16MHz), 
           .D(n31709));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n32350));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n32353));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1]_c [1]), .C(clk16MHz), 
           .D(n31712));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n59243));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21][0] ), .C(clk16MHz), 
           .D(n32632));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21][1] ), .C(clk16MHz), 
           .D(n32363));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21][2] ), .C(clk16MHz), 
           .D(n59263));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21][3] ), .C(clk16MHz), 
           .D(n59265));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21][4] ), .C(clk16MHz), 
           .D(n59255));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21][5] ), .C(clk16MHz), 
           .D(n59309));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n59297));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21][7] ), .C(clk16MHz), 
           .D(n59305));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22]_c [0]), .C(clk16MHz), 
           .D(n32624));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n32387));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n32390));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22][3] ), .C(clk16MHz), 
           .D(n32393));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n32396));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22][5] ), .C(clk16MHz), 
           .D(n32403));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n32406));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22][7] ), .C(clk16MHz), 
           .D(n32409));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n32413));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n32416));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1]_c [2]), .C(clk16MHz), 
           .D(n59395));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1]_c [3]), .C(clk16MHz), 
           .D(n31718));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n31721));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n32491));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n59159));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n31724));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
           .D(n31727));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n31730));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2]_c [0]), .C(clk16MHz), 
           .D(n24_adj_5604));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
           .D(n31736));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
           .D(n31739));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n32569), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n32568), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n32567), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n32566), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n32565), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n32564), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n32563), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n32562), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n32561), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n32560), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n32559), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n32558), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n32557), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n32556), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n32555), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n32554), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n32553), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n32552), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n32551), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n32550), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n32549), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n32548), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n32547), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n32546), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n32545), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n32544), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n32543), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n32542), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n32541), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n32540), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n32539), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n32538), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n32537), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n32536), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n32535), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n32534), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n32533), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n32532), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n32531), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n32530), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n32529), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n32528), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n32527), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n32526), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n32525), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n32524), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n32523), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n32522), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n32521), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n32520), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n32519), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n32518), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n32517), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n32516), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n32515), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n32514), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n32513), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n32512), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n32511), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n32510), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n32509), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n32508), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n32507), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n32506), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n32505), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n32504), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n32503), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n32502), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n32501), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n32500), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n32499), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n32498), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n32497), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n32496), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n32495), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n32494), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
           .D(n31742));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n32489));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n32488));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n32487));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n32486));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n32485));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n32484));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n32483));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n32482));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n32481));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n32480));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n32479));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n32478));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n32477));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n32476));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n32475));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n32474));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n32473));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n32472));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n32471));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n32470));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n32469));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n32468));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n32467));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(\control_mode[1] ), .C(clk16MHz), .D(n32466));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode_c[2]), .C(clk16MHz), .D(n32465));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
           .D(n31745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode_c[3]), .C(clk16MHz), .D(n32463));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n32462));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n32461));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk16MHz), .D(n32460));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(\control_mode[7] ), .C(clk16MHz), .D(n32459));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n32458));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n32457));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n37917));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n32455));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1345 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n39602), .I3(\FRAME_MATCHER.i[0] ), .O(n30619));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1345.LUT_INIT = 16'hbfff;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2887), .D(n2_adj_5605), .S(n59926));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n32454));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n32453));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n32452));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n32451));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n32450));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n32449));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n32448));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n32447));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n32446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n32445));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n32444));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n32443), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n32442), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n32441), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n32440), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n32439), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n32438), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n32437), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n32436), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n32435), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n32434), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n32433), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n32432), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n32431), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n32430), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n32429), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n32428), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n32427), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n32426), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n32425), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n32424), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n32423), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n32422), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n32421), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
           .D(n31748));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
           .D(n31751));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n31754));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_0__3__I_0_2_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_758));   // verilog/coms.v(77[16:27])
    defparam data_in_frame_0__3__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n31757));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19524_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [1]), 
            .I3(\data_in_frame[19] [1]), .O(n4945[1]));   // verilog/coms.v(148[4] 304[11])
    defparam i19524_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3]_c [1]), .C(clk16MHz), 
           .D(n59453));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i17641_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [2]), 
            .I3(\data_in_frame[19] [2]), .O(n4945[2]));   // verilog/coms.v(148[4] 304[11])
    defparam i17641_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i48723_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n79), .I3(\FRAME_MATCHER.i[0] ), .O(n67702));   // verilog/coms.v(157[7:23])
    defparam i48723_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_4_lut_adj_1346 (.I0(n60259), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [7]), .I3(n4_adj_5606), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i2_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n31703));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1347 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n60130), .I3(\FRAME_MATCHER.i[0] ), .O(n60134));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1347.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n59771), .I3(\FRAME_MATCHER.i[0] ), .O(n59777));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1348.LUT_INIT = 16'hfbff;
    SB_LUT4 i13983_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n32174));
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3]_c [2]), .C(clk16MHz), 
           .D(n59415));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13986_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n32177));
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFR \FRAME_MATCHER.i_2043__i1  (.Q(\FRAME_MATCHER.i[1] ), .C(clk16MHz), 
            .D(n30347), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i2  (.Q(\FRAME_MATCHER.i[2] ), .C(clk16MHz), 
            .D(n30349), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk16MHz), 
            .D(n30351), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n30353), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk16MHz), 
            .D(n30355), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n30357), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n30359), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n30361), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n30363), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n30365), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n30367), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n30369), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n30371), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n30373), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n30375), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n30377), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n30379), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n30381), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n30383), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n30385), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n30387), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n30389), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n30391), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n30393), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n30395), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n30397), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n30399), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n30401), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n30403), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n30405), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n30407), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_2_lut_adj_1349 (.I0(\data_in_frame[1]_c [0]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n60248));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1349.LUT_INIT = 16'h6666;
    SB_LUT4 i13989_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n32180));
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n31766));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n31696), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3]_c [4]), .C(clk16MHz), 
           .D(n59457));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3][5] ), .C(clk16MHz), 
           .D(n31772));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13992_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n32183));
    defparam i13992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n31695));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(\control_mode[0] ), .C(clk16MHz), .D(n31694));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n31693));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n31692), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n31691), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n31690), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n31689), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3]_c [6]), .C(clk16MHz), 
           .D(n31775));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3]_c [7]), .C(clk16MHz), 
           .D(n31778));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13995_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n32186));
    defparam i13995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_772));   // verilog/coms.v(81[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13998_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n32189));
    defparam i13998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14001_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n32192));
    defparam i14001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n59465));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i4_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3][3] ), 
            .I3(\data_in_frame[19] [3]), .O(n4945[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n31784));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i19437_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [4]), 
            .I3(\data_in_frame[19] [4]), .O(n4945[4]));   // verilog/coms.v(148[4] 304[11])
    defparam i19437_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i14004_3_lut_4_lut (.I0(n41173), .I1(n59771), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n32195));
    defparam i14004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n31787));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i6_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3][5] ), 
            .I3(\data_in_frame[19] [5]), .O(n4945[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i7_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [6]), 
            .I3(\data_in_frame[19] [6]), .O(n4945[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_adj_1350 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60259));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1350.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1351 (.I0(\data_in_frame[0] [5]), .I1(Kp_23__N_767), 
            .I2(\data_in_frame[1]_c [0]), .I3(GND_net), .O(n26984));   // verilog/coms.v(80[16:27])
    defparam i1_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1352 (.I0(n29010), .I1(n26984), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[2] [7]), .O(n60700));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1353 (.I0(\data_in_frame[5] [4]), .I1(n60528), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n28106));
    defparam i2_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1354 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3]_c [1]), 
            .I2(\data_in_frame[5] [1]), .I3(GND_net), .O(n60227));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60456));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60640));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60326));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60767));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1359 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[3]_c [6]), .I3(\data_in_frame[3][3] ), .O(n64245));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1360 (.I0(n64245), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[3][5] ), .I3(\data_in_frame[3]_c [4]), .O(n64247));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1361 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[2]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n64253));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1362 (.I0(n60767), .I1(n60326), .I2(n60640), 
            .I3(n60456), .O(n64257));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1363 (.I0(n60227), .I1(n64257), .I2(n64253), 
            .I3(n64247), .O(n64261));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1364 (.I0(n60332), .I1(n54798), .I2(n60459), 
            .I3(n64261), .O(n64269));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1365 (.I0(n28106), .I1(n60700), .I2(n64269), 
            .I3(n64267), .O(n62503));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1366 (.I0(n54762), .I1(n62503), .I2(n60609), 
            .I3(n64085), .O(n60488));
    defparam i1_4_lut_adj_1366.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60241));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_adj_1368 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(ID[2]), .I3(ID[1]), .O(n6_adj_5607));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1368.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1369 (.I0(ID[7]), .I1(\data_in_frame[0] [3]), .I2(\data_in_frame[0] [7]), 
            .I3(ID[3]), .O(n6_adj_5608));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1369.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1370 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [4]), 
            .I2(ID[0]), .I3(ID[4]), .O(n5_adj_5609));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1370.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1371 (.I0(ID[6]), .I1(\data_in_frame[0] [5]), .I2(\data_in_frame[0] [6]), 
            .I3(ID[5]), .O(n5_adj_5610));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1371.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1372 (.I0(n5_adj_5610), .I1(n5_adj_5609), .I2(n6_adj_5608), 
            .I3(n6_adj_5607), .O(n32_adj_5590));
    defparam i1_4_lut_adj_1372.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1373 (.I0(n60772), .I1(n60308), .I2(\data_in_frame[8] [1]), 
            .I3(n60891), .O(n10_adj_5611));
    defparam i4_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1374 (.I0(n60773), .I1(n60538), .I2(n10_adj_5611), 
            .I3(n60224), .O(n15_adj_5612));
    defparam i2_4_lut_adj_1374.LUT_INIT = 16'h2882;
    SB_LUT4 i1_3_lut_adj_1375 (.I0(n32_adj_5590), .I1(\data_in_frame[8] [0]), 
            .I2(n60271), .I3(GND_net), .O(n14_adj_5613));
    defparam i1_3_lut_adj_1375.LUT_INIT = 16'h1414;
    SB_LUT4 i9_4_lut_adj_1376 (.I0(n28213), .I1(n55607), .I2(n28782), 
            .I3(n4_adj_5597), .O(n22));
    defparam i9_4_lut_adj_1376.LUT_INIT = 16'h0004;
    SB_LUT4 i8_4_lut_adj_1377 (.I0(n15_adj_5612), .I1(Kp_23__N_974), .I2(n7_adj_5600), 
            .I3(\data_in_frame[8] [6]), .O(n21_adj_5614));
    defparam i8_4_lut_adj_1377.LUT_INIT = 16'h0802;
    SB_LUT4 i10_4_lut_adj_1378 (.I0(n28299), .I1(n28812), .I2(n29193), 
            .I3(n14_adj_5613), .O(n23_adj_5615));
    defparam i10_4_lut_adj_1378.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1379 (.I0(n23_adj_5615), .I1(n28337), .I2(n21_adj_5614), 
            .I3(n22), .O(n6_adj_5616));
    defparam i1_4_lut_adj_1379.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut_adj_1380 (.I0(n28357), .I1(n55742), .I2(n28342), 
            .I3(n6_adj_5616), .O(n35072));
    defparam i4_4_lut_adj_1380.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut_adj_1381 (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n35072), .I3(GND_net), .O(n31_adj_5617));   // verilog/TinyFPGA_B.v(4[10:13])
    defparam i1_3_lut_adj_1381.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13133_4_lut (.I0(n2887), .I1(LED_c), .I2(n31_adj_5617), .I3(n60119), 
            .O(n31324));   // verilog/coms.v(130[12] 305[6])
    defparam i13133_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i16893_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n35084));   // verilog/coms.v(118[11:12])
    defparam i16893_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i20023_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[17]_c [4]), .O(n4945[20]));   // verilog/coms.v(148[4] 304[11])
    defparam i20023_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i22_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[17] [5]), .O(n4945[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1382 (.I0(\data_out_frame[17] [3]), .I1(n62343), 
            .I2(GND_net), .I3(GND_net), .O(n60836));
    defparam i1_2_lut_adj_1382.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1383 (.I0(n60744), .I1(\data_out_frame[15] [2]), 
            .I2(n60909), .I3(\data_out_frame[14] [7]), .O(n14_adj_5618));
    defparam i6_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1384 (.I0(\data_out_frame[14] [6]), .I1(n60836), 
            .I2(n60531), .I3(\data_out_frame[17] [2]), .O(n13_adj_5619));
    defparam i5_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1385 (.I0(\data_out_frame[19] [4]), .I1(n13_adj_5619), 
            .I2(n14_adj_5618), .I3(GND_net), .O(n55907));
    defparam i1_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60441));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(n35084), 
            .I3(GND_net), .O(n5_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 mux_1087_i1_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3] [0]), 
            .I3(\data_in_frame[19] [0]), .O(n4945[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_out_frame[15] [0]), .I1(n55744), 
            .I2(GND_net), .I3(GND_net), .O(n60531));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1388 (.I0(n28456), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[12] [4]), 
            .O(n29117));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1389 (.I0(\data_out_frame[18] [6]), .I1(n60739), 
            .I2(GND_net), .I3(GND_net), .O(n60876));
    defparam i1_2_lut_adj_1389.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1390 (.I0(n55748), .I1(n60876), .I2(n60405), 
            .I3(n55783), .O(n55567));
    defparam i3_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i24_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[17] [7]), .O(n4945[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i3_3_lut_adj_1391 (.I0(n29117), .I1(n60452), .I2(n60879), 
            .I3(GND_net), .O(n8_adj_5620));
    defparam i3_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1392 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[16] [6]), 
            .I2(n8_adj_5620), .I3(n60858), .O(n28907));
    defparam i1_4_lut_adj_1392.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1393 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60517));
    defparam i1_2_lut_adj_1393.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1394 (.I0(n60643), .I1(n28968), .I2(\data_out_frame[11] [3]), 
            .I3(n60830), .O(n10_adj_5621));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1395 (.I0(\data_out_frame[14] [0]), .I1(n60388), 
            .I2(n28427), .I3(\data_out_frame[11] [6]), .O(n29047));
    defparam i3_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1396 (.I0(\data_out_frame[13] [5]), .I1(n27445), 
            .I2(GND_net), .I3(GND_net), .O(n29148));
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_c));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1397 (.I0(\data_out_frame[10] [1]), .I1(n60709), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5622));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1397.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1398 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(n60349), .I3(n6_adj_5622), .O(n1510));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1399 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[12] [7]), 
            .I2(n60861), .I3(n60235), .O(n13_adj_5623));   // verilog/coms.v(77[16:27])
    defparam i5_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1400 (.I0(n13_adj_5623), .I1(n55800), .I2(n12_adj_5624), 
            .I3(\data_out_frame[12] [6]), .O(n55744));   // verilog/coms.v(77[16:27])
    defparam i7_4_lut_adj_1400.LUT_INIT = 16'h9669;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(74[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1401 (.I0(\data_out_frame[9] [4]), .I1(n1312), 
            .I2(GND_net), .I3(GND_net), .O(n60388));
    defparam i1_2_lut_adj_1401.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1402 (.I0(\data_out_frame[11] [7]), .I1(n60736), 
            .I2(n60188), .I3(n28873), .O(n62099));
    defparam i3_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1403 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[7] [4]), .O(n60709));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5481));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48693_2_lut (.I0(\data_out_frame[3][3] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67669));
    defparam i48693_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\data_out_frame[12] [1]), .I1(n62099), 
            .I2(GND_net), .I3(GND_net), .O(n60544));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51978 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[1]), .O(n71343));
    defparam byte_transmit_counter_0__bdd_4_lut_51978.LUT_INIT = 16'he4aa;
    SB_LUT4 n71343_bdd_4_lut (.I0(n71343), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71346));
    defparam n71343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1087_i23_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[17][6] ), .O(n4945[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i4_4_lut_adj_1405 (.I0(n60544), .I1(\data_out_frame[12] [0]), 
            .I2(\data_out_frame[5] [4]), .I3(n60709), .O(n10_adj_5625));
    defparam i4_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1406 (.I0(n60168), .I1(n55852), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n60485));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(\data_out_frame[10] [0]), .I1(n28427), 
            .I2(GND_net), .I3(GND_net), .O(n28873));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60655));
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_223_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n60555), .I3(n60762), .O(n3_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_out_frame[25] [5]), .I1(n60480), 
            .I2(GND_net), .I3(GND_net), .O(n60555));
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1410 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n28968));
    defparam i2_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1411 (.I0(\data_out_frame[5] [1]), .I1(n60317), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n28427));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_adj_1411.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1087_i10_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[18][1] ), .O(n4945[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[8][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n60345));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1087_i11_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [2]), 
            .I3(\data_in_frame[18] [2]), .O(n4945[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[7] [0]), .I3(n29177), .O(n46));   // verilog/coms.v(78[16:27])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1413 (.I0(\data_out_frame[23] [4]), .I1(n54859), 
            .I2(n60818), .I3(GND_net), .O(n8_adj_5626));
    defparam i3_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_222_i3_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5626), .I3(n60555), 
            .O(n3_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_222_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i17_4_lut_adj_1414 (.I0(\data_out_frame[4] [4]), .I1(n60209), 
            .I2(n60712), .I3(\data_out_frame[6] [3]), .O(n44));   // verilog/coms.v(78[16:27])
    defparam i17_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1415 (.I0(\data_out_frame[7] [2]), .I1(n60706), 
            .I2(\data_out_frame[4] [6]), .I3(n60255), .O(n45));   // verilog/coms.v(78[16:27])
    defparam i18_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i12_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [3]), 
            .I3(\data_in_frame[18][3] ), .O(n4945[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i16_4_lut_adj_1416 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[8][5] ), 
            .I2(\data_out_frame[9] [0]), .I3(n60317), .O(n43));   // verilog/coms.v(78[16:27])
    defparam i16_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1417 (.I0(n60397), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[9] [5]), .I3(n1130), .O(n42));   // verilog/coms.v(78[16:27])
    defparam i15_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));   // verilog/coms.v(78[16:27])
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[7] [6]), .I1(n28968), .I2(\data_out_frame[7] [1]), 
            .I3(\data_out_frame[5] [4]), .O(n47));   // verilog/coms.v(78[16:27])
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5430));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_4_lut (.I0(n47), .I1(n52), .I2(n41_adj_5627), .I3(n42), 
            .O(n55852));   // verilog/coms.v(78[16:27])
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i4_3_lut (.I0(\data_out_frame[4] [3]), 
            .I1(\data_out_frame[5] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_adj_5429));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1418 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8][5] ), 
            .I2(n55852), .I3(n28031), .O(n10_adj_5628));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1419 (.I0(\data_out_frame[4] [2]), .I1(n10_adj_5628), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n62234));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i45122_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64617));
    defparam i45122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45123_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64618));
    defparam i45123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45342_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64837));
    defparam i45342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45341_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64836));
    defparam i45341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45113_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64608));
    defparam i45113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45114_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64609));
    defparam i45114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1420 (.I0(n62234), .I1(n28427), .I2(\data_out_frame[10] [0]), 
            .I3(n60345), .O(n60235));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1420.LUT_INIT = 16'h9669;
    SB_LUT4 i45117_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64612));
    defparam i45117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1087_i13_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [4]), 
            .I3(\data_in_frame[18]_c [4]), .O(n4945[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i14_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [5]), 
            .I3(\data_in_frame[18][5] ), .O(n4945[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i15_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[18] [6]), .O(n4945[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_4_lut_adj_1421 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [7]), 
            .I2(\control_mode[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5427));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1421.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1422 (.I0(n55800), .I1(n60867), .I2(GND_net), 
            .I3(GND_net), .O(n60839));
    defparam i1_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 i45116_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64611));
    defparam i45116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45092_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64587));
    defparam i45092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45093_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64588));
    defparam i45093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45096_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64591));
    defparam i45096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45095_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64590));
    defparam i45095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48682_2_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67667));
    defparam i48682_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1423 (.I0(n60839), .I1(n28024), .I2(n60235), 
            .I3(n40_adj_5629), .O(n14_adj_5630));
    defparam i6_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i19925_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2] [7]), 
            .I3(\data_in_frame[18][7] ), .O(n4945[15]));   // verilog/coms.v(148[4] 304[11])
    defparam i19925_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i7_4_lut_adj_1424 (.I0(\data_out_frame[13] [1]), .I1(n14_adj_5630), 
            .I2(n10_adj_5631), .I3(n60168), .O(n62343));
    defparam i7_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1425 (.I0(n60715), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[11] [0]), .I3(n60355), .O(n15_adj_5632));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1426 (.I0(n15_adj_5632), .I1(\data_out_frame[6] [6]), 
            .I2(n14_adj_5633), .I3(\data_out_frame[8][4] ), .O(n28056));   // verilog/coms.v(77[16:43])
    defparam i8_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60643));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 i45404_3_lut (.I0(\data_out_frame[8][1] ), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64899));
    defparam i45404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45405_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64900));
    defparam i45405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45402_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64897));
    defparam i45402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45401_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64896));
    defparam i45401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45101_3_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64596));
    defparam i45101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45102_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64597));
    defparam i45102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45399_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64894));
    defparam i45399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48476_2_lut (.I0(\data_out_frame[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67668));
    defparam i48476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(\data_out_frame[7] [1]), .I1(n28446), 
            .I2(GND_net), .I3(GND_net), .O(n28888));
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h6666;
    SB_LUT4 i45398_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64893));
    defparam i45398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45128_3_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64623));
    defparam i45128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45129_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64624));
    defparam i45129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45354_3_lut (.I0(\data_out_frame[26] [5]), .I1(\data_out_frame[27] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64849));
    defparam i45354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_221_i3_2_lut (.I0(n60286), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_221_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i45353_3_lut (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[25] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64848));
    defparam i45353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48681_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n67742));
    defparam i48681_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i45389_3_lut (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64884));
    defparam i45389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45390_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64885));
    defparam i45390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45372_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64867));
    defparam i45372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45371_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64866));
    defparam i45371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45125_3_lut (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64620));
    defparam i45125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45126_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64621));
    defparam i45126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1429 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28453));
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h6666;
    SB_LUT4 i45366_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64861));
    defparam i45366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45333_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64828));
    defparam i45333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45367_4_lut (.I0(n64861), .I1(n67742), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[0]), .O(n64862));
    defparam i45367_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i45332_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64827));
    defparam i45332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45302_3_lut (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64797));
    defparam i45302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45303_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64798));
    defparam i45303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20062_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1]_c [0]), 
            .I3(\data_in_frame[17]_c [0]), .O(n4945[16]));   // verilog/coms.v(148[4] 304[11])
    defparam i20062_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i45135_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64630));
    defparam i45135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45134_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64629));
    defparam i45134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1430 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[4] [7]), 
            .I2(n60546), .I3(\data_out_frame[6] [7]), .O(n7_adj_5634));
    defparam i2_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i45365_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64860));
    defparam i45365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1431 (.I0(n7_adj_5634), .I1(n28453), .I2(n1312), 
            .I3(n28888), .O(n54796));
    defparam i4_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i45297_3_lut (.I0(n71592), .I1(n71580), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n64792));
    defparam i45297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1432 (.I0(n29177), .I1(\data_out_frame[9] [2]), 
            .I2(n1130), .I3(n60643), .O(n10_adj_5635));
    defparam i4_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_220_i3_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n60567), .I3(n55840), .O(n3_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1433 (.I0(n28745), .I1(n54796), .I2(GND_net), 
            .I3(GND_net), .O(n55769));
    defparam i1_2_lut_adj_1433.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(n28056), .I1(n62343), .I2(GND_net), 
            .I3(GND_net), .O(n55750));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h9999;
    SB_LUT4 i19867_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1]_c [1]), 
            .I3(\data_in_frame[17]_c [1]), .O(n4945[17]));   // verilog/coms.v(148[4] 304[11])
    defparam i19867_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i45298_3_lut (.I0(n64791), .I1(n64792), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n64793));
    defparam i45298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5636));   // verilog/coms.v(88[17:28])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1435 (.I0(\FRAME_MATCHER.state[3] ), .I1(n55840), 
            .I2(n8_adj_5637), .I3(n60558), .O(n3_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1435.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1436 (.I0(n9_adj_5636), .I1(n60335), .I2(n62457), 
            .I3(n28441), .O(n60405));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1436.LUT_INIT = 16'h9669;
    SB_LUT4 i6_3_lut (.I0(n64793), .I1(n71556), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(tx_data[2]));   // verilog/coms.v(105[12:33])
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19864_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1]_c [2]), 
            .I3(\data_in_frame[17]_c [2]), .O(n4945[18]));   // verilog/coms.v(148[4] 304[11])
    defparam i19864_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i4_4_lut_adj_1437 (.I0(\data_out_frame[16] [6]), .I1(n54970), 
            .I2(n60405), .I3(n29259), .O(n10_adj_5638));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1438 (.I0(\data_out_frame[18] [7]), .I1(n55783), 
            .I2(n10_adj_5638), .I3(\data_out_frame[16] [4]), .O(n60739));
    defparam i1_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1439 (.I0(n60842), .I1(n28615), .I2(n55750), 
            .I3(n55769), .O(n40_adj_5639));
    defparam i16_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i20032_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[1]_c [3]), 
            .I3(\data_in_frame[17]_c [3]), .O(n4945[19]));   // verilog/coms.v(148[4] 304[11])
    defparam i20032_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i14_4_lut_adj_1440 (.I0(n55856), .I1(n60655), .I2(\data_out_frame[14] [6]), 
            .I3(\data_out_frame[14] [4]), .O(n38_adj_5640));
    defparam i14_4_lut_adj_1440.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1441 (.I0(\data_out_frame[11] [5]), .I1(n55577), 
            .I2(\data_out_frame[11] [4]), .I3(n55985), .O(n39_adj_5641));
    defparam i15_4_lut_adj_1441.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1442 (.I0(\data_out_frame[10] [5]), .I1(n55744), 
            .I2(n29259), .I3(n60206), .O(n37_adj_5642));
    defparam i13_4_lut_adj_1442.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1443 (.I0(n29148), .I1(n1699), .I2(\data_out_frame[14] [1]), 
            .I3(n54834), .O(n42_adj_5643));
    defparam i18_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n37_adj_5642), .I1(n39_adj_5641), .I2(n38_adj_5640), 
            .I3(n40_adj_5639), .O(n46_adj_5644));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1444 (.I0(n1563), .I1(\data_out_frame[11] [1]), 
            .I2(n28427), .I3(n29017), .O(n41_adj_5645));
    defparam i17_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1445 (.I0(n41_adj_5645), .I1(\data_out_frame[15] [4]), 
            .I2(n46_adj_5644), .I3(n42_adj_5643), .O(n10_adj_5646));
    defparam i1_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51820 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[1]), .O(n71331));
    defparam byte_transmit_counter_0__bdd_4_lut_51820.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1446 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[15] [3]), .I3(n10_adj_5646), .O(n16_adj_5647));
    defparam i7_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1447 (.I0(n60517), .I1(n16_adj_5647), .I2(n12_adj_5648), 
            .I3(n29148), .O(n62457));
    defparam i8_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1448 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n28441));
    defparam i1_2_lut_adj_1448.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_218_i3_4_lut (.I0(n55732), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5649), .I3(n60552), .O(n3_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i4_4_lut_adj_1449 (.I0(n7_adj_5650), .I1(\data_out_frame[19] [1]), 
            .I2(n62457), .I3(n60739), .O(n60879));
    defparam i4_4_lut_adj_1449.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1087_i9_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[2]_c [0]), 
            .I3(\data_in_frame[18][0] ), .O(n4945[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i19385_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(\data_in_frame[3]_c [7]), 
            .I3(\data_in_frame[19] [7]), .O(n4945[7]));   // verilog/coms.v(148[4] 304[11])
    defparam i19385_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i3_4_lut_adj_1450 (.I0(\data_out_frame[23] [1]), .I1(n28961), 
            .I2(\data_out_frame[22] [7]), .I3(n61784), .O(n60824));
    defparam i3_4_lut_adj_1450.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[20] [0]), .I1(n55462), 
            .I2(GND_net), .I3(GND_net), .O(n60903));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1452 (.I0(n60352), .I1(n60520), .I2(n60703), 
            .I3(n60824), .O(n62217));
    defparam i3_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1453 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(n62217), .I3(GND_net), .O(n14_adj_5651));
    defparam i5_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1454 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8][6] ), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n60209));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1455 (.I0(n60903), .I1(n54842), .I2(\data_out_frame[18] [3]), 
            .I3(n55514), .O(n15_adj_5652));
    defparam i6_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1456 (.I0(n15_adj_5652), .I1(n55273), .I2(n14_adj_5651), 
            .I3(n55985), .O(n60567));
    defparam i8_4_lut_adj_1456.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_out_frame[4] [7]), .I1(n60633), 
            .I2(GND_net), .I3(GND_net), .O(n60830));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1458 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n29017));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1458.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60355));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1460 (.I0(\data_out_frame[9] [2]), .I1(n60355), 
            .I2(\data_out_frame[13] [4]), .I3(\data_out_frame[7] [1]), .O(n12_adj_5653));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1461 (.I0(n29017), .I1(n12_adj_5653), .I2(n60830), 
            .I3(n40_adj_5629), .O(n55577));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60188));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1463 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28020));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1463.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1464 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60546));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1464.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1465 (.I0(n28020), .I1(n60188), .I2(n1191), .I3(\data_out_frame[5] [4]), 
            .O(n1168));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1466 (.I0(n60329), .I1(\data_out_frame[23] [0]), 
            .I2(n28483), .I3(GND_net), .O(n14_adj_5654));
    defparam i5_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1467 (.I0(n60627), .I1(n60452), .I2(n60903), 
            .I3(n60912), .O(n15_adj_5655));
    defparam i6_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(n1168), .I1(n60633), .I2(GND_net), 
            .I3(GND_net), .O(n28697));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60268));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i5673_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1964), 
            .I2(n61999), .I3(n4452), .O(n23514));   // verilog/coms.v(148[4] 304[11])
    defparam i5673_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(\data_out_frame[10] [7]), .I1(n28031), 
            .I2(GND_net), .I3(GND_net), .O(n60861));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1471 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8][6] ), 
            .I2(\data_out_frame[8][5] ), .I3(GND_net), .O(n60715));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1472 (.I0(n15_adj_5655), .I1(n60498), .I2(n14_adj_5654), 
            .I3(n60812), .O(n55732));
    defparam i8_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1473 (.I0(n60567), .I1(\data_out_frame[25] [4]), 
            .I2(n60499), .I3(n60818), .O(n60286));
    defparam i3_4_lut_adj_1473.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1474 (.I0(n60715), .I1(n60861), .I2(\data_out_frame[13] [3]), 
            .I3(n60268), .O(n12_adj_5656));   // verilog/coms.v(100[12:26])
    defparam i5_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1475 (.I0(\data_out_frame[11] [2]), .I1(n12_adj_5656), 
            .I2(n60915), .I3(n28697), .O(n28615));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1476 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n28031));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1477 (.I0(n23514), .I1(n1964), .I2(n25071), .I3(n4_adj_5657), 
            .O(n29420));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1477.LUT_INIT = 16'hbbba;
    SB_LUT4 i6_4_lut_adj_1478 (.I0(n60824), .I1(n54742), .I2(n60482), 
            .I3(\data_out_frame[21] [0]), .O(n14_adj_5658));
    defparam i6_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_out_frame[20] [7]), .I1(n55746), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5659));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(\data_in_frame[18][3] ), .I1(n55319), 
            .I2(\data_in_frame[18][5] ), .I3(GND_net), .O(n60802));
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\data_in_frame[18][3] ), .I1(n55319), 
            .I2(n54931), .I3(\data_in_frame[22][5] ), .O(n62141));
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1482 (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[10] [5]), .I3(n1191), .O(n60365));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1483 (.I0(\data_out_frame[8][4] ), .I1(n60867), 
            .I2(n60724), .I3(n60365), .O(n1522));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60349));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60727));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h6666;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2073));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1486 (.I0(n9_adj_5659), .I1(n14_adj_5658), .I2(n55732), 
            .I3(n55838), .O(n55840));
    defparam i7_4_lut_adj_1486.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1487 (.I0(\data_out_frame[24] [7]), .I1(n54792), 
            .I2(n55732), .I3(\data_out_frame[22] [6]), .O(n60558));
    defparam i3_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n60712));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60397));
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1490 (.I0(n60255), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [7]), .I3(n60736), .O(n10_adj_5660));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(n60799), .I1(n60480), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5661));
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1492 (.I0(n60558), .I1(n60570), .I2(n55840), 
            .I3(n60286), .O(n12_adj_5662));
    defparam i5_4_lut_adj_1492.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_217_i3_4_lut (.I0(n55802), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5662), .I3(n8_adj_5661), .O(n3_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i5_3_lut_adj_1493 (.I0(\data_out_frame[10] [2]), .I1(n10_adj_5660), 
            .I2(\data_out_frame[10] [1]), .I3(GND_net), .O(n1513));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1493.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1494 (.I0(n60712), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[4] [0]), .I3(n60727), .O(n10_adj_5663));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60724));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60618));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1497 (.I0(\data_out_frame[8][1] ), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n60255));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1497.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1498 (.I0(n60618), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[8][3] ), .I3(n60724), .O(n10_adj_5664));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1499 (.I0(n60255), .I1(n10_adj_5664), .I2(\data_out_frame[10] [3]), 
            .I3(GND_net), .O(n1519));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_adj_1499.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[12] [6]), .I1(n1522), 
            .I2(GND_net), .I3(GND_net), .O(n60909));
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1501 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(\data_out_frame[14] [7]), .I3(GND_net), .O(n60842));
    defparam i2_3_lut_adj_1501.LUT_INIT = 16'h9696;
    SB_LUT4 i44802_4_lut (.I0(n1964), .I1(n1967), .I2(n3303), .I3(n1970), 
            .O(n64282));   // verilog/coms.v(139[4] 141[7])
    defparam i44802_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60552));
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1503 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n60214));
    defparam i2_3_lut_adj_1503.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1504 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60335));
    defparam i1_2_lut_adj_1504.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1505 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1967), 
            .I2(n64282), .I3(n62119), .O(n58999));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1505.LUT_INIT = 16'hb3a0;
    SB_LUT4 select_787_Select_216_i3_4_lut (.I0(n60552), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60793), .I3(n60283), .O(n3_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_216_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i51425_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[4] [0]), .I2(n30673), 
            .I3(GND_net), .O(n59465));   // verilog/coms.v(94[13:20])
    defparam i51425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13587_3_lut (.I0(\data_in_frame[3]_c [7]), .I1(rx_data[7]), 
            .I2(n30671), .I3(GND_net), .O(n31778));   // verilog/coms.v(130[12] 305[6])
    defparam i13587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1506 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[25] [1]), .I3(\data_out_frame[25] [6]), 
            .O(n60799));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i13584_3_lut (.I0(\data_in_frame[3]_c [6]), .I1(rx_data[6]), 
            .I2(n30671), .I3(GND_net), .O(n31775));   // verilog/coms.v(130[12] 305[6])
    defparam i13584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1507 (.I0(\data_out_frame[25] [3]), .I1(n60799), 
            .I2(\data_out_frame[25] [4]), .I3(GND_net), .O(n60793));
    defparam i2_3_lut_adj_1507.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1508 (.I0(n60214), .I1(n60646), .I2(\data_out_frame[16] [7]), 
            .I3(GND_net), .O(n55179));
    defparam i2_3_lut_adj_1508.LUT_INIT = 16'h9696;
    SB_LUT4 i20061_3_lut (.I0(\control_mode[0] ), .I1(\data_in_frame[1]_c [0]), 
            .I2(n25151), .I3(GND_net), .O(n31694));
    defparam i20061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[15] [4]), .O(n9_adj_5484));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i51424_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[3]_c [4]), 
            .I2(n30671), .I3(GND_net), .O(n59457));   // verilog/coms.v(94[13:20])
    defparam i51424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_adj_1509 (.I0(n54978), .I1(n60570), .I2(n60793), 
            .I3(GND_net), .O(n8_adj_5665));
    defparam i3_3_lut_adj_1509.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_out_frame[17] [2]), .I1(n60452), 
            .I2(GND_net), .I3(GND_net), .O(n28070));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1511 (.I0(\data_out_frame[21] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(n60703), .I3(n6_adj_5666), .O(n54859));
    defparam i4_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[9] [0]), .I3(n60411), .O(n26_adj_5581));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1512 (.I0(\data_out_frame[21] [4]), .I1(n28070), 
            .I2(n60445), .I3(n6_adj_5667), .O(n62192));
    defparam i4_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_215_i3_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5665), .I3(n60685), 
            .O(n3_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(n28907), .I1(n55567), .I2(GND_net), 
            .I3(GND_net), .O(n60498));
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(n62192), .I1(n54859), .I2(GND_net), 
            .I3(GND_net), .O(n60466));
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h9999;
    SB_LUT4 i5678_4_lut (.I0(n1968), .I1(\FRAME_MATCHER.state[3] ), .I2(n1970), 
            .I3(n27855), .O(n23519));   // verilog/coms.v(148[4] 304[11])
    defparam i5678_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(\data_out_frame[21] [5]), .I1(n55907), 
            .I2(GND_net), .I3(GND_net), .O(n60159));
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1516 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n60232));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1516.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(n60764), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5668));
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1518 (.I0(n60159), .I1(n60466), .I2(\data_out_frame[25] [6]), 
            .I3(n60499), .O(n12_adj_5669));
    defparam i5_4_lut_adj_1518.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_208_i3_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n12_adj_5669), .I3(n8_adj_5668), 
            .O(n3_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_208_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_787_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1519 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n60787));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1519.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1520 (.I0(\data_in_frame[10] [5]), .I1(n28782), 
            .I2(n28213), .I3(\data_in_frame[12] [7]), .O(n60885));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1521 (.I0(rx_data[2]), .I1(\data_in_frame[3]_c [2]), 
            .I2(n30671), .I3(GND_net), .O(n59415));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1521.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1522 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [5]), 
            .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1522.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_4_lut_adj_1523 (.I0(\data_in_frame[10] [5]), .I1(n28782), 
            .I2(n28299), .I3(\data_in_frame[12] [4]), .O(n28224));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1524 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [3]), 
            .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1524.LUT_INIT = 16'ha088;
    SB_LUT4 i51423_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[3]_c [1]), 
            .I2(n30671), .I3(GND_net), .O(n59453));   // verilog/coms.v(94[13:20])
    defparam i51423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(n29078), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [4]), .I3(\data_in_frame[9] [3]), .O(n28332));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 i19663_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n25151), .I3(GND_net), .O(n32453));
    defparam i19663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5605));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut (.I0(n28782), .I1(n4_adj_5597), .I2(n55742), 
            .I3(n28824), .O(n64121));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19868_3_lut (.I0(control_mode_c[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n25151), .I3(GND_net), .O(n32463));
    defparam i19868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19866_3_lut (.I0(control_mode_c[2]), .I1(\data_in_frame[1]_c [2]), 
            .I2(n25151), .I3(GND_net), .O(n32465));
    defparam i19866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20060_3_lut (.I0(\control_mode[1] ), .I1(\data_in_frame[1]_c [1]), 
            .I2(n25151), .I3(GND_net), .O(n32466));
    defparam i20060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2062));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19346_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n25082), .I3(GND_net), .O(n32473));
    defparam i19346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21447_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n25082), .I3(GND_net), .O(n32476));
    defparam i21447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1526 (.I0(\data_in_frame[1]_c [1]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[5] [3]), .O(n60459));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i18905_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6]_c [5]), 
            .I2(n25082), .I3(GND_net), .O(n32485));
    defparam i18905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18915_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6]_c [4]), 
            .I2(n25082), .I3(GND_net), .O(n32486));
    defparam i18915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2061));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1527 (.I0(\data_in_frame[1]_c [1]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[3]_c [2]), .O(n60528));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 equal_314_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_5670));   // verilog/coms.v(157[7:23])
    defparam equal_314_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1528 (.I0(n28836), .I1(n4_adj_5467), .I2(\data_in_frame[15] [7]), 
            .I3(n60435), .O(n62101));
    defparam i2_3_lut_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i22817_4_lut (.I0(n8), .I1(\FRAME_MATCHER.i [31]), .I2(n27746), 
            .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i22817_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i23079_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(GND_net), .O(n41173));
    defparam i23079_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i41564_2_lut_3_lut (.I0(n3489), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n61010));
    defparam i41564_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1529 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(n55744), .I3(\data_out_frame[19] [3]), .O(n6_adj_5667));
    defparam i1_2_lut_3_lut_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1530 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(n55793), .I3(GND_net), .O(n60435));
    defparam i1_2_lut_3_lut_adj_1530.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_3_lut_4_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [2]), .I3(n60365), .O(n12_adj_5624));   // verilog/coms.v(88[17:63])
    defparam i4_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1531 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(\FRAME_MATCHER.i [5]), .O(n65));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1531.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1532 (.I0(\FRAME_MATCHER.i [4]), .I1(n27873), .I2(GND_net), 
            .I3(GND_net), .O(n27746));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1532.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1533 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n39602), .O(n30627));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1533.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1534 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n59771), .O(n59773));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1534.LUT_INIT = 16'hfffd;
    SB_LUT4 i48717_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n79), .O(n67698));   // verilog/coms.v(157[7:23])
    defparam i48717_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1535 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[6] [1]), .O(n28024));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1536 (.I0(Kp_23__N_748), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n55362));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1536.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1537 (.I0(\data_out_frame[20] [3]), .I1(n55464), 
            .I2(n60523), .I3(n54865), .O(n54974));
    defparam i1_2_lut_3_lut_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1538 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n27855), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n4_adj_5657));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1538.LUT_INIT = 16'hfff4;
    SB_LUT4 equal_305_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam equal_305_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i22815_4_lut (.I0(n5_adj_5672), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i22815_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i2_3_lut_4_lut_adj_1539 (.I0(\FRAME_MATCHER.i [4]), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(\FRAME_MATCHER.i [3]), 
            .O(n89));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1539.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1540 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1]_c [2]), 
            .I2(\data_in_frame[3]_c [4]), .I3(n60377), .O(n28357));
    defparam i1_2_lut_3_lut_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1541 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(n28715), .O(n54798));
    defparam i1_2_lut_3_lut_4_lut_adj_1541.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n60058));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut_4_lut_adj_1542 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[17]_c [4]), .I3(\data_in_frame[15] [2]), 
            .O(n64103));
    defparam i1_3_lut_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1543 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n60721));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1543.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1544 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n60361));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1544.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_adj_1545 (.I0(n27855), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n29976));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut_adj_1545.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1546 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n25071));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1546.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_1547 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n60888));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1548 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n55300), .I3(n55895), .O(n55754));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i32_3_lut (.I0(n30669), .I1(rx_data[0]), .I2(\data_in_frame[2]_c [0]), 
            .I3(GND_net), .O(n24_adj_5604));   // verilog/coms.v(94[13:20])
    defparam i32_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i2_4_lut_adj_1549 (.I0(n4452), .I1(n25071), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n29976), .O(n62594));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1549.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1550 (.I0(n27864), .I1(n1970), .I2(n1968), .I3(n62594), 
            .O(n29417));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1550.LUT_INIT = 16'hbaaa;
    SB_LUT4 i22629_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n40721));
    defparam i22629_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5673));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1552 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5674));
    defparam i1_4_lut_adj_1552.LUT_INIT = 16'ha8a0;
    SB_LUT4 i23111_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5674), .I3(n4_adj_5673), .O(n41206));
    defparam i23111_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i2_2_lut_adj_1553 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5675));
    defparam i2_2_lut_adj_1553.LUT_INIT = 16'heeee;
    SB_LUT4 i13631_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n31822));   // verilog/coms.v(130[12] 305[6])
    defparam i13631_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13512_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n31703));   // verilog/coms.v(130[12] 305[6])
    defparam i13512_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1554 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5676));
    defparam i6_4_lut_adj_1554.LUT_INIT = 16'hfeff;
    SB_LUT4 i13632_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n31823));   // verilog/coms.v(130[12] 305[6])
    defparam i13632_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13633_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n31824));   // verilog/coms.v(130[12] 305[6])
    defparam i13633_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13634_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n31825));   // verilog/coms.v(130[12] 305[6])
    defparam i13634_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1555 (.I0(\data_in[3] [6]), .I1(n14_adj_5676), 
            .I2(n10_adj_5675), .I3(\data_in[2] [1]), .O(n27904));
    defparam i7_4_lut_adj_1555.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1556 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n27904), .I3(\data_in[0] [5]), .O(n20_adj_5677));
    defparam i8_4_lut_adj_1556.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1557 (.I0(n27759), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5678));
    defparam i7_4_lut_adj_1557.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_4_lut_adj_1558 (.I0(n38177), .I1(\control_mode[1] ), 
            .I2(\control_mode[0] ), .I3(control_update), .O(n30039));   // verilog/coms.v(130[12] 305[6])
    defparam i1_3_lut_4_lut_adj_1558.LUT_INIT = 16'hbf00;
    SB_LUT4 i13635_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n31826));   // verilog/coms.v(130[12] 305[6])
    defparam i13635_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19646_3_lut (.I0(n30709), .I1(rx_data[0]), .I2(\data_in_frame[22]_c [0]), 
            .I3(GND_net), .O(n32624));   // verilog/coms.v(94[13:20])
    defparam i19646_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_4_lut_adj_1559 (.I0(\data_in_frame[21][7] ), .I1(n30619), 
            .I2(n30708), .I3(rx_data[7]), .O(n59305));
    defparam i12_4_lut_adj_1559.LUT_INIT = 16'h3a0a;
    SB_LUT4 i14_4_lut_adj_1560 (.I0(\data_in_frame[21] [6]), .I1(n61124), 
            .I2(n30708), .I3(rx_data[6]), .O(n59297));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1560.LUT_INIT = 16'h3a0a;
    SB_LUT4 i44967_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [3]), .O(n64453));
    defparam i44967_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i13636_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n31827));   // verilog/coms.v(130[12] 305[6])
    defparam i13636_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13637_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n31828));   // verilog/coms.v(130[12] 305[6])
    defparam i13637_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_3_lut_adj_1561 (.I0(n64453), .I1(n19_adj_5678), .I2(n20_adj_5677), 
            .I3(GND_net), .O(n1964));
    defparam i11_3_lut_adj_1561.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1562 (.I0(\data_in[2] [4]), .I1(n27904), .I2(n28014), 
            .I3(\data_in[1] [5]), .O(n18_adj_5679));
    defparam i7_4_lut_adj_1562.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1563 (.I0(\data_in[0] [6]), .I1(n18_adj_5679), 
            .I2(\data_in[3] [0]), .I3(n27913), .O(n20_adj_5680));
    defparam i9_4_lut_adj_1563.LUT_INIT = 16'hfffd;
    SB_LUT4 i13638_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n31829));   // verilog/coms.v(130[12] 305[6])
    defparam i13638_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13639_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n31830));   // verilog/coms.v(130[12] 305[6])
    defparam i13639_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13640_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n31831));   // verilog/coms.v(130[12] 305[6])
    defparam i13640_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13641_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n31832));   // verilog/coms.v(130[12] 305[6])
    defparam i13641_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13642_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n31833));   // verilog/coms.v(130[12] 305[6])
    defparam i13642_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13643_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n31834));   // verilog/coms.v(130[12] 305[6])
    defparam i13643_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13644_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n31835));   // verilog/coms.v(130[12] 305[6])
    defparam i13644_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13645_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n31836));   // verilog/coms.v(130[12] 305[6])
    defparam i13645_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13646_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n31837));   // verilog/coms.v(130[12] 305[6])
    defparam i13646_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13647_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n31838));   // verilog/coms.v(130[12] 305[6])
    defparam i13647_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1564 (.I0(n38177), .I1(\control_mode[1] ), 
            .I2(\control_mode[0] ), .I3(GND_net), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1564.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1565 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18]_c [4]), 
            .I2(\data_in_frame[18][5] ), .I3(GND_net), .O(n60673));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1565.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5682));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1566 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18]_c [4]), 
            .I2(\data_in_frame[20] [5]), .I3(GND_net), .O(n60147));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1566.LUT_INIT = 16'h9696;
    SB_LUT4 i13648_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n31839));   // verilog/coms.v(130[12] 305[6])
    defparam i13648_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13649_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n31840));   // verilog/coms.v(130[12] 305[6])
    defparam i13649_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13650_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n31841));   // verilog/coms.v(130[12] 305[6])
    defparam i13650_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13651_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n31842));   // verilog/coms.v(130[12] 305[6])
    defparam i13651_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1567 (.I0(n15_adj_5682), .I1(n20_adj_5680), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1967));
    defparam i10_4_lut_adj_1567.LUT_INIT = 16'hfeff;
    SB_LUT4 i13652_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n31843));   // verilog/coms.v(130[12] 305[6])
    defparam i13652_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13653_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n31844));   // verilog/coms.v(130[12] 305[6])
    defparam i13653_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13654_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n31845));   // verilog/coms.v(130[12] 305[6])
    defparam i13654_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13655_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n31846));   // verilog/coms.v(130[12] 305[6])
    defparam i13655_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1568 (.I0(\data_in[3] [2]), .I1(\data_in[2] [0]), 
            .I2(\data_in[1] [2]), .I3(\data_in[1] [6]), .O(n10_adj_5683));
    defparam i4_4_lut_adj_1568.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(\data_in[0] [1]), .I1(\data_in[3] [7]), 
            .I2(n10_adj_5683), .I3(\data_in[2] [6]), .O(n6_adj_5684));   // verilog/coms.v(139[7:86])
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'hfbff;
    SB_LUT4 i13656_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n31847));   // verilog/coms.v(130[12] 305[6])
    defparam i13656_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13661_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n31852));   // verilog/coms.v(130[12] 305[6])
    defparam i13661_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13660_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n31851));   // verilog/coms.v(130[12] 305[6])
    defparam i13660_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13659_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n31850));   // verilog/coms.v(130[12] 305[6])
    defparam i13659_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1570 (.I0(\data_in[0] [5]), .I1(\data_in[1] [3]), 
            .I2(\data_in[2] [5]), .I3(n6_adj_5684), .O(n27913));   // verilog/coms.v(139[7:86])
    defparam i4_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1571 (.I0(n62765), .I1(\data_in_frame[19] [4]), 
            .I2(n28505), .I3(GND_net), .O(n60295));
    defparam i1_2_lut_3_lut_adj_1571.LUT_INIT = 16'h6969;
    SB_LUT4 i11_3_lut_adj_1572 (.I0(\data_in_frame[18]_c [4]), .I1(rx_data[4]), 
            .I2(n30702), .I3(GND_net), .O(n59161));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1572.LUT_INIT = 16'hcaca;
    SB_LUT4 i13658_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n31849));   // verilog/coms.v(130[12] 305[6])
    defparam i13658_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13657_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n31848));   // verilog/coms.v(130[12] 305[6])
    defparam i13657_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1573 (.I0(n62765), .I1(\data_in_frame[19] [4]), 
            .I2(n62188), .I3(\data_in_frame[19] [5]), .O(n60688));
    defparam i2_3_lut_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1574 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5685));
    defparam i4_4_lut_adj_1574.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1575 (.I0(\data_in[3] [4]), .I1(n10_adj_5685), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n28014));
    defparam i5_3_lut_adj_1575.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1576 (.I0(\data_in_frame[19] [3]), .I1(n62765), 
            .I2(n60587), .I3(n60162), .O(n26256));
    defparam i1_2_lut_3_lut_4_lut_adj_1576.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1577 (.I0(\data_in[0] [3]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [0]), .I3(GND_net), .O(n14_adj_5686));
    defparam i5_3_lut_adj_1577.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1578 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(n28014), .I3(\data_in[1] [5]), .O(n15_adj_5687));
    defparam i6_4_lut_adj_1578.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1579 (.I0(n15_adj_5687), .I1(\data_in[1] [0]), 
            .I2(n14_adj_5686), .I3(\data_in[2] [2]), .O(n27759));
    defparam i8_4_lut_adj_1579.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1580 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n27759), .O(n16_adj_5688));
    defparam i6_4_lut_adj_1580.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1581 (.I0(\control_mode[1] ), .I1(n38177), 
            .I2(\control_mode[0] ), .I3(GND_net), .O(n15_adj_6));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1581.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1582 (.I0(\control_mode[1] ), .I1(n38177), 
            .I2(\control_mode[0] ), .I3(GND_net), .O(n15_adj_7));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1582.LUT_INIT = 16'hefef;
    SB_LUT4 i7_4_lut_adj_1583 (.I0(n27913), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [3]), .O(n17_adj_5691));
    defparam i7_4_lut_adj_1583.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\current[15] ), 
            .I2(\data_out_frame[21] [7]), .I3(\FRAME_MATCHER.i_31__N_2509 ), 
            .O(n26));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd800;
    SB_LUT4 i9_4_lut_adj_1584 (.I0(n17_adj_5691), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5688), .I3(\data_in[3] [1]), .O(n1970));
    defparam i9_4_lut_adj_1584.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_4_lut_4_lut_adj_1585 (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I1(\current[15] ), .I2(\data_out_frame[21] [5]), .I3(\FRAME_MATCHER.i_31__N_2509 ), 
            .O(n2_adj_5352));
    defparam i1_4_lut_4_lut_adj_1585.LUT_INIT = 16'hd800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64823), .I3(n64821), .O(n7));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i366_2_lut (.I0(n1967), .I1(n1964), .I2(GND_net), .I3(GND_net), 
            .O(n1968));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64865), .I3(n64863), .O(n7_adj_5401));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1586 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n35070));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1586.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n64811), .I3(n64809), .O(n7_adj_5359));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_4_lut_adj_1587 (.I0(n41206), .I1(n62063), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n40721), .O(n6_adj_5693));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1587.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1588 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n61010), .O(n79));
    defparam i3_4_lut_adj_1588.LUT_INIT = 16'hefff;
    SB_LUT4 i1_3_lut_4_lut_adj_1589 (.I0(\data_in_frame[18][7] ), .I1(\data_in_frame[18] [6]), 
            .I2(n60274), .I3(n60673), .O(n61920));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1589.LUT_INIT = 16'h6996;
    SB_LUT4 i12519_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n40778), 
            .I2(n39602), .I3(reset), .O(n30709));   // verilog/coms.v(157[7:23])
    defparam i12519_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i3_4_lut_adj_1590 (.I0(n35070), .I1(n6_adj_5693), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n71718));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1590.LUT_INIT = 16'hefee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1591 (.I0(\FRAME_MATCHER.i[0] ), .I1(n40778), 
            .I2(n61010), .I3(n10_adj_5670), .O(n30637));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1591.LUT_INIT = 16'hffbf;
    SB_LUT4 i12_4_lut_adj_1592 (.I0(\data_in_frame[17]_c [4]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[4]), .O(n59233));
    defparam i12_4_lut_adj_1592.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1593 (.I0(\FRAME_MATCHER.i [5]), .I1(n89), 
            .I2(n3489), .I3(GND_net), .O(n39602));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1593.LUT_INIT = 16'h4040;
    SB_LUT4 i12_4_lut_adj_1594 (.I0(\data_in_frame[17]_c [3]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[3]), .O(n59237));
    defparam i12_4_lut_adj_1594.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1595 (.I0(\data_in_frame[17]_c [2]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[2]), .O(n59251));
    defparam i12_4_lut_adj_1595.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1596 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n60118), .I3(GND_net), .O(n60119));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1596.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1597 (.I0(\data_in_frame[18][7] ), .I1(\data_in_frame[18] [6]), 
            .I2(n28517), .I3(GND_net), .O(n60385));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1597.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1598 (.I0(\data_in_frame[17]_c [1]), .I1(n30627), 
            .I2(n30700), .I3(rx_data[1]), .O(n59247));
    defparam i12_4_lut_adj_1598.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1599 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3489));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1599.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1600 (.I0(\FRAME_MATCHER.i [5]), .I1(n89), 
            .I2(n3489), .I3(n8_c), .O(n30635));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1600.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1601 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[1] ), 
            .I2(\FRAME_MATCHER.i[2] ), .I3(n59771), .O(n59779));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1601.LUT_INIT = 16'hffbf;
    SB_LUT4 i2_3_lut_4_lut_adj_1602 (.I0(n1967), .I1(n1964), .I2(n1970), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n62063));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1602.LUT_INIT = 16'h8000;
    SB_LUT4 i14_4_lut_adj_1603 (.I0(\data_in_frame[17]_c [0]), .I1(n7_adj_5694), 
            .I2(n30700), .I3(n4_adj_5695), .O(n59223));   // verilog/coms.v(94[13:20])
    defparam i14_4_lut_adj_1603.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_adj_1604 (.I0(n60584), .I1(n60807), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[14] [6]), .O(n60245));
    defparam i1_2_lut_4_lut_adj_1604.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1605 (.I0(n60584), .I1(n60807), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[16] [5]), .O(n60747));
    defparam i1_2_lut_4_lut_adj_1605.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5602));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1606 (.I0(\data_in_frame[14] [2]), .I1(n62168), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n60420));
    defparam i1_2_lut_3_lut_adj_1606.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1607 (.I0(\data_in_frame[14] [2]), .I1(n62168), 
            .I2(n62398), .I3(GND_net), .O(n27587));
    defparam i1_2_lut_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i45327_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64822));
    defparam i45327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45328_4_lut (.I0(n64822), .I1(n60052), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n64823));
    defparam i45328_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i45326_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64821));
    defparam i45326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5586));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1608 (.I0(n28745), .I1(n29047), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n60596));
    defparam i2_3_lut_4_lut_adj_1608.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [3]), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_4_lut_adj_1610 (.I0(\data_in_frame[19] [3]), .I1(n60810), 
            .I2(n60295), .I3(\data_in_frame[21][5] ), .O(n60851));
    defparam i2_3_lut_4_lut_adj_1610.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1611 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n41206), .O(n27855));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1611.LUT_INIT = 16'ha8aa;
    SB_LUT4 select_787_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5576));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'ha088;
    SB_LUT4 select_789_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5579));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1613 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n28809), .I3(\data_in_frame[14] [0]), .O(n28677));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1613.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_4_lut_adj_1614 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27873), .I3(\FRAME_MATCHER.i[1] ), .O(n5_adj_5672));
    defparam i1_3_lut_4_lut_adj_1614.LUT_INIT = 16'hfefc;
    SB_LUT4 select_789_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 n71331_bdd_4_lut (.I0(n71331), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(byte_transmit_counter[1]), 
            .O(n71334));
    defparam n71331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1615 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n60118));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1615.LUT_INIT = 16'hfefe;
    SB_LUT4 i12118_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3489), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n30308));   // verilog/coms.v(158[12:15])
    defparam i12118_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 select_787_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1616 (.I0(n28836), .I1(\data_in_frame[12] [5]), 
            .I2(n28392), .I3(\data_in_frame[13] [0]), .O(n60462));
    defparam i1_2_lut_3_lut_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5572));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5571));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5570));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5569));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_787_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5568));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5567));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1617 (.I0(\data_in_frame[8] [3]), .I1(n60538), 
            .I2(n4_adj_5597), .I3(\data_in_frame[10] [4]), .O(n28392));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5566));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(n60773), .I1(n28812), .I2(\data_in_frame[9] [2]), 
            .I3(\data_in_frame[11] [5]), .O(n11_adj_5574));   // verilog/coms.v(76[16:42])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5565));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5564));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_3_lut_4_lut (.I0(n60298), .I1(\data_out_frame[12] [1]), .I2(n62099), 
            .I3(\data_out_frame[18] [1]), .O(n23_c));
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5563));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5562));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1618 (.I0(\data_out_frame[21] [2]), .I1(n28907), 
            .I2(n55567), .I3(GND_net), .O(n60499));
    defparam i1_2_lut_3_lut_adj_1618.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1619 (.I0(n55179), .I1(n55783), .I2(\data_out_frame[16] [0]), 
            .I3(\data_out_frame[16] [1]), .O(n6_adj_5666));
    defparam i1_2_lut_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5561));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1620 (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[20] [3]), 
            .I2(n26026), .I3(n54865), .O(n54978));
    defparam i1_2_lut_4_lut_adj_1620.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(n55783), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n60858));
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5560));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1622 (.I0(\data_out_frame[12] [5]), .I1(n1519), 
            .I2(\data_out_frame[14] [7]), .I3(n60909), .O(n60646));
    defparam i1_2_lut_4_lut_adj_1622.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1623 (.I0(\data_out_frame[15] [4]), .I1(n28056), 
            .I2(n28615), .I3(GND_net), .O(n28460));
    defparam i1_2_lut_3_lut_adj_1623.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5559));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5558));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5557));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5556));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1624 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n60736));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1624.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5555));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5554));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [0]), 
            .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5553));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5552));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5551));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5550));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1626 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[6] [7]), .I3(n1168), .O(n60915));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5549));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5548));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5547));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5546));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5545));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1627 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[8][6] ), .I3(\data_out_frame[4] [2]), .O(n40_adj_5629));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5544));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5543));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1628 (.I0(n55746), .I1(\data_out_frame[23] [2]), 
            .I2(\data_out_frame[21] [0]), .I3(\data_out_frame[23] [3]), 
            .O(n60818));
    defparam i2_3_lut_4_lut_adj_1628.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1629 (.I0(\data_out_frame[13] [7]), .I1(n54834), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n54842));
    defparam i1_2_lut_3_lut_adj_1629.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_52008 (.I0(byte_transmit_counter[1]), 
            .I1(n64629), .I2(n64630), .I3(byte_transmit_counter[2]), .O(n71319));
    defparam byte_transmit_counter_1__bdd_4_lut_52008.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5542));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5541));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n7_adj_5650));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[14] [5]), 
            .I2(n1655), .I3(\data_out_frame[15] [0]), .O(n12_adj_5648));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n71319_bdd_4_lut (.I0(n71319), .I1(n64798), .I2(n64797), .I3(byte_transmit_counter[2]), 
            .O(n71322));
    defparam n71319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[12] [5]), 
            .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1631 (.I0(\data_out_frame[12] [1]), .I1(n62099), 
            .I2(n60206), .I3(GND_net), .O(n54970));
    defparam i1_2_lut_3_lut_adj_1631.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1632 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [3]), 
            .I2(n1513), .I3(n60744), .O(n29259));
    defparam i1_2_lut_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut (.I0(n1168), .I1(n60633), .I2(n10_adj_5635), 
            .I3(n28446), .O(n28745));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14102_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n32293));
    defparam i14102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14487_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n32678));
    defparam i14487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14490_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n32681));
    defparam i14490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5527));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14493_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n32684));
    defparam i14493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1633 (.I0(\data_out_frame[6] [6]), .I1(n60546), 
            .I2(\data_out_frame[6] [7]), .I3(n1168), .O(n29177));
    defparam i1_2_lut_4_lut_adj_1633.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1634 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[12] [7]), 
            .I2(n28968), .I3(GND_net), .O(n10_adj_5631));
    defparam i2_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14496_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n32687));
    defparam i14496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1635 (.I0(\data_out_frame[13] [7]), .I1(n54834), 
            .I2(n60815), .I3(GND_net), .O(n6_adj_5449));
    defparam i1_2_lut_3_lut_adj_1635.LUT_INIT = 16'h9696;
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[9] [6]), .O(n41_adj_5627));   // verilog/coms.v(78[16:27])
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1636 (.I0(n28024), .I1(\data_out_frame[8][3] ), 
            .I2(\data_out_frame[8][4] ), .I3(GND_net), .O(n60706));
    defparam i1_2_lut_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5521));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14499_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n32690));
    defparam i14499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13495_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n31686));
    defparam i13495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13492_3_lut_4_lut (.I0(n8), .I1(n60130), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n31683));
    defparam i13492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1637 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[10] [0]), 
            .I2(n28427), .I3(n60485), .O(n55800));
    defparam i1_3_lut_4_lut_adj_1637.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_4_lut_4_lut_adj_1638 (.I0(n41236), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n59159));
    defparam i11_4_lut_4_lut_adj_1638.LUT_INIT = 16'hfd20;
    SB_LUT4 i14300_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n32491));
    defparam i14300_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12140_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30330));   // verilog/coms.v(109[34:55])
    defparam i12140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1639 (.I0(n28024), .I1(n60345), .I2(n55800), 
            .I3(n60867), .O(n55856));
    defparam i1_2_lut_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i14225_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n32416));
    defparam i14225_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14222_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n32413));
    defparam i14222_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45369_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64864));
    defparam i45369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45370_4_lut (.I0(n64864), .I1(n30330), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n64865));
    defparam i45370_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 select_787_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1640 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [1]), 
            .I2(n10_adj_5621), .I3(n28888), .O(n27445));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1640.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i45368_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n64863));
    defparam i45368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(\data_in_frame[23] [5]), 
            .I3(rx_data[5]), .O(n59105));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i14068_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n32259));
    defparam i14068_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14071_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n32262));
    defparam i14071_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14031_3_lut_4_lut (.I0(n41236), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n32222));
    defparam i14031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5508));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1641 (.I0(n39602), .I1(\FRAME_MATCHER.i[0] ), 
            .I2(rx_data[0]), .I3(GND_net), .O(n4_adj_5695));
    defparam i1_2_lut_3_lut_adj_1641.LUT_INIT = 16'h8080;
    SB_LUT4 i48535_2_lut (.I0(n71586), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67792));
    defparam i48535_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5507));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1642 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n54742), .I3(GND_net), .O(n60417));
    defparam i1_2_lut_3_lut_adj_1642.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_71_i2_4_lut (.I0(\data_out_frame[8][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [1]), 
            .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_70_i2_4_lut (.I0(\data_out_frame[8][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_69_i2_4_lut (.I0(\data_out_frame[8][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_68_i2_4_lut (.I0(\data_out_frame[8][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_67_i2_4_lut (.I0(\data_out_frame[8][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_66_i2_4_lut (.I0(\data_out_frame[8][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_65_i2_4_lut (.I0(\data_out_frame[8][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1644 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[16] [5]), .I3(\data_out_frame[18] [6]), 
            .O(n6));
    defparam i1_2_lut_3_lut_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1645 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1] [4]), 
            .I2(n60488), .I3(\data_in_frame[3][5] ), .O(n60848));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1645.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13880_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n32071));
    defparam i13880_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14141_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n32332));
    defparam i14141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [6]), 
            .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'ha088;
    SB_LUT4 i13883_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n32074));
    defparam i13883_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5494));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13886_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n32077));
    defparam i13886_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5489));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1647 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n29010));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1647.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13889_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n32080));
    defparam i13889_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14138_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n32329));
    defparam i14138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14135_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n32326));
    defparam i14135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14132_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n32323));
    defparam i14132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14129_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n32320));
    defparam i14129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut_adj_1648 (.I0(n30621), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n59117));
    defparam i11_4_lut_4_lut_adj_1648.LUT_INIT = 16'hfe10;
    SB_LUT4 i14122_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n32313));
    defparam i14122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14119_3_lut_4_lut (.I0(n30621), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n32310));
    defparam i14119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut_adj_1649 (.I0(n30635), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n59243));
    defparam i11_4_lut_4_lut_adj_1649.LUT_INIT = 16'hfe10;
    SB_LUT4 i14162_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n32353));
    defparam i14162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14159_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n32350));
    defparam i14159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1650 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n60197));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1650.LUT_INIT = 16'h9696;
    SB_LUT4 i13892_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n32083));
    defparam i13892_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [3]), 
            .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'ha088;
    SB_LUT4 i14156_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n32347));
    defparam i14156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14153_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n32344));
    defparam i14153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14150_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n32341));
    defparam i14150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14147_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n32338));
    defparam i14147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14144_3_lut_4_lut (.I0(n30635), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n32335));
    defparam i14144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13539_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n31730));
    defparam i13539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13536_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n31727));
    defparam i13536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [7]), 
            .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'ha088;
    SB_LUT4 i13895_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n32086));
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51437_2_lut_3_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n70932));   // verilog/coms.v(99[12:25])
    defparam i51437_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13533_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n31724));
    defparam i13533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13898_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n32089));
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13530_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n31721));
    defparam i13530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1653 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1]_c [2]), 
            .I2(\data_in_frame[3]_c [4]), .I3(GND_net), .O(n28266));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1653.LUT_INIT = 16'h9696;
    SB_LUT4 i13901_3_lut_4_lut (.I0(n8_adj_8), .I1(n59771), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n32092));
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13527_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n31718));
    defparam i13527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n35070), .O(n6_adj_5603));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_4_lut_adj_1654 (.I0(n30655), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[1]_c [2]), .O(n59395));
    defparam i11_4_lut_4_lut_adj_1654.LUT_INIT = 16'hfe10;
    SB_LUT4 i13521_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[1]_c [1]), .O(n31712));
    defparam i13521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6][6] ), 
            .I2(\data_in_frame[6]_c [5]), .I3(GND_net), .O(n60217));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13518_3_lut_4_lut (.I0(n30655), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[1]_c [0]), .O(n31709));
    defparam i13518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1656 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n39603), .I3(\FRAME_MATCHER.i[0] ), .O(n30702));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1656.LUT_INIT = 16'h0020;
    SB_LUT4 i13092_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n31283));   // verilog/coms.v(130[12] 305[6])
    defparam i13092_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_787_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1657 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n60130), .I3(\FRAME_MATCHER.i[0] ), .O(n30669));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1657.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_4_lut_adj_1658 (.I0(\data_in_frame[6]_c [4]), .I1(Kp_23__N_875), 
            .I2(Kp_23__N_878), .I3(\data_in_frame[6]_c [5]), .O(Kp_23__N_974));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1659 (.I0(Kp_23__N_767), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[3] [0]), .O(n28947));   // verilog/coms.v(80[16:27])
    defparam i2_3_lut_4_lut_adj_1659.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1660 (.I0(\data_in_frame[5] [4]), .I1(n60528), 
            .I2(\data_in_frame[5] [5]), .I3(\data_in_frame[7] [6]), .O(n60377));
    defparam i1_2_lut_4_lut_adj_1660.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1661 (.I0(\data_in_frame[3]_c [6]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[1] [5]), .O(n60262));   // verilog/coms.v(18[27:29])
    defparam i2_3_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1662 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [6]), 
            .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1663 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [5]), 
            .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1663.LUT_INIT = 16'ha088;
    SB_LUT4 equal_304_i7_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5694));   // verilog/coms.v(157[7:23])
    defparam equal_304_i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_310_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_8));   // verilog/coms.v(157[7:23])
    defparam equal_310_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1664 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n39602), .I3(\FRAME_MATCHER.i[0] ), .O(n30623));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1664.LUT_INIT = 16'hffdf;
    SB_LUT4 select_787_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1665 (.I0(\data_in_frame[21][2] ), .I1(n55952), 
            .I2(n54912), .I3(\data_in_frame[23] [4]), .O(n62732));
    defparam i2_3_lut_4_lut_adj_1665.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1666 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [2]), 
            .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [0]), 
            .I2(\control_mode[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'ha088;
    SB_LUT4 i48689_2_lut (.I0(n71598), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67740));
    defparam i48689_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [7]), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_adj_1669 (.I0(n55903), .I1(\data_in_frame[15] [5]), 
            .I2(n55754), .I3(\data_in_frame[17][6] ), .O(n60679));
    defparam i1_2_lut_4_lut_adj_1669.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1670 (.I0(\data_in_frame[7] [1]), .I1(n55176), 
            .I2(n10_adj_5584), .I3(\data_in_frame[11] [5]), .O(n60759));
    defparam i5_3_lut_4_lut_adj_1670.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [6]), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1672 (.I0(\data_in_frame[10] [0]), .I1(n60561), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n60807));
    defparam i1_2_lut_3_lut_adj_1672.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1673 (.I0(\data_in_frame[8] [1]), .I1(n28249), 
            .I2(n10_adj_5577), .I3(\data_in_frame[5] [6]), .O(n54800));
    defparam i5_3_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1674 (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(n59771), .I3(\FRAME_MATCHER.i[0] ), .O(n59772));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1674.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_3_lut_adj_1675 (.I0(\data_out_frame[16] [3]), .I1(n62023), 
            .I2(\data_out_frame[21] [1]), .I3(GND_net), .O(n60352));
    defparam i1_2_lut_3_lut_adj_1675.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1676 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[3]_c [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[8] [1]), .O(n60314));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1] [5]), 
            .I2(n60184), .I3(GND_net), .O(n60203));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1678 (.I0(\data_out_frame[16] [3]), .I1(n62023), 
            .I2(n54970), .I3(GND_net), .O(n60900));
    defparam i1_2_lut_3_lut_adj_1678.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1679 (.I0(n28337), .I1(n28266), .I2(n60377), 
            .I3(Kp_23__N_1085), .O(n60561));
    defparam i1_2_lut_4_lut_adj_1679.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1680 (.I0(n28337), .I1(n28266), .I2(n60377), 
            .I3(GND_net), .O(n28824));
    defparam i1_2_lut_3_lut_adj_1680.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1681 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(n28213), .I3(n28299), .O(n64095));
    defparam i1_3_lut_4_lut_adj_1681.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1682 (.I0(n29193), .I1(\data_in_frame[8] [7]), 
            .I2(Kp_23__N_993), .I3(\data_in_frame[8] [6]), .O(n29250));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13077_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n31268));   // verilog/coms.v(130[12] 305[6])
    defparam i13077_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i51593_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n41206), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i51593_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 select_787_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1683 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(n60921), .O(n60827));
    defparam i1_2_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1684 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_974), .I3(GND_net), .O(n28122));
    defparam i1_2_lut_3_lut_adj_1684.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1685 (.I0(n55903), .I1(n60897), .I2(\data_in_frame[17] [7]), 
            .I3(\data_in_frame[17][6] ), .O(n60339));
    defparam i2_3_lut_4_lut_adj_1685.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51801 (.I0(byte_transmit_counter[1]), 
            .I1(n64827), .I2(n64828), .I3(byte_transmit_counter[2]), .O(n71289));
    defparam byte_transmit_counter_1__bdd_4_lut_51801.LUT_INIT = 16'he4aa;
    SB_LUT4 n71289_bdd_4_lut (.I0(n71289), .I1(n64621), .I2(n64620), .I3(byte_transmit_counter[2]), 
            .O(n71292));
    defparam n71289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51810 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[20] [2]), .I2(\data_out_frame[21] [2]), 
            .I3(byte_transmit_counter[4]), .O(n71283));
    defparam byte_transmit_counter_0__bdd_4_lut_51810.LUT_INIT = 16'he4aa;
    SB_LUT4 n71283_bdd_4_lut (.I0(n71283), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[4] [2]), .I3(byte_transmit_counter[4]), 
            .O(n71286));
    defparam n71283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51776 (.I0(byte_transmit_counter[1]), 
            .I1(n64866), .I2(n64867), .I3(byte_transmit_counter[2]), .O(n71277));
    defparam byte_transmit_counter_1__bdd_4_lut_51776.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1686 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n60329));
    defparam i1_2_lut_3_lut_adj_1686.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1687 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1964), .I3(n1967), .O(n27864));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1687.LUT_INIT = 16'h4000;
    SB_LUT4 i49200_2_lut (.I0(n71610), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67748));
    defparam i49200_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1688 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(n55291), .I3(n26026), .O(n55740));
    defparam i2_3_lut_4_lut_adj_1688.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1689 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[16] [2]), 
            .I2(n60694), .I3(n26207), .O(n54794));
    defparam i2_3_lut_4_lut_adj_1689.LUT_INIT = 16'h6996;
    SB_LUT4 i12133_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30323));   // verilog/coms.v(109[34:55])
    defparam i12133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1690 (.I0(\data_in_frame[19] [6]), .I1(n62765), 
            .I2(\data_in_frame[19] [4]), .I3(n28505), .O(n60621));
    defparam i1_2_lut_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1691 (.I0(n28332), .I1(n60721), .I2(n60827), 
            .I3(GND_net), .O(n60756));
    defparam i1_2_lut_3_lut_adj_1691.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1692 (.I0(\data_in_frame[12] [6]), .I1(n28213), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[10] [7]), .O(n6_adj_5472));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1692.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1693 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[14] [2]), 
            .I2(n62168), .I3(n28677), .O(n60676));
    defparam i1_2_lut_4_lut_adj_1693.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1694 (.I0(n28548), .I1(\data_in_frame[14] [2]), 
            .I2(n62168), .I3(\data_in_frame[16] [4]), .O(n28517));
    defparam i1_2_lut_4_lut_adj_1694.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13789_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n31980));
    defparam i13789_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13793_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n31984));
    defparam i13793_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1695 (.I0(\data_out_frame[20] [2]), .I1(n55737), 
            .I2(\data_out_frame[22] [3]), .I3(n60291), .O(n61840));
    defparam i2_3_lut_4_lut_adj_1695.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1696 (.I0(n60652), .I1(n10_adj_5468), .I2(n61964), 
            .I3(n60602), .O(n64151));
    defparam i1_2_lut_4_lut_adj_1696.LUT_INIT = 16'h9669;
    SB_LUT4 i13796_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n31987));
    defparam i13796_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1697 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[14] [5]), .I3(GND_net), .O(n60174));
    defparam i1_2_lut_3_lut_adj_1697.LUT_INIT = 16'h9696;
    SB_LUT4 i13799_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n31990));
    defparam i13799_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71277_bdd_4_lut (.I0(n71277), .I1(n64885), .I2(n64884), .I3(byte_transmit_counter[2]), 
            .O(n71280));
    defparam n71277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1698 (.I0(\data_out_frame[20] [2]), .I1(n55737), 
            .I2(n26026), .I3(\data_out_frame[20] [3]), .O(n55879));
    defparam i1_2_lut_3_lut_4_lut_adj_1698.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12089_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n30278));   // verilog/coms.v(109[34:55])
    defparam i12089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1699 (.I0(n55903), .I1(\data_in_frame[15] [5]), 
            .I2(n55754), .I3(GND_net), .O(n28130));
    defparam i1_2_lut_3_lut_adj_1699.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n64817), .I1(n64815), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n7_c));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i13802_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n31993));
    defparam i13802_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13805_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n31996));
    defparam i13805_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1700 (.I0(n29204), .I1(\data_in_frame[14] [7]), 
            .I2(n60200), .I3(\data_in_frame[12] [6]), .O(n61788));
    defparam i2_3_lut_4_lut_adj_1700.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48729_2_lut (.I0(n71634), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n67736));
    defparam i48729_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50225_3_lut (.I0(n71604), .I1(n71334), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n69720));
    defparam i50225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13808_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n31999));
    defparam i13808_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13811_3_lut_4_lut (.I0(n8), .I1(n59771), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n32002));
    defparam i13811_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1701 (.I0(\data_in_frame[18][1] ), .I1(\data_in_frame[18][3] ), 
            .I2(\data_in_frame[18][0] ), .I3(\data_in_frame[17] [5]), .O(n64159));
    defparam i1_3_lut_4_lut_adj_1701.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1702 (.I0(n55428), .I1(\data_in_frame[17]_c [0]), 
            .I2(n60587), .I3(\data_in_frame[19] [2]), .O(n60162));
    defparam i2_3_lut_4_lut_adj_1702.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1703 (.I0(n54824), .I1(n28548), .I2(n10_adj_5466), 
            .I3(n55864), .O(n54869));
    defparam i5_3_lut_4_lut_adj_1703.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1704 (.I0(n54869), .I1(n60385), .I2(\data_in_frame[19] [0]), 
            .I3(n29130), .O(n55952));
    defparam i1_2_lut_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1705 (.I0(n28548), .I1(n60873), .I2(n60747), 
            .I3(n60731), .O(n6_adj_5465));
    defparam i1_2_lut_4_lut_adj_1705.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1706 (.I0(\data_in_frame[0] [5]), .I1(n28715), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[0] [6]), .O(n22_adj_5698));
    defparam i5_4_lut_adj_1706.LUT_INIT = 16'h1221;
    SB_LUT4 select_787_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_51771 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[4]), .O(n71271));
    defparam byte_transmit_counter_0__bdd_4_lut_51771.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1707 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(n60879), .I3(GND_net), .O(n60703));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1707.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1708 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n60445));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1709 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(\data_out_frame[14] [4]), .I3(GND_net), .O(n60374));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1709.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_adj_1710 (.I0(n32_adj_5590), .I1(Kp_23__N_748), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n20_adj_5699));
    defparam i3_3_lut_adj_1710.LUT_INIT = 16'h1414;
    SB_LUT4 n71271_bdd_4_lut (.I0(n71271), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[6] [2]), .I3(byte_transmit_counter[4]), 
            .O(n71274));
    defparam n71271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1711 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n60744), .I3(GND_net), .O(n1655));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1711.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1712 (.I0(n60349), .I1(n10_adj_5663), .I2(\data_out_frame[6] [1]), 
            .I3(n1519), .O(n28456));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1712.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1713 (.I0(\data_out_frame[21] [5]), .I1(n55907), 
            .I2(n10_adj_5456), .I3(n55796), .O(n60682));
    defparam i5_3_lut_4_lut_adj_1713.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1714 (.I0(n60349), .I1(n10_adj_5663), .I2(\data_out_frame[6] [1]), 
            .I3(\data_out_frame[12] [4]), .O(n60744));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1714.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1715 (.I0(\data_out_frame[15] [4]), .I1(n28056), 
            .I2(n28615), .I3(n60153), .O(n60154));
    defparam i1_2_lut_4_lut_adj_1715.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1716 (.I0(n1964), .I1(n4452), .I2(n1967), 
            .I3(n1970), .O(n61999));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1716.LUT_INIT = 16'h2000;
    SB_LUT4 select_787_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1964), .I1(n4452), .I2(n4_adj_5657), 
            .I3(\FRAME_MATCHER.i_31__N_2514 ), .O(n62119));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i2_3_lut_4_lut_adj_1717 (.I0(\data_out_frame[17] [5]), .I1(n28056), 
            .I2(n62343), .I3(\data_out_frame[15] [3]), .O(n60153));
    defparam i2_3_lut_4_lut_adj_1717.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1718 (.I0(\data_out_frame[4] [0]), .I1(n60618), 
            .I2(\data_out_frame[10] [6]), .I3(n1130), .O(n14_adj_5633));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1718.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1719 (.I0(\FRAME_MATCHER.i[0] ), .I1(n7_adj_5694), 
            .I2(n61010), .I3(n10_adj_5670), .O(n30655));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1719.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_3_lut_adj_1720 (.I0(\data_out_frame[18] [3]), .I1(n61794), 
            .I2(n55464), .I3(GND_net), .O(n28483));
    defparam i1_2_lut_3_lut_adj_1720.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1721 (.I0(\data_out_frame[15] [5]), .I1(n55577), 
            .I2(n28615), .I3(GND_net), .O(n55783));
    defparam i1_2_lut_3_lut_adj_1721.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1722 (.I0(\data_out_frame[15] [5]), .I1(n55577), 
            .I2(n28056), .I3(\data_out_frame[15] [4]), .O(n55830));
    defparam i1_2_lut_3_lut_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1723 (.I0(\data_out_frame[13] [6]), .I1(n28745), 
            .I2(n54796), .I3(GND_net), .O(n60815));
    defparam i1_2_lut_3_lut_adj_1723.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1724 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n28446));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1724.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1725 (.I0(\data_out_frame[13] [7]), .I1(n54834), 
            .I2(\data_out_frame[15] [7]), .I3(n60596), .O(n6_adj_5448));
    defparam i1_2_lut_4_lut_adj_1725.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_2_lut_4_lut_adj_1726 (.I0(n55760), .I1(n60298), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[21] [6]), .O(n15_c));
    defparam i4_2_lut_4_lut_adj_1726.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1727 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n60633));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1727.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1728 (.I0(n37239), .I1(n22_adj_5698), .I2(\data_in_frame[0] [7]), 
            .I3(n60248), .O(n28_adj_5700));
    defparam i11_4_lut_adj_1728.LUT_INIT = 16'h0440;
    SB_LUT4 select_787_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1729 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1]_c [1]), .I3(\data_in_frame[1]_c [2]), 
            .O(n26_adj_5701));
    defparam i9_4_lut_adj_1729.LUT_INIT = 16'h8400;
    SB_LUT4 i8_4_lut_adj_1730 (.I0(n70932), .I1(\data_in_frame[2]_c [0]), 
            .I2(\data_in_frame[0] [0]), .I3(Kp_23__N_748), .O(n25_adj_5702));
    defparam i8_4_lut_adj_1730.LUT_INIT = 16'h1441;
    SB_LUT4 i12_4_lut_adj_1731 (.I0(n28690), .I1(n28157), .I2(n55362), 
            .I3(\data_in_frame[1] [5]), .O(n29_adj_5703));
    defparam i12_4_lut_adj_1731.LUT_INIT = 16'h1000;
    SB_LUT4 i14_4_lut_adj_1732 (.I0(\data_in_frame[1]_c [3]), .I1(n28_adj_5700), 
            .I2(n20_adj_5699), .I3(\data_in_frame[1] [6]), .O(n31_adj_5704));
    defparam i14_4_lut_adj_1732.LUT_INIT = 16'h8000;
    SB_LUT4 i16_4_lut_adj_1733 (.I0(n31_adj_5704), .I1(n29_adj_5703), .I2(n25_adj_5702), 
            .I3(n26_adj_5701), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1733.LUT_INIT = 16'h8000;
    SB_LUT4 select_787_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[25] [1]), .I1(n54978), .I2(n55802), 
            .I3(\data_out_frame[25] [2]), .O(n8_adj_5637));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1734 (.I0(\data_out_frame[25] [1]), .I1(n54978), 
            .I2(n55879), .I3(\data_out_frame[22] [4]), .O(n8_adj_5649));
    defparam i3_3_lut_4_lut_adj_1734.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1735 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[7] [4]), .O(n60317));
    defparam i2_3_lut_4_lut_adj_1735.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1736 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [3]), 
            .I2(n28446), .I3(n28020), .O(n1312));
    defparam i2_3_lut_4_lut_adj_1736.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i41582_3_lut_4_lut (.I0(n10_adj_5670), .I1(n61010), .I2(n8_adj_8), 
            .I3(reset), .O(n30671));
    defparam i41582_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1737 (.I0(n60482), .I1(n54876), .I2(GND_net), 
            .I3(GND_net), .O(n60627));
    defparam i1_2_lut_3_lut_adj_1737.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_4_lut_adj_1738 (.I0(\data_out_frame[10] [1]), .I1(n60727), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[10] [6]), 
            .O(n60168));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1738.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1739 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [1]), .I3(\data_out_frame[20] [2]), 
            .O(n28961));
    defparam i1_2_lut_4_lut_adj_1739.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1740 (.I0(n10_adj_5670), .I1(n61010), .I2(reset), 
            .I3(GND_net), .O(n60130));
    defparam i1_2_lut_3_lut_adj_1740.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1741 (.I0(n60388), .I1(n10_adj_5625), .I2(n1563), 
            .I3(\data_out_frame[14] [2]), .O(n60427));
    defparam i1_2_lut_4_lut_adj_1741.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1742 (.I0(n60388), .I1(n10_adj_5625), .I2(n1563), 
            .I3(\data_out_frame[14] [2]), .O(n55985));
    defparam i1_2_lut_4_lut_adj_1742.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1743 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[17] [0]), .I3(n60374), .O(n60452));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1743.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1744 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(\data_out_frame[14] [3]), .I3(GND_net), .O(n60206));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1744.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1745 (.I0(\data_out_frame[12] [2]), .I1(n1510), 
            .I2(n55985), .I3(n60374), .O(n55748));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1745.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1746 (.I0(\data_out_frame[20] [0]), .I1(n55462), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n60482));
    defparam i1_2_lut_3_lut_adj_1746.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1747 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\data_out_frame[1][5] ), .I3(GND_net), .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1747.LUT_INIT = 16'ha8a8;
    SB_LUT4 i2_3_lut_4_lut_adj_1748 (.I0(n55273), .I1(n61794), .I2(\data_out_frame[18] [3]), 
            .I3(\data_out_frame[18] [4]), .O(n54792));
    defparam i2_3_lut_4_lut_adj_1748.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1749 (.I0(\data_out_frame[15] [6]), .I1(n55577), 
            .I2(n60778), .I3(GND_net), .O(n55760));
    defparam i1_2_lut_3_lut_adj_1749.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1750 (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[17] [6]), .I3(\data_out_frame[19] [7]), 
            .O(n6_c));
    defparam i1_2_lut_4_lut_adj_1750.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1751 (.I0(\data_out_frame[23] [5]), .I1(n62192), 
            .I2(n54859), .I3(GND_net), .O(n60762));
    defparam i1_2_lut_3_lut_adj_1751.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_4_lut_adj_1752 (.I0(\data_out_frame[15] [1]), .I1(n60531), 
            .I2(\data_out_frame[17] [2]), .I3(n29117), .O(n55796));
    defparam i2_3_lut_4_lut_adj_1752.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1753 (.I0(\data_out_frame[16] [3]), .I1(n62023), 
            .I2(\data_out_frame[21] [1]), .I3(n55781), .O(n8_adj_5426));
    defparam i1_2_lut_4_lut_adj_1753.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1754 (.I0(n60150), .I1(n60627), .I2(n60414), 
            .I3(n55802), .O(n62281));
    defparam i2_3_lut_4_lut_adj_1754.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1755 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [4]), 
            .I2(n28483), .I3(GND_net), .O(n55802));
    defparam i1_2_lut_3_lut_adj_1755.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i22686_2_lut (.I0(\FRAME_MATCHER.i[1] ), .I1(\FRAME_MATCHER.i[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n40778));
    defparam i22686_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1756 (.I0(n61010), .I1(\FRAME_MATCHER.i [3]), .I2(reset), 
            .I3(n9_adj_5705), .O(n59771));   // verilog/coms.v(157[7:23])
    defparam i3_4_lut_adj_1756.LUT_INIT = 16'hfff7;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51766 (.I0(byte_transmit_counter[1]), 
            .I1(n64848), .I2(n64849), .I3(byte_transmit_counter[4]), .O(n71247));
    defparam byte_transmit_counter_1__bdd_4_lut_51766.LUT_INIT = 16'he4aa;
    SB_LUT4 n71247_bdd_4_lut (.I0(n71247), .I1(n64624), .I2(n64623), .I3(byte_transmit_counter[4]), 
            .O(n71250));
    defparam n71247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51743 (.I0(byte_transmit_counter[1]), 
            .I1(n64893), .I2(n64894), .I3(byte_transmit_counter[2]), .O(n71241));
    defparam byte_transmit_counter_1__bdd_4_lut_51743.LUT_INIT = 16'he4aa;
    SB_LUT4 n71241_bdd_4_lut (.I0(n71241), .I1(n64597), .I2(n64596), .I3(byte_transmit_counter[2]), 
            .O(n71244));
    defparam n71241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51738 (.I0(byte_transmit_counter[1]), 
            .I1(n64896), .I2(n64897), .I3(byte_transmit_counter[2]), .O(n71235));
    defparam byte_transmit_counter_1__bdd_4_lut_51738.LUT_INIT = 16'he4aa;
    SB_LUT4 n71235_bdd_4_lut (.I0(n71235), .I1(n64900), .I2(n64899), .I3(byte_transmit_counter[2]), 
            .O(n71238));
    defparam n71235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(Kp_23__N_1748), .I1(n41), .I2(reset), 
            .I3(GND_net), .O(n25151));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_787_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1757 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5705));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1757.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1758 (.I0(n3489), .I1(n8_c), .I2(GND_net), .I3(GND_net), 
            .O(n60135));
    defparam i1_2_lut_adj_1758.LUT_INIT = 16'hdddd;
    SB_LUT4 i41580_4_lut (.I0(reset), .I1(n10_adj_5670), .I2(n60135), 
            .I3(n161), .O(n30673));
    defparam i41580_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1759 (.I0(n55179), .I1(n60441), .I2(\data_out_frame[21] [7]), 
            .I3(n60854), .O(n60265));
    defparam i2_3_lut_4_lut_adj_1759.LUT_INIT = 16'h6996;
    SB_LUT4 i45296_3_lut_4_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[1]), 
            .I2(n64862), .I3(n64860), .O(n64791));
    defparam i45296_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_4_lut_adj_1760 (.I0(n55179), .I1(n60441), .I2(n55796), 
            .I3(\data_out_frame[23] [4]), .O(n60764));
    defparam i2_3_lut_4_lut_adj_1760.LUT_INIT = 16'h6996;
    SB_LUT4 i21052_3_lut_4_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[1]), 
            .I2(n64844), .I3(n64842), .O(n39176));
    defparam i21052_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_787_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n61840), .I2(n60685), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5414));
    defparam select_787_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h6900;
    SB_LUT4 select_787_Select_213_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n61840), .I2(n60514), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5413));
    defparam select_787_Select_213_i3_3_lut_4_lut.LUT_INIT = 16'h9600;
    SB_LUT4 i11_4_lut_4_lut_adj_1761 (.I0(n30637), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[6]_c [4]), .O(n59373));
    defparam i11_4_lut_4_lut_adj_1761.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_211_i3_3_lut_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\data_out_frame[24] [2]), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n60682), .O(n3_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_211_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i13761_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n31952));
    defparam i13761_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13764_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n31955));
    defparam i13764_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13768_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n31959));
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13771_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n31962));
    defparam i13771_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13775_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n31966));
    defparam i13775_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1762 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\data_out_frame[0][2] ), .I3(GND_net), .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1762.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13778_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n31969));
    defparam i13778_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13782_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n31973));
    defparam i13782_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13785_3_lut_4_lut (.I0(n41173), .I1(n60130), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n31976));
    defparam i13785_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51733 (.I0(byte_transmit_counter[1]), 
            .I1(n64590), .I2(n64591), .I3(byte_transmit_counter[2]), .O(n71211));
    defparam byte_transmit_counter_1__bdd_4_lut_51733.LUT_INIT = 16'he4aa;
    SB_LUT4 n71211_bdd_4_lut (.I0(n71211), .I1(n64588), .I2(n64587), .I3(byte_transmit_counter[2]), 
            .O(n71214));
    defparam n71211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51715 (.I0(byte_transmit_counter[1]), 
            .I1(n64611), .I2(n64612), .I3(byte_transmit_counter[2]), .O(n71205));
    defparam byte_transmit_counter_1__bdd_4_lut_51715.LUT_INIT = 16'he4aa;
    SB_LUT4 n71205_bdd_4_lut (.I0(n71205), .I1(n64609), .I2(n64608), .I3(byte_transmit_counter[2]), 
            .O(n71208));
    defparam n71205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1763 (.I0(\data_in_frame[5] [6]), .I1(n28266), 
            .I2(\data_in_frame[1] [4]), .I3(n60262), .O(n28761));   // verilog/coms.v(18[27:29])
    defparam i2_3_lut_4_lut_adj_1763.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51710 (.I0(byte_transmit_counter[1]), 
            .I1(n64836), .I2(n64837), .I3(byte_transmit_counter[2]), .O(n71199));
    defparam byte_transmit_counter_1__bdd_4_lut_51710.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1764 (.I0(\data_in_frame[5] [6]), .I1(n28266), 
            .I2(n60848), .I3(GND_net), .O(n60271));   // verilog/coms.v(18[27:29])
    defparam i1_2_lut_3_lut_adj_1764.LUT_INIT = 16'h9696;
    SB_LUT4 n71199_bdd_4_lut (.I0(n71199), .I1(n64618), .I2(n64617), .I3(byte_transmit_counter[2]), 
            .O(n71202));
    defparam n71199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1765 (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[1]_c [1]), 
            .I2(\data_in_frame[3][3] ), .I3(\data_in_frame[0] [7]), .O(n28702));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1765.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1766 (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n60197), .I3(n60241), .O(Kp_23__N_767));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1766.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1767 (.I0(n28690), .I1(n70932), .I2(Kp_23__N_748), 
            .I3(GND_net), .O(n64267));
    defparam i1_2_lut_3_lut_adj_1767.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1768 (.I0(n28690), .I1(n70932), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n54762));
    defparam i1_2_lut_3_lut_adj_1768.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1769 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n28690));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1769.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1770 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n4_adj_5606));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1770.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1771 (.I0(\data_out_frame[18] [4]), .I1(n55273), 
            .I2(n60482), .I3(n54876), .O(n55267));
    defparam i1_2_lut_3_lut_4_lut_adj_1771.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1772 (.I0(\data_in_frame[6]_c [4]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[6] [7]), .I3(n60821), .O(n64085));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1772.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1773 (.I0(\data_in_frame[6]_c [4]), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_872), .I3(GND_net), .O(n60308));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1773.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_4_lut_adj_1774 (.I0(n30637), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[6]_c [5]), .O(n59379));
    defparam i11_4_lut_4_lut_adj_1774.LUT_INIT = 16'hfe10;
    SB_LUT4 i13904_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n32095));
    defparam i13904_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(n28031), .I3(\data_out_frame[5] [7]), .O(n60867));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_51705 (.I0(byte_transmit_counter[1]), 
            .I1(n64584), .I2(n64585), .I3(byte_transmit_counter[2]), .O(n71193));
    defparam byte_transmit_counter_1__bdd_4_lut_51705.LUT_INIT = 16'he4aa;
    SB_LUT4 i13907_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n32098));
    defparam i13907_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13910_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n32101));
    defparam i13910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n71193_bdd_4_lut (.I0(n71193), .I1(n64582), .I2(n64581), .I3(byte_transmit_counter[2]), 
            .O(n71196));
    defparam n71193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13913_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n32104));
    defparam i13913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13919_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n32110));
    defparam i13919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [0]), 
            .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'ha088;
    SB_LUT4 i13755_3_lut_4_lut (.I0(n30637), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[6][6] ), .O(n31946));
    defparam i13755_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13924_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n32115));
    defparam i13924_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13927_3_lut_4_lut (.I0(n8_c), .I1(n59771), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n32118));
    defparam i13927_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1776 (.I0(\data_in_frame[4] [4]), .I1(n70932), 
            .I2(n28715), .I3(\data_in_frame[6] [7]), .O(n60772));
    defparam i1_2_lut_3_lut_4_lut_adj_1776.LUT_INIT = 16'h9669;
    uart_tx tx (.n1(n1), .tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data[7:1], 
            \tx_data[0] }), .r_SM_Main({r_SM_Main}), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n59789(n59789), .GND_net(GND_net), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n63279(n63279), .n27(n27), .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), 
            .r_Clock_Count({r_Clock_Count}), .VCC_net(VCC_net), .n32272(n32272), 
            .n71737(n71737), .n30087(n30087), .n31705(n31705), .tx_active(tx_active), 
            .n5233(n5233), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), .n29(n29), .n23(n23), 
            .n61776(n61776), .n6(n6_adj_9), .n60925(n60925), .n63255(n63255), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.baudrate({baudrate}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n27889(n27889), .r_SM_Main({r_SM_Main_adj_23}), .clk16MHz(clk16MHz), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29(n29), .n23(n23), .r_Clock_Count({r_Clock_Count_adj_24}), 
            .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), 
            .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), 
            .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), 
            .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), 
            .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_21 ), 
            .n59798(n59798), .n63269(n63269), .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), 
            .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), .n5230(n5230), .n32278(n32278), 
            .n55993(n55993), .rx_data_ready(rx_data_ready), .n30084(n30084), 
            .n32606(n32606), .rx_data({rx_data}), .n32605(n32605), .n32604(n32604), 
            .n32603(n32603), .n32600(n32600), .n32599(n32599), .n32598(n32598), 
            .n32286(n32286), .n60086(n60086), .n4(n4), .n6(n6_adj_22), 
            .n30080(n30080), .n60927(n60927), .n63257(n63257), .n63621(n63621), 
            .n63605(n63605), .n63549(n63549), .n63515(n63515), .n63551(n63551), 
            .n63641(n63641), .n63587(n63587), .n63623(n63623)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n1, tx_o, clk16MHz, tx_data, r_SM_Main, \r_Bit_Index[0] , 
            n59789, GND_net, \r_SM_Main_2__N_3545[0] , n63279, n27, 
            \r_SM_Main_2__N_3536[1] , r_Clock_Count, VCC_net, n32272, 
            n71737, n30087, n31705, tx_active, n5233, \o_Rx_DV_N_3488[12] , 
            \o_Rx_DV_N_3488[24] , n29, n23, n61776, n6, n60925, 
            n63255, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output n1;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output n59789;
    input GND_net;
    input \r_SM_Main_2__N_3545[0] ;
    input n63279;
    input n27;
    input \r_SM_Main_2__N_3536[1] ;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n32272;
    input n71737;
    output n30087;
    input n31705;
    output tx_active;
    input n5233;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n29;
    input n23;
    input n61776;
    output n6;
    output n60925;
    output n63255;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n3, n27401;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n24197;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n24196;
    wire [8:0]n41;
    
    wire n53680, n53679, n53678, n53677, n61072, n53676, n53675, 
        n53674, n53673, o_Tx_Serial_N_3598, n3_adj_5315, n31418;
    wire [2:0]n460;
    
    wire n31396, n64845, n64846, n64606, n64605, n67691, n67688, 
        n63247, n63253, n71325;
    
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n24197), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59789));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6339_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n63279), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n24196));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i6339_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i6340_3_lut (.I0(n24196), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n24197));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i6340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2056_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n53680), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2056_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n53679), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_9 (.CI(n53679), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n53680));
    SB_LUT4 r_Clock_Count_2056_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n53678), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_8 (.CI(n53678), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n53679));
    SB_LUT4 r_Clock_Count_2056_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n53677), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i41625_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n61072));
    defparam i41625_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY r_Clock_Count_2056_add_4_7 (.CI(n53677), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n53678));
    SB_LUT4 r_Clock_Count_2056_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n53676), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_6 (.CI(n53676), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n53677));
    SB_LUT4 r_Clock_Count_2056_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n53675), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_5 (.CI(n53675), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n53676));
    SB_LUT4 r_Clock_Count_2056_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n53674), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_4 (.CI(n53674), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n53675));
    SB_LUT4 r_Clock_Count_2056_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n53673), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_3 (.CI(n53673), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n53674));
    SB_LUT4 r_Clock_Count_2056_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n53673));
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3598), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5315), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n27401), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_2056__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n31418));   // verilog/uart_tx.v(119[34:51])
    SB_LUT4 i51604_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3536[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n31418));
    defparam i51604_4_lut.LUT_INIT = 16'h1115;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n32272));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n71737));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n30087), 
            .D(n460[1]), .R(n31396));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n30087), 
            .D(n460[2]), .R(n31396));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n31705));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i45350_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64845));
    defparam i45350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45351_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64846));
    defparam i45351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45111_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64606));
    defparam i45111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45110_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n64605));
    defparam i45110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49174_3_lut (.I0(n5233), .I1(\o_Rx_DV_N_3488[12] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n67691));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49174_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i49171_4_lut (.I0(n67691), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67688));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i49171_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n67688), .I1(n61776), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5315));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n61776), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i2336_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2336_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5233), .I2(n59789), 
            .I3(GND_net), .O(n63247));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), .I3(n63247), 
            .O(n63253));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n63253), .I1(n61072), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n31396));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h0323;
    SB_LUT4 i2329_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2329_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i41486_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n60925));
    defparam i41486_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(n59789), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n63255));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i51694_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n30087));
    defparam i51694_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n64605), 
            .I2(n64606), .I3(r_Bit_Index[2]), .O(n71325));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71325_bdd_4_lut (.I0(n71325), .I1(n64846), .I2(n64845), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3598));
    defparam n71325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n27401));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (baudrate, GND_net, VCC_net, n27889, r_SM_Main, clk16MHz, 
            r_Rx_Data, RX_N_2, \o_Rx_DV_N_3488[24] , n27, n29, n23, 
            r_Clock_Count, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \r_Bit_Index[0] , n59798, n63269, \r_SM_Main_2__N_3446[1] , 
            \o_Rx_DV_N_3488[0] , n5230, n32278, n55993, rx_data_ready, 
            n30084, n32606, rx_data, n32605, n32604, n32603, n32600, 
            n32599, n32598, n32286, n60086, n4, n6, n30080, n60927, 
            n63257, n63621, n63605, n63549, n63515, n63551, n63641, 
            n63587, n63623) /* synthesis syn_module_defined=1 */ ;
    input [31:0]baudrate;
    input GND_net;
    input VCC_net;
    output n27889;
    output [2:0]r_SM_Main;
    input clk16MHz;
    output r_Rx_Data;
    input RX_N_2;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n29;
    output n23;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0] ;
    output n59798;
    input n63269;
    input \r_SM_Main_2__N_3446[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n5230;
    input n32278;
    input n55993;
    output rx_data_ready;
    output n30084;
    input n32606;
    output [7:0]rx_data;
    input n32605;
    input n32604;
    input n32603;
    input n32600;
    input n32599;
    input n32598;
    input n32286;
    input n60086;
    output n4;
    output n6;
    output n30080;
    output n60927;
    output n63257;
    input n63621;
    output n63605;
    input n63549;
    output n63515;
    output n63551;
    output n63641;
    output n63587;
    output n63623;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n70771, n2597, n70772, n42, n960, n70404, n21, n19, 
        n17, n9, n68090, n43, n16, n67997, n69176, n70228, n43_adj_5043, 
        n69496, n70478, n959, n70405, n8, n70481, n37, n69174, 
        n2599;
    wire [23:0]n8189;
    wire [23:0]n294;
    
    wire n2716, n45, n24, n3172;
    wire [23:0]n8319;
    
    wire n3274, n7, n68124;
    wire [23:0]n8241;
    
    wire n2845, n858, n53406, n13, n11, n69096, n15, n69090, 
        n53407, n25, n23_c, n70482, n60967, n48, n31, n29_c, 
        n27_c, n69818, n63911, n27999, n63953, n63909, n27951, 
        n63151, n538, n61262, n37_adj_5044, n35, n33, n70700, 
        n64527, n64477, n60980, n64561, n64517, n64383, n64385, 
        n64567, n41, n1602, n12, n2488;
    wire [23:0]n8163;
    
    wire n2608;
    wire [23:0]n8215;
    
    wire n2713, n2977, n53405, n2725, n2714, n63157, n48_adj_5045, 
        n4_c, n70382, n2867, n53404, n70383, n68036, n10, n30, 
        n2715, n2754, n53403, n68055, n68042, n70747, n2638, n53402, 
        n1116, n70249, n70893, n70894, n1742, n6_c;
    wire [23:0]n7903;
    
    wire n1266, n70384, n2609, n2726, n64323, n48_adj_5046;
    wire [23:0]n7929;
    
    wire n1413;
    wire [23:0]n7955;
    
    wire n1557, n70385, n68007, n1879, n2717, n2519, n53401, n69860, 
        n70247, n39, n70829, n41_adj_5047, n68009, n63703, n64467, 
        n70530;
    wire [23:0]n7981;
    
    wire n1698, n40, n63119;
    wire [23:0]n8007;
    
    wire n1836, n45_adj_5048, n69846, n1408, n63137, n1560, n3151, 
        n3253, n21_adj_5049, n70532, n64063, n63925, n63921, n63127, 
        n62087, n23_adj_5050, n2600, n2724, n25_adj_5051, n64529;
    wire [23:0]n8033;
    
    wire n1971, n3050;
    wire [23:0]n8293;
    
    wire n3155, n3053, n3158, n33_adj_5052, n64533, n48_adj_5053, 
        n3054, n3159;
    wire [23:0]n8059;
    
    wire n2103, n31_adj_5054, n2718, n37_adj_5055, n3051, n3156, 
        n37_adj_5056, n63973, n63897, n63899, n1414, n67826, n37_adj_5057, 
        n3052, n3157, n36, n68454, n39_adj_5058, n35_adj_5059, n2598, 
        n3059, n3164, n64397, n63845, n64539, n3058, n3163, n21_adj_5060, 
        n19_adj_5061, n17_adj_5062, n2729, n69482, n63713, n40931, 
        n63107, n27987, n62097, n23_adj_5063, n3065, n3170, n69998, 
        n3066, n3171, n9_adj_5064, n3056, n3161, n40933, n63419, 
        n3057, n3162, n43_adj_5065, n25_adj_5066, n27_adj_5067, n63437, 
        n64487, n64479, n64559, n3064, n3169, n11_adj_5068, n3060, 
        n3165, n61773, n19_adj_5069, n3061, n3166, n3062, n3167, 
        n3055, n3160, n3063, n3168, n13_adj_5070, n31_adj_5071, 
        n29_adj_5072, n27_adj_5073, n69994, n15_adj_5074, n17_adj_5075, 
        n27896, n29_adj_5076, n64067, n63705, n63701, n63723, n2397, 
        n53400, n63709, n63711, n63707, n63725, n2013, n27990, 
        n2602, n2719, n48_adj_5077, n64069, n64065, n28002, n68167, 
        n2603, n2720, n35_adj_5078, n33_adj_5079, n68456, n69234, 
        n69864, n69862, n2272, n53399, n68169, n6_adj_5080, n70390, 
        n63767, n3, n2144, n53398, n14, n32, n70391, r_Rx_Data_R, 
        n68161, n2730, n14_adj_5081, n12_adj_5082, n68156, n70745, 
        n67592, n70239, n63841, n67593, n70159, n60961, n8_adj_5083, 
        n70392, n70160, n70393, n52857, n68186, n69221, n10_adj_5084, 
        n69858, n2721, n53397, n70237, n2604, n2605, n2722, n70213, 
        n52856, n63131, n2606, n2723, n70891, n53396, n53395, 
        n2610, n2727, n2611, n2728, n53394, n70386, n52855, n63187, 
        n2612, n70911, n70912, n1459, n53393, n1460, n53392, n2607, 
        n3154, n70906, n60965, n3153, n70678, n2476, n2596, n1011, 
        n53391, n2477, n3152, n70679, n2481, n2601, n52854;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n2478, n856, n53390;
    wire [7:0]n1;
    
    wire n53641, n53640, n53639, n3084, n2479, n53638, n53637, 
        n3049, n22, n40_adj_5092, n53636, n68439, n53635, n52853, 
        n63185, n698, n53389, n52852, n63183, n3188, n41_adj_5095, 
        n3048, n2480, n803, n9625, n24106, n46, n20, n68431, 
        n70230, n39_adj_5096, n52851, n53388, n52850, n63181, n2482, 
        n69188, n2484, n2483, n31_adj_5097, n52849, n63179, n33_adj_5098, 
        n35_adj_5099, n2485, n2486, n27_adj_5100, n29_adj_5101, n63149, 
        n61266, n9796, n24124, n46_adj_5102, n2490, n1111, n2489, 
        n19_adj_5103, n21_adj_5104, n52848, n63129, n2491, n18, 
        n26, n2363;
    wire [23:0]n8137;
    
    wire n52847, n63177, n16_adj_5105, n68473, n70652, n53387, n2353, 
        n52846, n53386, n52845, n53385, n2357, n61270, n52844, 
        n39_adj_5106, n53384, n52843, n2354, n53383, n52842, n45_adj_5107, 
        n2355, n53382, n53381, n43_adj_5108, n53380, n70653, n70473, 
        n70336, n70708, n69186, n70710, n63143, n48_adj_5109, n53379, 
        n1261, n2356, n41_adj_5110, n2358, n2360, n2359, n33_adj_5111, 
        n1552, n35_adj_5112, n63861, n3_adj_5113, n37_adj_5114, n63865, 
        n5, n63869, n1693, n2365, n8_adj_5115, n2366, n59836, 
        n21_adj_5116;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n23_adj_5117, n1831, n2362, n2361, n1966, n29_adj_5118, 
        n31_adj_5119, n64439, n2098, n2101, n41_adj_5120, n2367, 
        n64545, n2487, n25_adj_5121, n2, n63975, n27_adj_5122, n10012, 
        n63923, n63961, n63983, n63979, n63981, n27975, n19_adj_5123, 
        n68612, n2108, n27_adj_5124, n68600, n70360, n33_adj_5125, 
        n31_adj_5126, n29_adj_5127, n68725, n18_adj_5128, n70171, 
        n70172, n30_adj_5129, n38_adj_5130, n61285, n68606, n69554, 
        n24_adj_5131, n26_adj_5132, n2109, n26_adj_5133, n69170, n53378, 
        n53377, n53376, n53375, n53374, n53373, n53372, n53371, 
        n22_adj_5134, n30_adj_5135, n63147, n53370, n53369, n20_adj_5136, 
        n68596, n70646, n53368, n70647, n52841, n53367, n53366, 
        n53365, n53364, n70185, n70485, n53363, n69560, n53362, 
        n53361, n53360, n70225, n53359, n53358, n53357, n53356, 
        n53355, n63145, n61274, n53354, n53353, n53352, n69168, 
        n53351, n53350, n53349, n53348, n70227, n53347, n53346, 
        n53345, n53344, n2364, n53343, n53342, n53341, n53340, 
        n61278;
    wire [23:0]n8111;
    
    wire n2227, n53339, n2228, n53338, n2229, n53337, n2230, n53336, 
        n2231, n53335, n2232, n53334, n52840, n2233, n53333, n3186, 
        n53488, n2234, n53332, n2235, n53331, n2236, n53330, n2237, 
        n53329, n3082, n53487, n35_adj_5137, n70186, n2238, n53328, 
        n2239, n53327, n2240, n53326, n63141, n61282;
    wire [23:0]n8085;
    
    wire n53325, n2099, n53324, n2100, n53323, n53322, n2102, 
        n53321, n53320, n2104, n53319, n2105, n53318, n2106, n53317, 
        n2107, n53316, n53315, n53314, n2110, n53313, n1967, n53312, 
        n1968, n53311, n1969, n53310, n1970, n53309, n53308, n1972, 
        n53307, n1973, n53306, n30202, n31416, n3_adj_5138, n1974, 
        n53305, n52839, n1975, n53304, n1976, n53303, n52838, 
        n1977, n53302, n53301, n1832, n53300, n1833, n53299, n52837, 
        n39_adj_5139, n68709, n28, n68706, n70640, n41_adj_5140, 
        n52836, n1834, n53298, n1835, n53297, n53486, n53296, 
        n52835, n1837, n53295, n53485, n1838, n53294, n52834, 
        n1839, n53293, n1840, n53292, n53484, n1841, n53291, n63139, 
        n61291, n53483, n39_adj_5141, n53482, n69148, n37_adj_5142, 
        n70840, n53481, n53480, n53280, n1694, n53279, n70841, 
        n70774, n1695, n53278, n1696, n53277, n53479, n1697, n53276, 
        n53478, n35_adj_5143, n53275, n53477, n1699, n53274, n1700, 
        n53273, n1701, n53272, n53476, n53475, n1702, n53474, 
        n53473, n53271, n1553, n53270, n48_adj_5144, n1554, n53269, 
        n53472, n53471, n1555, n53268, n53470, n1556, n53267, 
        n67678, n67684, n53469, n53468, n67675, n53467, n53466, 
        n61250, n67681, n53266, n3046, n53465, n31_adj_5145, n3047, 
        n53464, n1558, n53265, n33_adj_5146, n53463, n1559, n53264, 
        n25_adj_5147, n27_adj_5148, n29_adj_5149, n53462, n53461, 
        n37_adj_5150, n29_adj_5151, n35_adj_5152, n31_adj_5153, n41_adj_5154, 
        n53460, n39_adj_5155, n29_adj_5156, n23_adj_5157, n31_adj_5158, 
        n33_adj_5159, n53263, n53459, n27_adj_5160, n68690, n68769, 
        n35_adj_5161, n33_adj_5162, n68680, n53262, n67631, n1409, 
        n53261, n53458, n30_adj_5163, n38_adj_5164, n22_adj_5165, 
        n26_adj_5166, n1410, n53260, n67628, n1411, n53259, n67625, 
        n28_adj_5167, n30_adj_5168, n70193, n70194, n1412, n53258, 
        n68753, n28_adj_5169, n68742, n70636, n69140, n53457, n26_adj_5170, 
        n37_adj_5171, n34, n53257, n70838, n24_adj_5172, n68674, 
        n70642, n39_adj_5173, n70643, n70839, n70776, n48_adj_5174, 
        n53256, n1415, n53255, n63211, n61300, n41_adj_5175, n70489, 
        n70368, n45_adj_5176, n39_adj_5177, n63217, n53254, n1262, 
        n53253, n68682, n70398, n43_adj_5178, n69158, n43_adj_5179, 
        n41_adj_5180, n1263, n53252, n1264, n53251, n1265, n53250, 
        n53249, n70630, n70631, n34_adj_5181, n1267, n53248, n70400, 
        n70401, n68845, n38_adj_5182, n63135, n61304, n53247, n23_adj_5183, 
        n44_adj_5184, n25_adj_5185, n27_adj_5186, n1112, n53246, n21_adj_5187, 
        n68641, n1113, n53245, n1114, n53244, n1115, n53243, n53242, 
        n63133, n61308, n53456, n53455, n53454, n53453, n53452, 
        n53451, n53450, n53449, n53448, n53447, n70910, n2938, 
        n63153, n53446, n70898, n2827, n2957, n68632, n27993, 
        n962, n53445;
    wire [2:0]n479;
    
    wire n31398, n63155, n61254;
    wire [23:0]n8267;
    
    wire n53444, n2939, n53443, n2940, n53442, n71751, n2941, 
        n53441, n2942, n53440, n2943, n53439, n26_adj_5188, n28_adj_5189, 
        n2944, n53438, n2945, n53437, n2946, n53436, n2947, n53435, 
        n2948, n53434, n2949, n53433, n2950, n53432, n2951, n53431, 
        n2952, n53430, n2953, n53429, n2954, n53428, n2955, n53427, 
        n2956, n53426, n53425, n61258, n53424, n2828, n53423, 
        n2829, n53422, n2830, n53421, n2831, n53420, n2832, n53419, 
        n2833, n53418, n2834, n53417, n2835, n53416, n2836, n53415, 
        n2837, n53414, n2838, n53413, n2839, n53412, n2840, n53411, 
        n2841, n53410, n41_adj_5190, n36_adj_5191, n38_adj_5192, n40_adj_5193, 
        n67837, n70741, n70742, n63965, n63873, n63697, n2842, 
        n53409, n63967, n2843, n53408, n70635, n2844, n43_adj_5194, 
        n33_adj_5195, n31_adj_5196, n39_adj_5197, n41_adj_5198, n37_adj_5199, 
        n63971, n43_adj_5200, n24_adj_5201, n32_adj_5202, n39_adj_5203, 
        n41_adj_5204, n38_adj_5205, n40_adj_5206, n42_adj_5207, n67845, 
        n70508, n70509, n22_adj_5208, n68630, n70644, n70645, n35_adj_5209, 
        n37_adj_5210, n70487, n29_adj_5211, n70362, n68793, n14_adj_5212, 
        n15_adj_5213, n20_adj_5214, n68635, n70743, n32_adj_5215, 
        n40_adj_5216, n28_adj_5217, n64461, n64459, n63919, n70195, 
        n70196, n69162, n70836, n70837, n68786, n30_adj_5218, n68784, 
        n70632, n69136, n70780, n70834, n70835, n12_adj_5219, n68351, 
        n14_adj_5220, n16_adj_5221, n68316, n18_adj_5222, n9789, n40_adj_5223, 
        n14_adj_5224, n68411, n16_adj_5225, n24096, n42_adj_5226, 
        n18_adj_5227, n68381, n20_adj_5228, n67662, n63941, n63883, 
        n24122, n44_adj_5229, n804, n44_adj_5230, n44_adj_5231, n68038, 
        n10_adj_5232, n14_adj_5233, n68241, n805, n16_adj_5234, n12_adj_5235, 
        n68286, n18_adj_5237, n68543, n20_adj_5238, n22_adj_5239, 
        n64503, n43_adj_5240, n37_adj_5241, n39_adj_5242, n41_adj_5243, 
        n32_adj_5244, n70199, n23_adj_5245, n70200, n67815, n68832, 
        n68555, n63237, n63243, n34_adj_5246, n70215, n63057, n25_adj_5248, 
        n67620, n67617, n69130, n70502, n70503, n70523, n63969, 
        n48_adj_5249, n64531, n35_adj_5250, n39_adj_5251, n33_adj_5252, 
        n43_adj_5253, n37_adj_5254, n63055, n17_adj_5255, n61294, 
        n68557, n27_adj_5256, n29_adj_5257, n68549, n70350, n32_adj_5258, 
        n16_adj_5259, n70197, n70165, n70198, n68817, n69706, n34_adj_5260, 
        n70217, n69133, n23_adj_5261, n70500, n70501, n25_adj_5262, 
        n70166, n48_adj_5263, n21_adj_5264, n63951, n27966, n28_adj_5265, 
        n70648, n70649, n15_adj_5266, n17_adj_5267, n19_adj_5268, 
        n31_adj_5269, n69504, n961, n11_adj_5270, n13_adj_5271, n68252, 
        n69310, n69908, n69902, n68254, n8_adj_5272, n70131, n70132, 
        n34_adj_5273, n63475, n68243, n70668, n69214, n64481, n70133, 
        n70134, n69284, n20_adj_5274, n69212, n70272, n70846, n69856, 
        n70915, n63503, n70916, n70908, n64557, n37_adj_5275, n70934, 
        n41_adj_5276, n35_adj_5277, n39_adj_5278, n29_adj_5279, n31_adj_5280, 
        n23_adj_5281, n25_adj_5282, n27_adj_5283, n17_adj_5284, n19_adj_5285, 
        n21_adj_5286, n33_adj_5287, n39_adj_5288, n37_adj_5289, n43_adj_5290, 
        n41_adj_5291, n25_adj_5292, n27_adj_5293, n29_adj_5294, n15_adj_5295, 
        n17_adj_5296, n19_adj_5297, n21_adj_5298, n23_adj_5299, n31_adj_5300, 
        n63819, n33_adj_5301, n35_adj_5302, n68397, n69426, n69974, 
        n69972, n68401, n12_adj_5303, n46_adj_5304, n48_adj_5305, 
        n63901, n63903, n63853, n70153, n27945, n38_adj_5306, n70154, 
        n68044, n68385, n42_adj_5307, n70504, n70626, n70505, n69196, 
        n24_adj_5308, n70654, n70655, n70471, n70328, n70832, n69194, 
        n70897, n13_adj_5309, n15_adj_5310, n68331, n69370, n69946, 
        n69942, n68335, n10_adj_5311, n70147, n70148, n42_adj_5312, 
        n36_adj_5313, n68318, n70664, n69202, n22_adj_5314, n70656, 
        n70657, n70469, n70316, n70844, n69200, n70913, n70914, 
        n61311;
    
    SB_LUT4 i51277_3_lut (.I0(n70771), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n70772));   // verilog/uart_rx.v(119[33:55])
    defparam i51277_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50909_3_lut (.I0(n42), .I1(baudrate[3]), .I2(n960), .I3(GND_net), 
            .O(n70404));   // verilog/uart_rx.v(119[33:55])
    defparam i50909_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48595_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n68090));
    defparam i48595_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48502_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n67997));
    defparam i48502_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50983_4_lut (.I0(n69176), .I1(n70228), .I2(n43_adj_5043), 
            .I3(n69496), .O(n70478));   // verilog/uart_rx.v(119[33:55])
    defparam i50983_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50910_3_lut (.I0(n70404), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n70405));   // verilog/uart_rx.v(119[33:55])
    defparam i50910_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49679_3_lut (.I0(n70481), .I1(baudrate[12]), .I2(n37), .I3(GND_net), 
            .O(n69174));   // verilog/uart_rx.v(119[33:55])
    defparam i49679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8189[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8319[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48629_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n68124));
    defparam i48629_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 add_2755_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n53406), 
            .O(n8241[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49601_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n68124), 
            .O(n69096));
    defparam i49601_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49595_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n69096), 
            .O(n69090));
    defparam i49595_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2755_3 (.CI(n53406), .I0(n2845), .I1(n858), .CO(n53407));
    SB_LUT4 i50987_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n69090), 
            .O(n70482));
    defparam i50987_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50711_3_lut (.I0(n70405), .I1(baudrate[5]), .I2(n60967), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i50711_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i50323_4_lut (.I0(n31), .I1(n29_c), .I2(n27_c), .I3(n70482), 
            .O(n69818));
    defparam i50323_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut (.I0(n63911), .I1(n27999), .I2(n63953), .I3(n63909), 
            .O(n27951));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2755_2_lut (.I0(n61262), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i51205_4_lut (.I0(n37_adj_5044), .I1(n35), .I2(n33), .I3(n69818), 
            .O(n70700));
    defparam i51205_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i45075_4_lut (.I0(n64527), .I1(n64477), .I2(n60980), .I3(baudrate[4]), 
            .O(n64561));
    defparam i45075_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51685_4_lut (.I0(n64517), .I1(n64383), .I2(n64561), .I3(n64385), 
            .O(n64567));
    defparam i51685_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2755_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53406));
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8163[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n53405), 
            .O(n8215[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8189[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8189[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63157), .I3(n48_adj_5045), .O(n4_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i50887_3_lut (.I0(n4_c), .I1(baudrate[13]), .I2(n27_c), .I3(GND_net), 
            .O(n70382));   // verilog/uart_rx.v(119[33:55])
    defparam i50887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n53404), 
            .O(n8215[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_19 (.CI(n53404), .I0(n2714), .I1(n2867), .CO(n53405));
    SB_LUT4 i50888_3_lut (.I0(n70382), .I1(baudrate[14]), .I2(n29_c), 
            .I3(GND_net), .O(n70383));   // verilog/uart_rx.v(119[33:55])
    defparam i50888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48541_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n68036));
    defparam i48541_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n53403), 
            .O(n8215[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_18 (.CI(n53403), .I0(n2715), .I1(n2754), .CO(n53404));
    SB_LUT4 i48547_4_lut (.I0(n33), .I1(n31), .I2(n29_c), .I3(n68055), 
            .O(n68042));
    defparam i48547_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51252_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n68036), 
            .O(n70747));   // verilog/uart_rx.v(119[33:55])
    defparam i51252_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2754_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n53402), 
            .O(n8215[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(n27951), .I1(n48), .I2(baudrate[0]), .I3(GND_net), 
            .O(n1116));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_CARRY add_2754_17 (.CI(n53402), .I0(n2716), .I1(n2638), .CO(n53403));
    SB_LUT4 i50754_3_lut (.I0(n70383), .I1(baudrate[15]), .I2(n31), .I3(GND_net), 
            .O(n70249));   // verilog/uart_rx.v(119[33:55])
    defparam i50754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51398_4_lut (.I0(n70249), .I1(n70747), .I2(n35), .I3(n68042), 
            .O(n70893));   // verilog/uart_rx.v(119[33:55])
    defparam i51398_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51399_3_lut (.I0(n70893), .I1(baudrate[18]), .I2(n37_adj_5044), 
            .I3(GND_net), .O(n70894));   // verilog/uart_rx.v(119[33:55])
    defparam i51399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7903[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50889_3_lut (.I0(n6_c), .I1(baudrate[10]), .I2(n21), .I3(GND_net), 
            .O(n70384));   // verilog/uart_rx.v(119[33:55])
    defparam i50889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8189[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51489_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n64323), .I2(n48_adj_5046), 
            .I3(baudrate[15]), .O(n294[9]));
    defparam i51489_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7929[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7955[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50890_3_lut (.I0(n70384), .I1(baudrate[11]), .I2(n23_c), 
            .I3(GND_net), .O(n70385));   // verilog/uart_rx.v(119[33:55])
    defparam i50890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48512_4_lut (.I0(n43), .I1(n25), .I2(n23_c), .I3(n68090), 
            .O(n68007));
    defparam i48512_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2754_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n53401), 
            .O(n8215[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50365_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n67997), 
            .O(n69860));   // verilog/uart_rx.v(119[33:55])
    defparam i50365_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50752_3_lut (.I0(n70385), .I1(baudrate[12]), .I2(n25), .I3(GND_net), 
            .O(n70247));   // verilog/uart_rx.v(119[33:55])
    defparam i50752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51334_3_lut (.I0(n70894), .I1(baudrate[19]), .I2(n39), .I3(GND_net), 
            .O(n70829));   // verilog/uart_rx.v(119[33:55])
    defparam i51334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48514_4_lut (.I0(n43), .I1(n41_adj_5047), .I2(n39), .I3(n70700), 
            .O(n68009));
    defparam i48514_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i44981_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n64323), .I2(n63703), 
            .I3(baudrate[15]), .O(n64467));
    defparam i44981_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51035_4_lut (.I0(n70247), .I1(n69860), .I2(n45), .I3(n68007), 
            .O(n70530));   // verilog/uart_rx.v(119[33:55])
    defparam i51035_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7981[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51296_3_lut (.I0(n70829), .I1(baudrate[20]), .I2(n41_adj_5047), 
            .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam i51296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63119));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8007[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(n69846), .I1(baudrate[8]), .I2(n1408), 
            .I3(n63137), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8319[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51037_4_lut (.I0(n40), .I1(n70530), .I2(n45), .I3(n68009), 
            .O(n70532));   // verilog/uart_rx.v(119[33:55])
    defparam i51037_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_989 (.I0(n64063), .I1(n63925), .I2(n63119), .I3(n63921), 
            .O(n63127));
    defparam i1_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i51607_4_lut (.I0(n63127), .I1(n70532), .I2(baudrate[23]), 
            .I3(n3253), .O(n62087));   // verilog/uart_rx.v(119[33:55])
    defparam i51607_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8189[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51477_2_lut_4_lut (.I0(n69846), .I1(baudrate[8]), .I2(n1408), 
            .I3(n64529), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i51477_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8033[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8293[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8293[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51451_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n64533), .I3(n48_adj_5053), .O(n294[19]));
    defparam i51451_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8293[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8059[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8293[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_990 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n63973));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_991 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n63897));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_992 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n63899));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'heeee;
    SB_LUT4 i48331_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n67826));   // verilog/uart_rx.v(119[33:55])
    defparam i48331_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8293[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48959_4_lut (.I0(n37_adj_5055), .I1(n25_adj_5051), .I2(n23_adj_5050), 
            .I3(n21_adj_5049), .O(n68454));
    defparam i48959_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i41534_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n60980));
    defparam i41534_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8189[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_16 (.CI(n53401), .I0(n2717), .I1(n2519), .CO(n53402));
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8293[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44911_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n64397));
    defparam i44911_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45053_4_lut (.I0(n64397), .I1(n63845), .I2(n63899), .I3(baudrate[9]), 
            .O(n64539));
    defparam i45053_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8293[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49987_4_lut (.I0(n19_adj_5061), .I1(n17_adj_5062), .I2(n2729), 
            .I3(baudrate[2]), .O(n69482));
    defparam i49987_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_4_lut_adj_993 (.I0(baudrate[17]), .I1(n63713), .I2(baudrate[2]), 
            .I3(n40931), .O(n63107));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_994 (.I0(n64517), .I1(n63107), .I2(n27987), .I3(n64477), 
            .O(n62097));
    defparam i1_4_lut_adj_994.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8293[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50503_4_lut (.I0(n25_adj_5051), .I1(n23_adj_5050), .I2(n21_adj_5049), 
            .I3(n69482), .O(n69998));
    defparam i50503_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8293[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8293[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_995 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n40933), .O(n63419));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8293[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_996 (.I0(n63419), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n63437));
    defparam i1_4_lut_adj_996.LUT_INIT = 16'h0002;
    SB_LUT4 i45073_4_lut (.I0(n64487), .I1(n64477), .I2(n64479), .I3(n64383), 
            .O(n64559));
    defparam i45073_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8293[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8293[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_997 (.I0(n64539), .I1(n64559), .I2(n60980), .I3(n63437), 
            .O(n61773));
    defparam i1_4_lut_adj_997.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8293[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8293[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8293[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8293[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50499_4_lut (.I0(n31_adj_5071), .I1(n29_adj_5072), .I2(n27_adj_5073), 
            .I3(n69998), .O(n69994));
    defparam i50499_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51577_3_lut (.I0(n27896), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n27889));   // verilog/uart_rx.v(119[33:55])
    defparam i51577_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n64067));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_999 (.I0(n63705), .I1(n63701), .I2(n63703), .I3(n64383), 
            .O(n63723));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2754_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n53400), 
            .O(n8215[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n64063));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(n63713), .I1(n63709), .I2(n63711), 
            .I3(n63707), .O(n63725));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1002 (.I0(n63725), .I1(n27990), .I2(n63723), 
            .I3(GND_net), .O(n27896));
    defparam i1_3_lut_adj_1002.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8189[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n61773), .I1(baudrate[2]), 
            .I2(n62097), .I3(GND_net), .O(n48_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1003 (.I0(n64067), .I1(n64069), .I2(n63921), 
            .I3(n64065), .O(n28002));
    defparam i1_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 i48672_4_lut (.I0(n29_adj_5076), .I1(n17_adj_5075), .I2(n15_adj_5074), 
            .I3(n13_adj_5070), .O(n68167));
    defparam i48672_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8189[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48961_4_lut (.I0(n37_adj_5055), .I1(n35_adj_5078), .I2(n33_adj_5079), 
            .I3(n69994), .O(n68456));
    defparam i48961_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49739_4_lut (.I0(n11_adj_5068), .I1(n9_adj_5064), .I2(n3171), 
            .I3(baudrate[2]), .O(n69234));
    defparam i49739_4_lut.LUT_INIT = 16'heffe;
    SB_CARRY add_2754_15 (.CI(n53400), .I0(n2718), .I1(n2397), .CO(n53401));
    SB_LUT4 i44838_2_lut (.I0(baudrate[17]), .I1(n27987), .I2(GND_net), 
            .I3(GND_net), .O(n64323));
    defparam i44838_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50369_4_lut (.I0(n17_adj_5075), .I1(n15_adj_5074), .I2(n13_adj_5070), 
            .I3(n69234), .O(n69864));
    defparam i50369_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51460_2_lut (.I0(n48_adj_5077), .I1(n27896), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i51460_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i50367_4_lut (.I0(n23_adj_5063), .I1(n21_adj_5060), .I2(n19_adj_5069), 
            .I3(n69864), .O(n69862));
    defparam i50367_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_2754_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n53399), 
            .O(n8215[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48674_4_lut (.I0(n29_adj_5076), .I1(n27_adj_5067), .I2(n25_adj_5066), 
            .I3(n69862), .O(n68169));
    defparam i48674_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50895_3_lut (.I0(n6_adj_5080), .I1(baudrate[13]), .I2(n29_adj_5076), 
            .I3(GND_net), .O(n70390));   // verilog/uart_rx.v(119[33:55])
    defparam i50895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(n63909), .I1(n63973), .I2(baudrate[16]), 
            .I3(n40931), .O(n63767));
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'h0100;
    SB_CARRY add_2754_14 (.CI(n53399), .I0(n2719), .I1(n2272), .CO(n53400));
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2754_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n53398), 
            .O(n8215[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14), .I1(baudrate[17]), 
            .I2(n37_adj_5057), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50896_3_lut (.I0(n70390), .I1(baudrate[14]), .I2(n31_adj_5054), 
            .I3(GND_net), .O(n70391));   // verilog/uart_rx.v(119[33:55])
    defparam i50896_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48666_4_lut (.I0(n35_adj_5059), .I1(n33_adj_5052), .I2(n31_adj_5054), 
            .I3(n68167), .O(n68161));
    defparam i48666_4_lut.LUT_INIT = 16'haaab;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51250_4_lut (.I0(n32), .I1(n12_adj_5082), .I2(n37_adj_5057), 
            .I3(n68156), .O(n70745));   // verilog/uart_rx.v(119[33:55])
    defparam i51250_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49336_3_lut (.I0(n61773), .I1(n62097), .I2(baudrate[2]), 
            .I3(GND_net), .O(n67592));   // verilog/uart_rx.v(119[33:55])
    defparam i49336_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i50744_3_lut (.I0(n70391), .I1(baudrate[15]), .I2(n33_adj_5052), 
            .I3(GND_net), .O(n70239));   // verilog/uart_rx.v(119[33:55])
    defparam i50744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49159_4_lut (.I0(n60980), .I1(n63767), .I2(n63911), .I3(n63841), 
            .O(n67593));   // verilog/uart_rx.v(119[33:55])
    defparam i49159_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i50664_3_lut (.I0(n14_adj_5081), .I1(baudrate[13]), .I2(n37_adj_5055), 
            .I3(GND_net), .O(n70159));   // verilog/uart_rx.v(119[33:55])
    defparam i50664_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_13 (.CI(n53398), .I0(n2720), .I1(n2144), .CO(n53399));
    SB_LUT4 div_37_i427_4_lut (.I0(n67593), .I1(n67592), .I2(n294[21]), 
            .I3(n64323), .O(n60961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i50897_3_lut (.I0(n8_adj_5083), .I1(baudrate[10]), .I2(n23_adj_5063), 
            .I3(GND_net), .O(n70392));   // verilog/uart_rx.v(119[33:55])
    defparam i50897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50665_3_lut (.I0(n70159), .I1(baudrate[14]), .I2(n39_adj_5058), 
            .I3(GND_net), .O(n70160));   // verilog/uart_rx.v(119[33:55])
    defparam i50665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50898_3_lut (.I0(n70392), .I1(baudrate[11]), .I2(n25_adj_5066), 
            .I3(GND_net), .O(n70393));   // verilog/uart_rx.v(119[33:55])
    defparam i50898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n52857), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49726_4_lut (.I0(n25_adj_5066), .I1(n23_adj_5063), .I2(n21_adj_5060), 
            .I3(n68186), .O(n69221));
    defparam i49726_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50363_3_lut (.I0(n10_adj_5084), .I1(baudrate[9]), .I2(n21_adj_5060), 
            .I3(GND_net), .O(n69858));   // verilog/uart_rx.v(119[33:55])
    defparam i50363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n53397), 
            .O(n8215[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_12 (.CI(n53397), .I0(n2721), .I1(n2013), .CO(n53398));
    SB_LUT4 i50742_3_lut (.I0(n70393), .I1(baudrate[12]), .I2(n27_adj_5067), 
            .I3(GND_net), .O(n70237));   // verilog/uart_rx.v(119[33:55])
    defparam i50742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8189[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8189[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50718_4_lut (.I0(n35_adj_5059), .I1(n33_adj_5052), .I2(n31_adj_5054), 
            .I3(n68169), .O(n70213));
    defparam i50718_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n63131), .I1(n27889), .I2(VCC_net), 
            .I3(n52856), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8189[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51396_4_lut (.I0(n70239), .I1(n70745), .I2(n37_adj_5057), 
            .I3(n68161), .O(n70891));   // verilog/uart_rx.v(119[33:55])
    defparam i51396_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n53396), 
            .O(n8215[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_11 (.CI(n53396), .I0(n2722), .I1(n1879), .CO(n53397));
    SB_LUT4 add_2754_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n53395), 
            .O(n8215[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8189[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_10 (.CI(n53395), .I0(n2723), .I1(n1742), .CO(n53396));
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8189[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_25 (.CI(n52856), .I0(n27889), .I1(VCC_net), 
            .CO(n52857));
    SB_LUT4 add_2754_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n53394), 
            .O(n8215[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50891_4_lut (.I0(n70237), .I1(n69858), .I2(n27_adj_5067), 
            .I3(n69221), .O(n70386));   // verilog/uart_rx.v(119[33:55])
    defparam i50891_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n63187), .I1(n64567), .I2(VCC_net), 
            .I3(n52855), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8189[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51416_4_lut (.I0(n70386), .I1(n70891), .I2(n37_adj_5057), 
            .I3(n70213), .O(n70911));   // verilog/uart_rx.v(119[33:55])
    defparam i51416_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2754_9 (.CI(n53394), .I0(n2724), .I1(n1602), .CO(n53395));
    SB_LUT4 i51417_3_lut (.I0(n70911), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n70912));   // verilog/uart_rx.v(119[33:55])
    defparam i51417_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n53393), 
            .O(n8215[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_8 (.CI(n53393), .I0(n2725), .I1(n1459), .CO(n53394));
    SB_CARRY sub_38_add_2_24 (.CI(n52855), .I0(n64567), .I1(VCC_net), 
            .CO(n52856));
    SB_LUT4 add_2754_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n53392), 
            .O(n8215[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8189[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_7 (.CI(n53392), .I0(n2726), .I1(n1460), .CO(n53393));
    SB_LUT4 i51411_3_lut (.I0(n70912), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n70906));   // verilog/uart_rx.v(119[33:55])
    defparam i51411_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i534_3_lut (.I0(n60961), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n60965));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i51183_3_lut (.I0(n70906), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n70678));   // verilog/uart_rx.v(119[33:55])
    defparam i51183_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8163[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n53391), 
            .O(n8215[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8163[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51184_3_lut (.I0(n70678), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n70679));   // verilog/uart_rx.v(119[33:55])
    defparam i51184_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50750_3_lut (.I0(n70679), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam i50750_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8163[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_6 (.CI(n53391), .I0(n2727), .I1(n1011), .CO(n53392));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n52854), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8163[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n53390), 
            .O(n8215[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n53641), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n53640), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_8 (.CI(n53640), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n53641));
    SB_LUT4 r_Clock_Count_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n53639), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8163[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY r_Clock_Count_2053_add_4_7 (.CI(n53639), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n53640));
    SB_LUT4 r_Clock_Count_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n53638), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_6 (.CI(n53638), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n53639));
    SB_LUT4 r_Clock_Count_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n53637), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8293[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45_adj_5048), .I3(GND_net), .O(n40_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY r_Clock_Count_2053_add_4_5 (.CI(n53637), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n53638));
    SB_LUT4 r_Clock_Count_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n53636), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_5 (.CI(n53390), .I0(n2728), .I1(n856), .CO(n53391));
    SB_LUT4 i48944_4_lut (.I0(n43_adj_5065), .I1(n41), .I2(n39_adj_5058), 
            .I3(n68454), .O(n68439));
    defparam i48944_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY r_Clock_Count_2053_add_4_4 (.CI(n53636), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n53637));
    SB_CARRY sub_38_add_2_23 (.CI(n52854), .I0(n294[21]), .I1(VCC_net), 
            .CO(n52855));
    SB_LUT4 r_Clock_Count_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n53635), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_22_lut (.I0(n63185), .I1(n294[20]), .I2(VCC_net), 
            .I3(n52853), .O(n63187)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_22 (.CI(n52853), .I0(n294[20]), .I1(VCC_net), 
            .CO(n52854));
    SB_CARRY r_Clock_Count_2053_add_4_3 (.CI(n53635), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n53636));
    SB_LUT4 add_2754_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n53389), 
            .O(n8215[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n53635));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n63183), .I1(n294[19]), .I2(VCC_net), 
            .I3(n52852), .O(n63185)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_21 (.CI(n52852), .I0(n294[19]), .I1(VCC_net), 
            .CO(n52853));
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8293[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8163[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4045_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9625), .I3(n24106), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i4045_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 i50735_4_lut (.I0(n40_adj_5092), .I1(n20), .I2(n45_adj_5048), 
            .I3(n68431), .O(n70230));   // verilog/uart_rx.v(119[33:55])
    defparam i50735_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2754_4 (.CI(n53389), .I0(n2729), .I1(n698), .CO(n53390));
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i639_4_lut (.I0(n60965), .I1(n294[19]), .I2(n46), .I3(baudrate[4]), 
            .O(n60967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n52851), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n52851), .I0(n294[18]), .I1(VCC_net), 
            .CO(n52852));
    SB_LUT4 add_2754_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n53388), 
            .O(n8215[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_19_lut (.I0(n63181), .I1(n294[17]), .I2(VCC_net), 
            .I3(n52850), .O(n63183)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8163[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49693_3_lut (.I0(n70160), .I1(baudrate[15]), .I2(n41), .I3(GND_net), 
            .O(n69188));   // verilog/uart_rx.v(119[33:55])
    defparam i49693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8163[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_19 (.CI(n52850), .I0(n294[17]), .I1(VCC_net), 
            .CO(n52851));
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8163[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_3 (.CI(n53388), .I0(n2730), .I1(n858), .CO(n53389));
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n63179), .I1(n294[16]), .I2(VCC_net), 
            .I3(n52849), .O(n63181)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_18 (.CI(n52849), .I0(n294[16]), .I1(VCC_net), 
            .CO(n52850));
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8163[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8163[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_2_lut (.I0(n61266), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4216_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9796), .I3(n24124), 
            .O(n46_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam i4216_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8163[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i742_4_lut (.I0(n60967), .I1(n294[18]), .I2(n46_adj_5102), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8163[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n63129), .I1(n294[15]), .I2(VCC_net), 
            .I3(n52848), .O(n63131)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n52848), .I0(n294[15]), .I1(VCC_net), 
            .CO(n52849));
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8163[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18), .I1(baudrate[9]), 
            .I2(n29_adj_5072), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53388));
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8137[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n63177), .I1(n294[14]), .I2(VCC_net), 
            .I3(n52847), .O(n63179)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n52847), .I0(n294[14]), .I1(VCC_net), 
            .CO(n52848));
    SB_LUT4 i51157_4_lut (.I0(n26), .I1(n16_adj_5105), .I2(n29_adj_5072), 
            .I3(n68473), .O(n70652));   // verilog/uart_rx.v(119[33:55])
    defparam i51157_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2753_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n53387), 
            .O(n8189[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8137[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n52846), .O(n63177)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_15 (.CI(n52846), .I0(n294[13]), .I1(VCC_net), 
            .CO(n52847));
    SB_LUT4 add_2753_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n53386), 
            .O(n8189[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n52845), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_18 (.CI(n53386), .I0(n2597), .I1(n2754), .CO(n53387));
    SB_LUT4 add_2753_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n53385), 
            .O(n8189[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8137[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_14 (.CI(n52845), .I0(n294[12]), .I1(VCC_net), 
            .CO(n52846));
    SB_LUT4 i41822_1_lut (.I0(n27987), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61270));
    defparam i41822_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2753_17 (.CI(n53385), .I0(n2598), .I1(n2638), .CO(n53386));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n52844), .O(n63129)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n52844), .I0(n294[11]), .I1(VCC_net), 
            .CO(n52845));
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n53384), 
            .O(n8189[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n52843), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8137[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2753_16 (.CI(n53384), .I0(n2599), .I1(n2519), .CO(n53385));
    SB_LUT4 add_2753_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n53383), 
            .O(n8189[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n52843), .I0(n294[10]), .I1(VCC_net), 
            .CO(n52844));
    SB_CARRY add_2753_15 (.CI(n53383), .I0(n2600), .I1(n2397), .CO(n53384));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n52842), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8137[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2753_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n53382), 
            .O(n8189[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_14 (.CI(n53382), .I0(n2601), .I1(n2272), .CO(n53383));
    SB_LUT4 add_2753_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n53381), 
            .O(n8189[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2753_13 (.CI(n53381), .I0(n2602), .I1(n2144), .CO(n53382));
    SB_LUT4 add_2753_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n53380), 
            .O(n8189[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_12 (.CI(n53380), .I0(n2603), .I1(n2013), .CO(n53381));
    SB_LUT4 i51158_3_lut (.I0(n70652), .I1(baudrate[10]), .I2(n31_adj_5071), 
            .I3(GND_net), .O(n70653));   // verilog/uart_rx.v(119[33:55])
    defparam i51158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50978_3_lut (.I0(n70653), .I1(baudrate[11]), .I2(n33_adj_5079), 
            .I3(GND_net), .O(n70473));   // verilog/uart_rx.v(119[33:55])
    defparam i50978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50841_4_lut (.I0(n43_adj_5065), .I1(n41), .I2(n39_adj_5058), 
            .I3(n68456), .O(n70336));
    defparam i50841_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51213_4_lut (.I0(n69188), .I1(n70230), .I2(n45_adj_5048), 
            .I3(n68439), .O(n70708));   // verilog/uart_rx.v(119[33:55])
    defparam i51213_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49691_3_lut (.I0(n70473), .I1(baudrate[12]), .I2(n35_adj_5078), 
            .I3(GND_net), .O(n69186));   // verilog/uart_rx.v(119[33:55])
    defparam i49691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51215_4_lut (.I0(n69186), .I1(n70708), .I2(n45_adj_5048), 
            .I3(n70336), .O(n70710));   // verilog/uart_rx.v(119[33:55])
    defparam i51215_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(n63143), .I1(n48_adj_5109), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h2222;
    SB_LUT4 add_2753_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n53379), 
            .O(n8189[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_11 (.CI(n53379), .I0(n2604), .I1(n1879), .CO(n53380));
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7903[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8137[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8137[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8137[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7929[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8137[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7955[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n63861));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5113));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(r_Clock_Count[3]), .I1(n3_adj_5113), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n63861), .O(n63865));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n63865), .O(n63869));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'hffde;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7981[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8137[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5115));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8137[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(r_Clock_Count[6]), .I1(n8_adj_5115), 
            .I2(n63869), .I3(\o_Rx_DV_N_3488[7] ), .O(n59836));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'hfdfe;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59798));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8007[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8137[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8137[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8033[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44953_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n59836), .I2(GND_net), 
            .I3(GND_net), .O(n64439));
    defparam i44953_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8059[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8137[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45059_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n64439), .O(n64545));
    defparam i45059_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n63269), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i1_4_lut_adj_1010 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n63975));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n64545), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n10012));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n10012), .I1(n2), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i1_3_lut_adj_1011 (.I0(n63923), .I1(n63973), .I2(n63961), 
            .I3(GND_net), .O(n63983));
    defparam i1_3_lut_adj_1011.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(n63983), .I1(n63979), .I2(n63981), 
            .I3(n63975), .O(n27975));
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49117_4_lut (.I0(n25_adj_5121), .I1(n23_adj_5117), .I2(n21_adj_5116), 
            .I3(n19_adj_5123), .O(n68612));
    defparam i49117_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49105_4_lut (.I0(n31_adj_5119), .I1(n29_adj_5118), .I2(n27_adj_5122), 
            .I3(n68612), .O(n68600));
    defparam i49105_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50865_4_lut (.I0(n37_adj_5114), .I1(n35_adj_5112), .I2(n33_adj_5111), 
            .I3(n68600), .O(n70360));
    defparam i50865_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49230_4_lut (.I0(n33_adj_5125), .I1(n31_adj_5126), .I2(n29_adj_5127), 
            .I3(n27_adj_5124), .O(n68725));
    defparam i49230_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50676_3_lut (.I0(n18_adj_5128), .I1(baudrate[13]), .I2(n41_adj_5110), 
            .I3(GND_net), .O(n70171));   // verilog/uart_rx.v(119[33:55])
    defparam i50676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50677_3_lut (.I0(n70171), .I1(baudrate[14]), .I2(n43_adj_5108), 
            .I3(GND_net), .O(n70172));   // verilog/uart_rx.v(119[33:55])
    defparam i50677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5129), .I1(baudrate[10]), 
            .I2(n41_adj_5120), .I3(GND_net), .O(n38_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22901_rep_3_2_lut (.I0(n8059[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n61285));   // verilog/uart_rx.v(119[33:55])
    defparam i22901_rep_3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50059_4_lut (.I0(n43_adj_5108), .I1(n41_adj_5110), .I2(n29_adj_5118), 
            .I3(n68606), .O(n69554));
    defparam i50059_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5131), .I1(baudrate[7]), 
            .I2(n29_adj_5118), .I3(GND_net), .O(n26_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n61285), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i49675_3_lut (.I0(n70172), .I1(baudrate[15]), .I2(n45_adj_5107), 
            .I3(GND_net), .O(n69170));   // verilog/uart_rx.v(119[33:55])
    defparam i49675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2753_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n53378), 
            .O(n8189[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_10 (.CI(n53378), .I0(n2605), .I1(n1742), .CO(n53379));
    SB_LUT4 add_2753_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n53377), 
            .O(n8189[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_9 (.CI(n53377), .I0(n2606), .I1(n1602), .CO(n53378));
    SB_LUT4 add_2753_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n53376), 
            .O(n8189[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_8 (.CI(n53376), .I0(n2607), .I1(n1459), .CO(n53377));
    SB_LUT4 add_2753_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n53375), 
            .O(n8189[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_7 (.CI(n53375), .I0(n2608), .I1(n1460), .CO(n53376));
    SB_LUT4 add_2753_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n53374), 
            .O(n8189[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_6 (.CI(n53374), .I0(n2609), .I1(n1011), .CO(n53375));
    SB_LUT4 add_2753_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n53373), 
            .O(n8189[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_5 (.CI(n53373), .I0(n2610), .I1(n856), .CO(n53374));
    SB_LUT4 add_2753_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n53372), 
            .O(n8189[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_4 (.CI(n53372), .I0(n2611), .I1(n698), .CO(n53373));
    SB_LUT4 add_2753_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n53371), 
            .O(n8189[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5134), .I1(baudrate[9]), 
            .I2(n33_adj_5111), .I3(GND_net), .O(n30_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2753_3 (.CI(n53371), .I0(n2612), .I1(n858), .CO(n53372));
    SB_LUT4 add_2753_2_lut (.I0(n61270), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2753_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53371));
    SB_LUT4 add_2752_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n53370), 
            .O(n8163[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2752_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n53369), 
            .O(n8163[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_17 (.CI(n53369), .I0(n2477), .I1(n2638), .CO(n53370));
    SB_LUT4 i51151_4_lut (.I0(n30_adj_5135), .I1(n20_adj_5136), .I2(n33_adj_5111), 
            .I3(n68596), .O(n70646));   // verilog/uart_rx.v(119[33:55])
    defparam i51151_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2752_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n53368), 
            .O(n8163[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_16 (.CI(n53368), .I0(n2478), .I1(n2519), .CO(n53369));
    SB_LUT4 i51152_3_lut (.I0(n70646), .I1(baudrate[10]), .I2(n35_adj_5112), 
            .I3(GND_net), .O(n70647));   // verilog/uart_rx.v(119[33:55])
    defparam i51152_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_11 (.CI(n52842), .I0(n294[9]), .I1(VCC_net), 
            .CO(n52843));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n52841), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2752_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n53367), 
            .O(n8163[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_15 (.CI(n53367), .I0(n2479), .I1(n2397), .CO(n53368));
    SB_LUT4 add_2752_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n53366), 
            .O(n8163[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_14 (.CI(n53366), .I0(n2480), .I1(n2272), .CO(n53367));
    SB_LUT4 add_2752_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n53365), 
            .O(n8163[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_13 (.CI(n53365), .I0(n2481), .I1(n2144), .CO(n53366));
    SB_LUT4 add_2752_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n53364), 
            .O(n8163[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50690_3_lut (.I0(n26_adj_5133), .I1(baudrate[6]), .I2(n33_adj_5125), 
            .I3(GND_net), .O(n70185));   // verilog/uart_rx.v(119[33:55])
    defparam i50690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50990_3_lut (.I0(n70647), .I1(baudrate[11]), .I2(n37_adj_5114), 
            .I3(GND_net), .O(n70485));   // verilog/uart_rx.v(119[33:55])
    defparam i50990_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_12 (.CI(n53364), .I0(n2482), .I1(n2013), .CO(n53365));
    SB_LUT4 add_2752_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n53363), 
            .O(n8163[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_11 (.CI(n53363), .I0(n2483), .I1(n1879), .CO(n53364));
    SB_LUT4 i50065_4_lut (.I0(n43_adj_5108), .I1(n41_adj_5110), .I2(n39_adj_5106), 
            .I3(n70360), .O(n69560));
    defparam i50065_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2752_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n53362), 
            .O(n8163[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_10 (.CI(n53362), .I0(n2484), .I1(n1742), .CO(n53363));
    SB_LUT4 add_2752_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n53361), 
            .O(n8163[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_9 (.CI(n53361), .I0(n2485), .I1(n1602), .CO(n53362));
    SB_LUT4 add_2752_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n53360), 
            .O(n8163[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50730_4_lut (.I0(n69170), .I1(n26_adj_5132), .I2(n45_adj_5107), 
            .I3(n69554), .O(n70225));   // verilog/uart_rx.v(119[33:55])
    defparam i50730_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2752_8 (.CI(n53360), .I0(n2486), .I1(n1459), .CO(n53361));
    SB_LUT4 add_2752_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n53359), 
            .O(n8163[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_7 (.CI(n53359), .I0(n2487), .I1(n1460), .CO(n53360));
    SB_LUT4 add_2752_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n53358), 
            .O(n8163[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_6 (.CI(n53358), .I0(n2488), .I1(n1011), .CO(n53359));
    SB_LUT4 add_2752_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n53357), 
            .O(n8163[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n52841), .I0(n294[8]), .I1(VCC_net), 
            .CO(n52842));
    SB_CARRY add_2752_5 (.CI(n53357), .I0(n2489), .I1(n856), .CO(n53358));
    SB_LUT4 add_2752_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n53356), 
            .O(n8163[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_4 (.CI(n53356), .I0(n2490), .I1(n698), .CO(n53357));
    SB_LUT4 add_2752_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n53355), 
            .O(n8163[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_3 (.CI(n53355), .I0(n2491), .I1(n858), .CO(n53356));
    SB_LUT4 add_2752_2_lut (.I0(n61274), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2752_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53355));
    SB_LUT4 add_2751_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n53354), 
            .O(n8137[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2751_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n53353), 
            .O(n8137[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_16 (.CI(n53353), .I0(n2354), .I1(n2519), .CO(n53354));
    SB_LUT4 add_2751_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n53352), 
            .O(n8137[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_15 (.CI(n53352), .I0(n2355), .I1(n2397), .CO(n53353));
    SB_LUT4 i49673_3_lut (.I0(n70485), .I1(baudrate[12]), .I2(n39_adj_5106), 
            .I3(GND_net), .O(n69168));   // verilog/uart_rx.v(119[33:55])
    defparam i49673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n53351), 
            .O(n8137[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_14 (.CI(n53351), .I0(n2356), .I1(n2272), .CO(n53352));
    SB_LUT4 add_2751_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n53350), 
            .O(n8137[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_13 (.CI(n53350), .I0(n2357), .I1(n2144), .CO(n53351));
    SB_LUT4 add_2751_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n53349), 
            .O(n8137[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_12 (.CI(n53349), .I0(n2358), .I1(n2013), .CO(n53350));
    SB_LUT4 add_2751_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n53348), 
            .O(n8137[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_11 (.CI(n53348), .I0(n2359), .I1(n1879), .CO(n53349));
    SB_LUT4 i50732_4_lut (.I0(n69168), .I1(n70225), .I2(n45_adj_5107), 
            .I3(n69560), .O(n70227));   // verilog/uart_rx.v(119[33:55])
    defparam i50732_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2751_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n53347), 
            .O(n8137[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_10 (.CI(n53347), .I0(n2360), .I1(n1742), .CO(n53348));
    SB_LUT4 add_2751_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n53346), 
            .O(n8137[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_9 (.CI(n53346), .I0(n2361), .I1(n1602), .CO(n53347));
    SB_LUT4 add_2751_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n53345), 
            .O(n8137[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_8 (.CI(n53345), .I0(n2362), .I1(n1459), .CO(n53346));
    SB_LUT4 add_2751_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n53344), 
            .O(n8137[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_7 (.CI(n53344), .I0(n2363), .I1(n1460), .CO(n53345));
    SB_LUT4 add_2751_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n53343), 
            .O(n8137[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_6 (.CI(n53343), .I0(n2364), .I1(n1011), .CO(n53344));
    SB_LUT4 add_2751_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n53342), 
            .O(n8137[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_5 (.CI(n53342), .I0(n2365), .I1(n856), .CO(n53343));
    SB_LUT4 add_2751_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n53341), 
            .O(n8137[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_4 (.CI(n53341), .I0(n2366), .I1(n698), .CO(n53342));
    SB_LUT4 add_2751_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n53340), 
            .O(n8137[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_3 (.CI(n53340), .I0(n2367), .I1(n858), .CO(n53341));
    SB_LUT4 add_2751_2_lut (.I0(n61278), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2751_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53340));
    SB_LUT4 add_2750_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n53339), 
            .O(n8111[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2750_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n53338), 
            .O(n8111[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_15 (.CI(n53338), .I0(n2228), .I1(n2397), .CO(n53339));
    SB_LUT4 add_2750_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n53337), 
            .O(n8111[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_14 (.CI(n53337), .I0(n2229), .I1(n2272), .CO(n53338));
    SB_LUT4 add_2750_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n53336), 
            .O(n8111[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_13 (.CI(n53336), .I0(n2230), .I1(n2144), .CO(n53337));
    SB_LUT4 add_2750_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n53335), 
            .O(n8111[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_12 (.CI(n53335), .I0(n2231), .I1(n2013), .CO(n53336));
    SB_LUT4 add_2750_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n53334), 
            .O(n8111[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n52840), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_11 (.CI(n53334), .I0(n2232), .I1(n1879), .CO(n53335));
    SB_LUT4 add_2750_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n53333), 
            .O(n8111[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n53488), 
            .O(n8319[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8111[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2750_10 (.CI(n53333), .I0(n2233), .I1(n1742), .CO(n53334));
    SB_LUT4 add_2750_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n53332), 
            .O(n8111[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_9 (.CI(n53332), .I0(n2234), .I1(n1602), .CO(n53333));
    SB_LUT4 add_2750_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n53331), 
            .O(n8111[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_8 (.CI(n53331), .I0(n2235), .I1(n1459), .CO(n53332));
    SB_LUT4 add_2750_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n53330), 
            .O(n8111[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_7 (.CI(n53330), .I0(n2236), .I1(n1460), .CO(n53331));
    SB_LUT4 add_2750_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n53329), 
            .O(n8111[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n53487), 
            .O(n8319[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_6 (.CI(n53329), .I0(n2237), .I1(n1011), .CO(n53330));
    SB_LUT4 i50691_3_lut (.I0(n70185), .I1(baudrate[7]), .I2(n35_adj_5137), 
            .I3(GND_net), .O(n70186));   // verilog/uart_rx.v(119[33:55])
    defparam i50691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n53328), 
            .O(n8111[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_5 (.CI(n53328), .I0(n2238), .I1(n856), .CO(n53329));
    SB_LUT4 add_2750_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n53327), 
            .O(n8111[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_4 (.CI(n53327), .I0(n2239), .I1(n698), .CO(n53328));
    SB_LUT4 add_2750_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n53326), 
            .O(n8111[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_3 (.CI(n53326), .I0(n2240), .I1(n858), .CO(n53327));
    SB_LUT4 add_2750_2_lut (.I0(n61282), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2750_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53326));
    SB_LUT4 add_2749_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n53325), 
            .O(n8085[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2749_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n53324), 
            .O(n8085[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_13 (.CI(n53324), .I0(n2099), .I1(n2272), .CO(n53325));
    SB_LUT4 add_2749_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n53323), 
            .O(n8085[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_12 (.CI(n53323), .I0(n2100), .I1(n2144), .CO(n53324));
    SB_LUT4 add_2749_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n53322), 
            .O(n8085[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_11 (.CI(n53322), .I0(n2101), .I1(n2013), .CO(n53323));
    SB_LUT4 add_2749_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n53321), 
            .O(n8085[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_10 (.CI(n53321), .I0(n2102), .I1(n1879), .CO(n53322));
    SB_LUT4 add_2749_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n53320), 
            .O(n8085[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_9 (.CI(n53320), .I0(n2103), .I1(n1742), .CO(n53321));
    SB_LUT4 add_2749_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n53319), 
            .O(n8085[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_8 (.CI(n53319), .I0(n2104), .I1(n1602), .CO(n53320));
    SB_CARRY sub_38_add_2_9 (.CI(n52840), .I0(n294[7]), .I1(VCC_net), 
            .CO(n52841));
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8111[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n53318), 
            .O(n8085[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_7 (.CI(n53318), .I0(n2105), .I1(n1459), .CO(n53319));
    SB_LUT4 add_2749_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n53317), 
            .O(n8085[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_6 (.CI(n53317), .I0(n2106), .I1(n1460), .CO(n53318));
    SB_LUT4 add_2749_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n53316), 
            .O(n8085[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_5 (.CI(n53316), .I0(n2107), .I1(n1011), .CO(n53317));
    SB_LUT4 add_2749_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n53315), 
            .O(n8085[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_4 (.CI(n53315), .I0(n2108), .I1(n856), .CO(n53316));
    SB_LUT4 add_2749_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n53314), 
            .O(n8085[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_3 (.CI(n53314), .I0(n2109), .I1(n698), .CO(n53315));
    SB_LUT4 add_2749_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8085[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n53314));
    SB_LUT4 add_2748_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n53313), 
            .O(n8059[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2748_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n53312), 
            .O(n8059[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_13 (.CI(n53312), .I0(n1967), .I1(n2144), .CO(n53313));
    SB_LUT4 add_2748_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n53311), 
            .O(n8059[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_12 (.CI(n53311), .I0(n1968), .I1(n2013), .CO(n53312));
    SB_LUT4 add_2748_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n53310), 
            .O(n8059[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_11 (.CI(n53310), .I0(n1969), .I1(n1879), .CO(n53311));
    SB_LUT4 add_2748_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n53309), 
            .O(n8059[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_10 (.CI(n53309), .I0(n1970), .I1(n1742), .CO(n53310));
    SB_LUT4 add_2748_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n53308), 
            .O(n8059[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_9 (.CI(n53308), .I0(n1971), .I1(n1602), .CO(n53309));
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8111[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n53307), 
            .O(n8059[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_8 (.CI(n53307), .I0(n1972), .I1(n1459), .CO(n53308));
    SB_LUT4 add_2748_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n53306), 
            .O(n8059[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_7 (.CI(n53306), .I0(n1973), .I1(n1460), .CO(n53307));
    SB_DFFESR r_Clock_Count_2053__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n30202), .D(n1[0]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5138), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2748_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n53305), 
            .O(n8059[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n52839), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_6 (.CI(n53305), .I0(n1974), .I1(n1011), .CO(n53306));
    SB_LUT4 add_2748_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n53304), 
            .O(n8059[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n52839), .I0(n294[6]), .I1(VCC_net), 
            .CO(n52840));
    SB_CARRY add_2748_5 (.CI(n53304), .I0(n1975), .I1(n856), .CO(n53305));
    SB_LUT4 add_2748_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n53303), 
            .O(n8059[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n52838), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_4 (.CI(n53303), .I0(n1976), .I1(n698), .CO(n53304));
    SB_LUT4 add_2748_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n53302), 
            .O(n8059[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_3 (.CI(n53302), .I0(n1977), .I1(n858), .CO(n53303));
    SB_CARRY add_2758_24 (.CI(n53487), .I0(n3152), .I1(n3082), .CO(n53488));
    SB_LUT4 add_2748_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8059[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53302));
    SB_LUT4 add_2747_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n53301), 
            .O(n8033[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n53300), 
            .O(n8033[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n52838), .I0(n294[5]), .I1(VCC_net), 
            .CO(n52839));
    SB_CARRY add_2747_12 (.CI(n53300), .I0(n1832), .I1(n2013), .CO(n53301));
    SB_LUT4 add_2747_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n53299), 
            .O(n8033[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n52837), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_11 (.CI(n53299), .I0(n1833), .I1(n1879), .CO(n53300));
    SB_LUT4 i49214_4_lut (.I0(n39_adj_5139), .I1(n37_adj_5056), .I2(n35_adj_5137), 
            .I3(n68725), .O(n68709));
    defparam i49214_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8111[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8111[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51145_4_lut (.I0(n38_adj_5130), .I1(n28), .I2(n41_adj_5120), 
            .I3(n68706), .O(n70640));   // verilog/uart_rx.v(119[33:55])
    defparam i51145_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_38_add_2_6 (.CI(n52837), .I0(n294[4]), .I1(VCC_net), 
            .CO(n52838));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n52836), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n53298), 
            .O(n8033[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_10 (.CI(n53298), .I0(n1834), .I1(n1742), .CO(n53299));
    SB_LUT4 add_2747_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n53297), 
            .O(n8033[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n53486), 
            .O(n8319[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_9 (.CI(n53297), .I0(n1835), .I1(n1602), .CO(n53298));
    SB_CARRY sub_38_add_2_5 (.CI(n52836), .I0(n294[3]), .I1(VCC_net), 
            .CO(n52837));
    SB_LUT4 add_2747_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n53296), 
            .O(n8033[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_8 (.CI(n53296), .I0(n1836), .I1(n1459), .CO(n53297));
    SB_CARRY add_2758_23 (.CI(n53486), .I0(n3153), .I1(n3188), .CO(n53487));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n52835), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n53295), 
            .O(n8033[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_7 (.CI(n53295), .I0(n1837), .I1(n1460), .CO(n53296));
    SB_LUT4 add_2758_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n53485), 
            .O(n8319[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n53294), 
            .O(n8033[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n52835), .I0(n294[2]), .I1(VCC_net), 
            .CO(n52836));
    SB_CARRY add_2747_6 (.CI(n53294), .I0(n1838), .I1(n1011), .CO(n53295));
    SB_CARRY add_2758_22 (.CI(n53485), .I0(n3154), .I1(n3084), .CO(n53486));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n52834), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n53293), 
            .O(n8033[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_5 (.CI(n53293), .I0(n1839), .I1(n856), .CO(n53294));
    SB_CARRY sub_38_add_2_3 (.CI(n52834), .I0(n294[1]), .I1(VCC_net), 
            .CO(n52835));
    SB_LUT4 add_2747_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n53292), 
            .O(n8033[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n62087), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n53484), 
            .O(n8319[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_4 (.CI(n53292), .I0(n1840), .I1(n698), .CO(n53293));
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n62087), .I1(GND_net), 
            .CO(n52834));
    SB_LUT4 add_2747_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n53291), 
            .O(n8033[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_3 (.CI(n53291), .I0(n1841), .I1(n858), .CO(n53292));
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8111[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2758_21 (.CI(n53484), .I0(n3155), .I1(n2977), .CO(n53485));
    SB_LUT4 add_2747_2_lut (.I0(n61291), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2747_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53291));
    SB_LUT4 add_2758_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n53483), 
            .O(n8319[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2758_20 (.CI(n53483), .I0(n3156), .I1(n2867), .CO(n53484));
    SB_LUT4 add_2758_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n53482), 
            .O(n8319[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_19 (.CI(n53482), .I0(n3157), .I1(n2754), .CO(n53483));
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8111[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Clock_Count_2053__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n30202), .D(n1[7]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n30202), .D(n1[6]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n30202), .D(n1[5]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n30202), .D(n1[4]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n30202), .D(n1[3]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n30202), .D(n1[2]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n30202), .D(n1[1]), .R(n31416));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i49653_3_lut (.I0(n70186), .I1(baudrate[8]), .I2(n37_adj_5056), 
            .I3(GND_net), .O(n69148));   // verilog/uart_rx.v(119[33:55])
    defparam i49653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51345_4_lut (.I0(n69148), .I1(n70640), .I2(n41_adj_5120), 
            .I3(n68709), .O(n70840));   // verilog/uart_rx.v(119[33:55])
    defparam i51345_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8111[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n53481), 
            .O(n8319[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_18 (.CI(n53481), .I0(n3158), .I1(n2638), .CO(n53482));
    SB_LUT4 add_2758_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n53480), 
            .O(n8319[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2746_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n53280), 
            .O(n8007[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_17 (.CI(n53480), .I0(n3159), .I1(n2519), .CO(n53481));
    SB_LUT4 add_2746_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n53279), 
            .O(n8007[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_10 (.CI(n53279), .I0(n1694), .I1(n1879), .CO(n53280));
    SB_LUT4 i51346_3_lut (.I0(n70840), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n70841));   // verilog/uart_rx.v(119[33:55])
    defparam i51346_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51279_3_lut (.I0(n70841), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n70774));   // verilog/uart_rx.v(119[33:55])
    defparam i51279_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2746_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n53278), 
            .O(n8007[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_9 (.CI(n53278), .I0(n1695), .I1(n1742), .CO(n53279));
    SB_LUT4 add_2746_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n53277), 
            .O(n8007[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n53479), 
            .O(n8319[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_16 (.CI(n53479), .I0(n3160), .I1(n2397), .CO(n53480));
    SB_CARRY add_2746_8 (.CI(n53277), .I0(n1696), .I1(n1602), .CO(n53278));
    SB_LUT4 add_2746_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n53276), 
            .O(n8007[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n53478), 
            .O(n8319[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_15 (.CI(n53478), .I0(n3161), .I1(n2272), .CO(n53479));
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2746_7 (.CI(n53276), .I0(n1697), .I1(n1459), .CO(n53277));
    SB_LUT4 add_2746_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n53275), 
            .O(n8007[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n53477), 
            .O(n8319[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_14 (.CI(n53477), .I0(n3162), .I1(n2144), .CO(n53478));
    SB_CARRY add_2746_6 (.CI(n53275), .I0(n1698), .I1(n1460), .CO(n53276));
    SB_LUT4 add_2746_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n53274), 
            .O(n8007[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_5 (.CI(n53274), .I0(n1699), .I1(n1011), .CO(n53275));
    SB_LUT4 add_2746_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n53273), 
            .O(n8007[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_4 (.CI(n53273), .I0(n1700), .I1(n856), .CO(n53274));
    SB_LUT4 add_2746_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n53272), 
            .O(n8007[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n53476), 
            .O(n8319[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_3 (.CI(n53272), .I0(n1701), .I1(n698), .CO(n53273));
    SB_CARRY add_2758_13 (.CI(n53476), .I0(n3163), .I1(n2013), .CO(n53477));
    SB_LUT4 add_2758_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n53475), 
            .O(n8319[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_12 (.CI(n53475), .I0(n3164), .I1(n1879), .CO(n53476));
    SB_LUT4 add_2746_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8007[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n53474), 
            .O(n8319[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_11 (.CI(n53474), .I0(n3165), .I1(n1742), .CO(n53475));
    SB_CARRY add_2746_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n53272));
    SB_LUT4 add_2758_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n53473), 
            .O(n8319[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n53271), 
            .O(n7981[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_10 (.CI(n53473), .I0(n3166), .I1(n1602), .CO(n53474));
    SB_LUT4 add_2745_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n53270), 
            .O(n7981[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_10 (.CI(n53270), .I0(n1553), .I1(n1742), .CO(n53271));
    SB_LUT4 i49659_3_lut (.I0(n70774), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam i49659_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2745_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n53269), 
            .O(n7981[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_9 (.CI(n53269), .I0(n1554), .I1(n1602), .CO(n53270));
    SB_LUT4 add_2758_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n53472), 
            .O(n8319[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_9 (.CI(n53472), .I0(n3167), .I1(n1459), .CO(n53473));
    SB_LUT4 add_2758_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n53471), 
            .O(n8319[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n53268), 
            .O(n7981[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_8 (.CI(n53471), .I0(n3168), .I1(n1460), .CO(n53472));
    SB_LUT4 add_2758_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n53470), 
            .O(n8319[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_8 (.CI(n53268), .I0(n1555), .I1(n1459), .CO(n53269));
    SB_LUT4 add_2745_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n53267), 
            .O(n7981[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49067_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5230), .I3(\o_Rx_DV_N_3488[8] ), .O(n67678));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49067_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i49163_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n59836), 
            .I3(r_SM_Main[0]), .O(n67684));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49163_4_lut.LUT_INIT = 16'h0100;
    SB_CARRY add_2745_7 (.CI(n53267), .I0(n1556), .I1(n1460), .CO(n53268));
    SB_CARRY add_2758_7 (.CI(n53470), .I0(n3169), .I1(n1011), .CO(n53471));
    SB_LUT4 add_2758_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n53469), 
            .O(n8319[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_6 (.CI(n53469), .I0(n3170), .I1(n856), .CO(n53470));
    SB_LUT4 i1_2_lut_adj_1013 (.I0(n63141), .I1(n48_adj_5046), .I2(GND_net), 
            .I3(GND_net), .O(n2367));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h2222;
    SB_LUT4 add_2758_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n53468), 
            .O(n8319[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_5 (.CI(n53468), .I0(n3171), .I1(n698), .CO(n53469));
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8111[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49064_4_lut (.I0(n67678), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67675));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49064_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2758_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n53467), 
            .O(n8319[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_4 (.CI(n53467), .I0(n3172), .I1(n858), .CO(n53468));
    SB_LUT4 add_2758_3_lut (.I0(n61250), .I1(GND_net), .I2(n538), .I3(n53466), 
            .O(n63157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8059[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8111[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49070_4_lut (.I0(n67684), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67681));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49070_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8085[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2758_3 (.CI(n53466), .I0(GND_net), .I1(n538), .CO(n53467));
    SB_CARRY add_2758_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n53466));
    SB_LUT4 add_2745_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n53266), 
            .O(n7981[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8085[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2745_6 (.CI(n53266), .I0(n1557), .I1(n1011), .CO(n53267));
    SB_LUT4 add_2757_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n53465), 
            .O(n8293[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n67681), .I1(n67675), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5138));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 add_2757_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n53464), 
            .O(n8293[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n53265), 
            .O(n7981[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8111[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2745_5 (.CI(n53265), .I0(n1558), .I1(n856), .CO(n53266));
    SB_CARRY add_2757_22 (.CI(n53464), .I0(n3047), .I1(n3188), .CO(n53465));
    SB_LUT4 add_2757_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n53463), 
            .O(n8293[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n53264), 
            .O(n7981[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8111[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2757_21 (.CI(n53463), .I0(n3048), .I1(n3084), .CO(n53464));
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8085[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2745_4 (.CI(n53264), .I0(n1559), .I1(n698), .CO(n53265));
    SB_LUT4 add_2757_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n53462), 
            .O(n8293[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_20 (.CI(n53462), .I0(n3049), .I1(n2977), .CO(n53463));
    SB_LUT4 add_2757_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n53461), 
            .O(n8293[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2757_19 (.CI(n53461), .I0(n3050), .I1(n2867), .CO(n53462));
    SB_LUT4 add_2757_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n53460), 
            .O(n8293[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2757_18 (.CI(n53460), .I0(n3051), .I1(n2754), .CO(n53461));
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2745_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n53263), 
            .O(n7981[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n53459), 
            .O(n8293[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49195_4_lut (.I0(n29_adj_5151), .I1(n27_adj_5148), .I2(n25_adj_5147), 
            .I3(n23_adj_5157), .O(n68690));
    defparam i49195_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49274_4_lut (.I0(n33_adj_5159), .I1(n31_adj_5158), .I2(n29_adj_5156), 
            .I3(n27_adj_5160), .O(n68769));
    defparam i49274_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49185_4_lut (.I0(n35_adj_5161), .I1(n33_adj_5162), .I2(n31_adj_5153), 
            .I3(n68690), .O(n68680));
    defparam i49185_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2745_3 (.CI(n53263), .I0(n1560), .I1(n858), .CO(n53264));
    SB_LUT4 add_2745_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7981[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53263));
    SB_LUT4 add_2744_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n53262), 
            .O(n7955[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49284_2_lut (.I0(n59836), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n67631));
    defparam i49284_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_2744_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n53261), 
            .O(n7955[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_17 (.CI(n53459), .I0(n3052), .I1(n2638), .CO(n53460));
    SB_CARRY add_2744_9 (.CI(n53261), .I0(n1409), .I1(n1602), .CO(n53262));
    SB_LUT4 add_2757_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n53458), 
            .O(n8293[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5163), .I1(baudrate[9]), 
            .I2(n41_adj_5154), .I3(GND_net), .O(n38_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2744_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n53260), 
            .O(n7955[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_8 (.CI(n53260), .I0(n1410), .I1(n1459), .CO(n53261));
    SB_LUT4 i49279_4_lut (.I0(n67631), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n67628));
    defparam i49279_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2744_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n53259), 
            .O(n7955[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48568_4_lut (.I0(n67628), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n67625));
    defparam i48568_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY add_2744_7 (.CI(n53259), .I0(n1411), .I1(n1460), .CO(n53260));
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5167), .I1(baudrate[7]), 
            .I2(n33_adj_5162), .I3(GND_net), .O(n30_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50698_3_lut (.I0(n26_adj_5166), .I1(baudrate[5]), .I2(n33_adj_5159), 
            .I3(GND_net), .O(n70193));   // verilog/uart_rx.v(119[33:55])
    defparam i50698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50699_3_lut (.I0(n70193), .I1(baudrate[6]), .I2(n35_adj_5152), 
            .I3(GND_net), .O(n70194));   // verilog/uart_rx.v(119[33:55])
    defparam i50699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2744_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n53258), 
            .O(n7955[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51610_4_lut (.I0(r_SM_Main[2]), .I1(n67625), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(r_SM_Main[1]), .O(n31416));
    defparam i51610_4_lut.LUT_INIT = 16'h0511;
    SB_CARRY add_2757_16 (.CI(n53458), .I0(n3053), .I1(n2519), .CO(n53459));
    SB_LUT4 i49258_4_lut (.I0(n39_adj_5155), .I1(n37_adj_5150), .I2(n35_adj_5152), 
            .I3(n68769), .O(n68753));
    defparam i49258_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51141_4_lut (.I0(n38_adj_5164), .I1(n28_adj_5169), .I2(n41_adj_5154), 
            .I3(n68742), .O(n70636));   // verilog/uart_rx.v(119[33:55])
    defparam i51141_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49645_3_lut (.I0(n70194), .I1(baudrate[7]), .I2(n37_adj_5150), 
            .I3(GND_net), .O(n69140));   // verilog/uart_rx.v(119[33:55])
    defparam i49645_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2744_6 (.CI(n53258), .I0(n1412), .I1(n1011), .CO(n53259));
    SB_LUT4 add_2757_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n53457), 
            .O(n8293[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5170), .I1(baudrate[9]), 
            .I2(n37_adj_5171), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2744_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n53257), 
            .O(n7955[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51343_4_lut (.I0(n69140), .I1(n70636), .I2(n41_adj_5154), 
            .I3(n68753), .O(n70838));   // verilog/uart_rx.v(119[33:55])
    defparam i51343_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51147_4_lut (.I0(n34), .I1(n24_adj_5172), .I2(n37_adj_5171), 
            .I3(n68674), .O(n70642));   // verilog/uart_rx.v(119[33:55])
    defparam i51147_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51148_3_lut (.I0(n70642), .I1(baudrate[10]), .I2(n39_adj_5173), 
            .I3(GND_net), .O(n70643));   // verilog/uart_rx.v(119[33:55])
    defparam i51148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51344_3_lut (.I0(n70838), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n70839));   // verilog/uart_rx.v(119[33:55])
    defparam i51344_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51281_3_lut (.I0(n70839), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n70776));   // verilog/uart_rx.v(119[33:55])
    defparam i51281_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49651_3_lut (.I0(n70776), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam i49651_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2744_5 (.CI(n53257), .I0(n1413), .I1(n856), .CO(n53258));
    SB_LUT4 add_2744_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n53256), 
            .O(n7955[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_4 (.CI(n53256), .I0(n1414), .I1(n698), .CO(n53257));
    SB_LUT4 add_2744_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n53255), 
            .O(n7955[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n59836), .I1(r_SM_Main[1]), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n63211));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'h1000;
    SB_CARRY add_2744_3 (.CI(n53255), .I0(n1415), .I1(n858), .CO(n53256));
    SB_LUT4 add_2744_2_lut (.I0(n61300), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i50994_3_lut (.I0(n70643), .I1(baudrate[11]), .I2(n41_adj_5175), 
            .I3(GND_net), .O(n70489));   // verilog/uart_rx.v(119[33:55])
    defparam i50994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50873_4_lut (.I0(n41_adj_5175), .I1(n39_adj_5173), .I2(n37_adj_5171), 
            .I3(n68680), .O(n70368));
    defparam i50873_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1015 (.I0(n64467), .I1(n48_adj_5174), .I2(n8059[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_1015.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n63211), .O(n63217));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h0100;
    SB_CARRY add_2744_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53255));
    SB_LUT4 add_2743_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n53254), 
            .O(n7929[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n53253), 
            .O(n7929[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_8 (.CI(n53253), .I0(n1262), .I1(n1459), .CO(n53254));
    SB_LUT4 i51471_4_lut (.I0(r_SM_Main[2]), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n63217), .O(n30202));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i51471_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i50903_4_lut (.I0(n30_adj_5168), .I1(n22_adj_5165), .I2(n33_adj_5162), 
            .I3(n68682), .O(n70398));   // verilog/uart_rx.v(119[33:55])
    defparam i50903_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49663_3_lut (.I0(n70489), .I1(baudrate[12]), .I2(n43_adj_5178), 
            .I3(GND_net), .O(n69158));   // verilog/uart_rx.v(119[33:55])
    defparam i49663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2743_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n53252), 
            .O(n7929[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_7 (.CI(n53252), .I0(n1263), .I1(n1460), .CO(n53253));
    SB_LUT4 add_2743_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n53251), 
            .O(n7929[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_6 (.CI(n53251), .I0(n1264), .I1(n1011), .CO(n53252));
    SB_LUT4 add_2743_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n53250), 
            .O(n7929[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_5 (.CI(n53250), .I0(n1265), .I1(n856), .CO(n53251));
    SB_LUT4 add_2743_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n53249), 
            .O(n7929[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51135_4_lut (.I0(n69158), .I1(n70398), .I2(n43_adj_5178), 
            .I3(n70368), .O(n70630));   // verilog/uart_rx.v(119[33:55])
    defparam i51135_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51136_3_lut (.I0(n70630), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n70631));   // verilog/uart_rx.v(119[33:55])
    defparam i51136_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51022_3_lut (.I0(n70631), .I1(baudrate[14]), .I2(n2227), 
            .I3(GND_net), .O(n48_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam i51022_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2743_4 (.CI(n53249), .I0(n1266), .I1(n698), .CO(n53250));
    SB_LUT4 add_2743_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n53248), 
            .O(n7929[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8085[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50905_3_lut (.I0(n34_adj_5181), .I1(baudrate[5]), .I2(n41_adj_5180), 
            .I3(GND_net), .O(n70400));   // verilog/uart_rx.v(119[33:55])
    defparam i50905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50906_3_lut (.I0(n70400), .I1(baudrate[6]), .I2(n43_adj_5179), 
            .I3(GND_net), .O(n70401));   // verilog/uart_rx.v(119[33:55])
    defparam i50906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49350_4_lut (.I0(n43_adj_5179), .I1(n41_adj_5180), .I2(n39_adj_5177), 
            .I3(n67826), .O(n68845));
    defparam i49350_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8111[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39_adj_5177), 
            .I3(GND_net), .O(n38_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2743_3 (.CI(n53248), .I0(n1267), .I1(n858), .CO(n53249));
    SB_LUT4 add_2743_2_lut (.I0(n61304), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2743_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53248));
    SB_LUT4 add_2742_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n53247), 
            .O(n7903[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50717_3_lut (.I0(n70401), .I1(baudrate[7]), .I2(n45_adj_5176), 
            .I3(GND_net), .O(n44_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam i50717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50351_4_lut (.I0(n44_adj_5184), .I1(n38_adj_5182), .I2(n45_adj_5176), 
            .I3(n68845), .O(n69846));   // verilog/uart_rx.v(119[33:55])
    defparam i50351_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7981[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2742_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n53246), 
            .O(n7903[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_7 (.CI(n53246), .I0(n1112), .I1(n1460), .CO(n53247));
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8007[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8033[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49146_4_lut (.I0(n27_adj_5186), .I1(n25_adj_5185), .I2(n23_adj_5183), 
            .I3(n21_adj_5187), .O(n68641));
    defparam i49146_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8059[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8085[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2742_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n53245), 
            .O(n7903[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_6 (.CI(n53245), .I0(n1113), .I1(n1011), .CO(n53246));
    SB_LUT4 add_2742_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n53244), 
            .O(n7903[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_5 (.CI(n53244), .I0(n1114), .I1(n856), .CO(n53245));
    SB_LUT4 add_2742_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n53243), 
            .O(n7903[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_4 (.CI(n53243), .I0(n1115), .I1(n698), .CO(n53244));
    SB_LUT4 add_2742_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n53242), 
            .O(n7903[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_3 (.CI(n53242), .I0(n1116), .I1(n858), .CO(n53243));
    SB_LUT4 add_2742_2_lut (.I0(n61308), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2742_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53242));
    SB_CARRY add_2757_15 (.CI(n53457), .I0(n3054), .I1(n2397), .CO(n53458));
    SB_LUT4 add_2757_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n53456), 
            .O(n8293[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_14 (.CI(n53456), .I0(n3055), .I1(n2272), .CO(n53457));
    SB_LUT4 add_2757_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n53455), 
            .O(n8293[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_13 (.CI(n53455), .I0(n3056), .I1(n2144), .CO(n53456));
    SB_LUT4 add_2757_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n53454), 
            .O(n8293[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_12 (.CI(n53454), .I0(n3057), .I1(n2013), .CO(n53455));
    SB_LUT4 add_2757_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n53453), 
            .O(n8293[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_11 (.CI(n53453), .I0(n3058), .I1(n1879), .CO(n53454));
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8085[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2757_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n53452), 
            .O(n8293[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_10 (.CI(n53452), .I0(n3059), .I1(n1742), .CO(n53453));
    SB_LUT4 add_2757_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n53451), 
            .O(n8293[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_9 (.CI(n53451), .I0(n3060), .I1(n1602), .CO(n53452));
    SB_LUT4 add_2757_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n53450), 
            .O(n8293[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_8 (.CI(n53450), .I0(n3061), .I1(n1459), .CO(n53451));
    SB_LUT4 add_2757_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n53449), 
            .O(n8293[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8085[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2757_7 (.CI(n53449), .I0(n3062), .I1(n1460), .CO(n53450));
    SB_LUT4 add_2757_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n53448), 
            .O(n8293[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_6 (.CI(n53448), .I0(n3063), .I1(n1011), .CO(n53449));
    SB_LUT4 add_2757_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n53447), 
            .O(n8293[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1017 (.I0(n70910), .I1(baudrate[20]), .I2(n2938), 
            .I3(n63153), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1017.LUT_INIT = 16'h7100;
    SB_LUT4 i51520_2_lut_4_lut (.I0(n70910), .I1(baudrate[20]), .I2(n2938), 
            .I3(n64527), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i51520_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2757_5 (.CI(n53447), .I0(n3064), .I1(n856), .CO(n53448));
    SB_LUT4 add_2757_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n53446), 
            .O(n8293[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1018 (.I0(n70898), .I1(baudrate[19]), .I2(n2827), 
            .I3(n63151), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1018.LUT_INIT = 16'h7100;
    SB_LUT4 i49137_4_lut (.I0(n33_adj_5146), .I1(n31_adj_5145), .I2(n29_adj_5149), 
            .I3(n68641), .O(n68632));
    defparam i49137_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51517_2_lut_4_lut (.I0(n70898), .I1(baudrate[19]), .I2(n2827), 
            .I3(n27993), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i51517_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63711), .I1(n64533), .I2(baudrate[0]), 
            .I3(n48_adj_5053), .O(n962));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_CARRY add_2757_4 (.CI(n53446), .I0(n3065), .I1(n698), .CO(n53447));
    SB_LUT4 add_2757_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n53445), 
            .O(n8293[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n32278));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .D(n55993));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n30084), 
            .D(n479[1]), .R(n31398));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2757_3 (.CI(n53445), .I0(n3066), .I1(n858), .CO(n53446));
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n30084), 
            .D(n479[2]), .R(n31398));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n32606));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n32605));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n32604));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n32603));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n32600));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n32599));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n32598));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2757_2_lut (.I0(n61254), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2757_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53445));
    SB_LUT4 add_2756_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n53444), 
            .O(n8267[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2756_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n53443), 
            .O(n8267[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_21 (.CI(n53443), .I0(n2939), .I1(n3084), .CO(n53444));
    SB_LUT4 add_2756_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n53442), 
            .O(n8267[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8085[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_20 (.CI(n53442), .I0(n2940), .I1(n2977), .CO(n53443));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n32286));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8033[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n71751));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2756_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n53441), 
            .O(n8267[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8059[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_19 (.CI(n53441), .I0(n2941), .I1(n2867), .CO(n53442));
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8085[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2756_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n53440), 
            .O(n8267[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_18 (.CI(n53440), .I0(n2942), .I1(n2754), .CO(n53441));
    SB_LUT4 add_2756_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n53439), 
            .O(n8267[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_17 (.CI(n53439), .I0(n2943), .I1(n2638), .CO(n53440));
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5188), .I1(baudrate[7]), 
            .I2(n31_adj_5145), .I3(GND_net), .O(n28_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2756_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n53438), 
            .O(n8267[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_16 (.CI(n53438), .I0(n2944), .I1(n2519), .CO(n53439));
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2756_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n53437), 
            .O(n8267[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_15 (.CI(n53437), .I0(n2945), .I1(n2397), .CO(n53438));
    SB_LUT4 add_2756_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n53436), 
            .O(n8267[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_14 (.CI(n53436), .I0(n2946), .I1(n2272), .CO(n53437));
    SB_LUT4 add_2756_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n53435), 
            .O(n8267[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_13 (.CI(n53435), .I0(n2947), .I1(n2144), .CO(n53436));
    SB_LUT4 add_2756_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n53434), 
            .O(n8267[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_12 (.CI(n53434), .I0(n2948), .I1(n2013), .CO(n53435));
    SB_LUT4 add_2756_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n53433), 
            .O(n8267[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_11 (.CI(n53433), .I0(n2949), .I1(n1879), .CO(n53434));
    SB_LUT4 add_2756_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n53432), 
            .O(n8267[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_10 (.CI(n53432), .I0(n2950), .I1(n1742), .CO(n53433));
    SB_LUT4 add_2756_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n53431), 
            .O(n8267[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_9 (.CI(n53431), .I0(n2951), .I1(n1602), .CO(n53432));
    SB_LUT4 add_2756_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n53430), 
            .O(n8267[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_8 (.CI(n53430), .I0(n2952), .I1(n1459), .CO(n53431));
    SB_LUT4 add_2756_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n53429), 
            .O(n8267[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_7 (.CI(n53429), .I0(n2953), .I1(n1460), .CO(n53430));
    SB_LUT4 add_2756_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n53428), 
            .O(n8267[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_6 (.CI(n53428), .I0(n2954), .I1(n1011), .CO(n53429));
    SB_LUT4 add_2756_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n53427), 
            .O(n8267[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_5 (.CI(n53427), .I0(n2955), .I1(n856), .CO(n53428));
    SB_LUT4 add_2756_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n53426), 
            .O(n8267[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8085[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2756_4 (.CI(n53426), .I0(n2956), .I1(n698), .CO(n53427));
    SB_LUT4 add_2756_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n53425), 
            .O(n8267[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_3 (.CI(n53425), .I0(n2957), .I1(n858), .CO(n53426));
    SB_LUT4 add_2756_2_lut (.I0(n61258), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2756_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53425));
    SB_LUT4 add_2755_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n53424), 
            .O(n8241[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2755_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n53423), 
            .O(n8241[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_20 (.CI(n53423), .I0(n2828), .I1(n2977), .CO(n53424));
    SB_LUT4 add_2755_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n53422), 
            .O(n8241[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_19 (.CI(n53422), .I0(n2829), .I1(n2867), .CO(n53423));
    SB_LUT4 add_2755_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n53421), 
            .O(n8241[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_18 (.CI(n53421), .I0(n2830), .I1(n2754), .CO(n53422));
    SB_LUT4 add_2755_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n53420), 
            .O(n8241[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_17 (.CI(n53420), .I0(n2831), .I1(n2638), .CO(n53421));
    SB_LUT4 add_2755_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n53419), 
            .O(n8241[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_16 (.CI(n53419), .I0(n2832), .I1(n2519), .CO(n53420));
    SB_LUT4 i1_3_lut_adj_1019 (.I0(n27975), .I1(n48_adj_5144), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1019.LUT_INIT = 16'hefef;
    SB_LUT4 add_2755_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n53418), 
            .O(n8241[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_15 (.CI(n53418), .I0(n2833), .I1(n2397), .CO(n53419));
    SB_LUT4 add_2755_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n53417), 
            .O(n8241[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_14 (.CI(n53417), .I0(n2834), .I1(n2272), .CO(n53418));
    SB_LUT4 add_2755_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n53416), 
            .O(n8241[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_13 (.CI(n53416), .I0(n2835), .I1(n2144), .CO(n53417));
    SB_LUT4 add_2755_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n53415), 
            .O(n8241[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_12 (.CI(n53415), .I0(n2836), .I1(n2013), .CO(n53416));
    SB_LUT4 add_2755_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n53414), 
            .O(n8241[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_11 (.CI(n53414), .I0(n2837), .I1(n1879), .CO(n53415));
    SB_LUT4 add_2755_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n53413), 
            .O(n8241[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_10 (.CI(n53413), .I0(n2838), .I1(n1742), .CO(n53414));
    SB_LUT4 add_2755_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n53412), 
            .O(n8241[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_9 (.CI(n53412), .I0(n2839), .I1(n1602), .CO(n53413));
    SB_LUT4 add_2755_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n53411), 
            .O(n8241[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_8 (.CI(n53411), .I0(n2840), .I1(n1459), .CO(n53412));
    SB_LUT4 add_2755_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n53410), 
            .O(n8241[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_7 (.CI(n53410), .I0(n2841), .I1(n1460), .CO(n53411));
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5192), .I1(baudrate[4]), 
            .I2(n41_adj_5190), .I3(GND_net), .O(n40_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51246_4_lut (.I0(n40_adj_5193), .I1(n36_adj_5191), .I2(n41_adj_5190), 
            .I3(n67837), .O(n70741));   // verilog/uart_rx.v(119[33:55])
    defparam i51246_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51247_3_lut (.I0(n70741), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n70742));   // verilog/uart_rx.v(119[33:55])
    defparam i51247_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(n63965), .I1(n63873), .I2(n63961), 
            .I3(baudrate[19]), .O(n63697));
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2755_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n53409), 
            .O(n8241[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1021 (.I0(n63697), .I1(n63923), .I2(n63967), 
            .I3(n63925), .O(n27990));
    defparam i1_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i41818_1_lut (.I0(n27990), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61266));
    defparam i41818_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2755_6 (.CI(n53409), .I0(n2842), .I1(n1011), .CO(n53410));
    SB_LUT4 add_2755_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n53408), 
            .O(n8241[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_5 (.CI(n53408), .I0(n2843), .I1(n856), .CO(n53409));
    SB_LUT4 i51140_3_lut (.I0(n70742), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n70635));   // verilog/uart_rx.v(119[33:55])
    defparam i51140_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2755_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n53407), 
            .O(n8241[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_4 (.CI(n53407), .I0(n2844), .I1(n698), .CO(n53408));
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7955[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7981[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8007[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8033[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8059[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8033[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8059[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8085[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8085[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n63971));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n63713));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49191_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i49191_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5201), .I1(baudrate[9]), 
            .I2(n35_adj_5143), .I3(GND_net), .O(n32_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7903[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7929[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7955[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7981[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8007[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45042_1_lut (.I0(n64527), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61258));
    defparam i45042_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5206), .I1(baudrate[4]), 
            .I2(n43_adj_5194), .I3(GND_net), .O(n42_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51013_4_lut (.I0(n42_adj_5207), .I1(n38_adj_5205), .I2(n43_adj_5194), 
            .I3(n67845), .O(n70508));   // verilog/uart_rx.v(119[33:55])
    defparam i51013_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51014_3_lut (.I0(n70508), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n70509));   // verilog/uart_rx.v(119[33:55])
    defparam i51014_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51149_4_lut (.I0(n32_adj_5202), .I1(n22_adj_5208), .I2(n35_adj_5143), 
            .I3(n68630), .O(n70644));   // verilog/uart_rx.v(119[33:55])
    defparam i51149_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7929[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7955[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7981[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51150_3_lut (.I0(n70644), .I1(baudrate[10]), .I2(n37_adj_5142), 
            .I3(GND_net), .O(n70645));   // verilog/uart_rx.v(119[33:55])
    defparam i51150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8007[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50992_3_lut (.I0(n70645), .I1(baudrate[11]), .I2(n39_adj_5141), 
            .I3(GND_net), .O(n70487));   // verilog/uart_rx.v(119[33:55])
    defparam i50992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50867_4_lut (.I0(n39_adj_5141), .I1(n37_adj_5142), .I2(n35_adj_5143), 
            .I3(n68632), .O(n70362));
    defparam i50867_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49298_4_lut (.I0(n35_adj_5209), .I1(n33_adj_5195), .I2(n31_adj_5196), 
            .I3(n29_adj_5211), .O(n68793));
    defparam i49298_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5212));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5230), 
            .O(n15_adj_5213));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5213), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5212), 
            .I3(n60086), .O(n71751));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i51248_4_lut (.I0(n28_adj_5189), .I1(n20_adj_5214), .I2(n31_adj_5145), 
            .I3(n68635), .O(n70743));   // verilog/uart_rx.v(119[33:55])
    defparam i51248_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5215), .I1(baudrate[9]), 
            .I2(n43_adj_5200), .I3(GND_net), .O(n40_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n63701));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n63705));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n63707));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n63709));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'heeee;
    SB_LUT4 i44975_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n64461));
    defparam i44975_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i45041_4_lut (.I0(n64461), .I1(n63965), .I2(n64459), .I3(n63919), 
            .O(n64527));
    defparam i45041_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i44899_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n64385));
    defparam i44899_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50700_3_lut (.I0(n28_adj_5217), .I1(baudrate[5]), .I2(n35_adj_5209), 
            .I3(GND_net), .O(n70195));   // verilog/uart_rx.v(119[33:55])
    defparam i50700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50701_3_lut (.I0(n70195), .I1(baudrate[6]), .I2(n37_adj_5210), 
            .I3(GND_net), .O(n70196));   // verilog/uart_rx.v(119[33:55])
    defparam i50701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n64383));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'heeee;
    SB_LUT4 i49667_3_lut (.I0(n70487), .I1(baudrate[12]), .I2(n41_adj_5140), 
            .I3(GND_net), .O(n69162));   // verilog/uart_rx.v(119[33:55])
    defparam i49667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45031_4_lut (.I0(n63707), .I1(n63703), .I2(n63705), .I3(n63701), 
            .O(n64517));
    defparam i45031_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51341_4_lut (.I0(n69162), .I1(n70743), .I2(n41_adj_5140), 
            .I3(n70362), .O(n70836));   // verilog/uart_rx.v(119[33:55])
    defparam i51341_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51342_3_lut (.I0(n70836), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n70837));   // verilog/uart_rx.v(119[33:55])
    defparam i51342_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49291_4_lut (.I0(n41_adj_5204), .I1(n39_adj_5203), .I2(n37_adj_5210), 
            .I3(n68793), .O(n68786));
    defparam i49291_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51137_4_lut (.I0(n40_adj_5216), .I1(n30_adj_5218), .I2(n43_adj_5200), 
            .I3(n68784), .O(n70632));   // verilog/uart_rx.v(119[33:55])
    defparam i51137_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49641_3_lut (.I0(n70196), .I1(baudrate[7]), .I2(n39_adj_5203), 
            .I3(GND_net), .O(n69136));   // verilog/uart_rx.v(119[33:55])
    defparam i49641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51285_3_lut (.I0(n70837), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n70780));   // verilog/uart_rx.v(119[33:55])
    defparam i51285_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51339_4_lut (.I0(n69136), .I1(n70632), .I2(n43_adj_5200), 
            .I3(n68786), .O(n70834));   // verilog/uart_rx.v(119[33:55])
    defparam i51339_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_adj_1029 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n63911));
    defparam i1_2_lut_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1030 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n63909));
    defparam i1_2_lut_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 i41806_1_lut (.I0(n27999), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61254));
    defparam i41806_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51340_3_lut (.I0(n70834), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n70835));   // verilog/uart_rx.v(119[33:55])
    defparam i51340_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48856_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n68351));
    defparam i48856_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51212_3_lut (.I0(n70780), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam i51212_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48821_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n68316));
    defparam i48821_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i4200_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9789));   // verilog/uart_rx.v(119[33:55])
    defparam i4200_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i4194_2_lut_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), 
            .I3(GND_net), .O(n40_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam i4194_2_lut_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48916_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n68411));
    defparam i48916_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45047_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n64529), 
            .I3(GND_net), .O(n64533));
    defparam i45047_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8111[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4031_2_lut_3_lut (.I0(n24096), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam i4031_2_lut_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48886_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n68381));
    defparam i48886_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49213_2_lut_3_lut (.I0(n27896), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n67662));   // verilog/uart_rx.v(119[33:55])
    defparam i49213_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_4_lut_adj_1031 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n63981));
    defparam i1_2_lut_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1032 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n63941));
    defparam i1_2_lut_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8059[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44973_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[29]), .O(n64459));
    defparam i44973_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n63883));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4209_2_lut_4_lut (.I0(n960), .I1(n9789), .I2(n24122), .I3(baudrate[3]), 
            .O(n44_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam i4209_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n63703));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'heeee;
    SB_LUT4 i4207_2_lut_3_lut (.I0(baudrate[3]), .I1(n24122), .I2(n9789), 
            .I3(GND_net), .O(n9796));   // verilog/uart_rx.v(119[33:55])
    defparam i4207_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i4038_2_lut_4_lut (.I0(n804), .I1(n40931), .I2(n24096), .I3(baudrate[2]), 
            .O(n44_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam i4038_2_lut_4_lut.LUT_INIT = 16'ha2fb;
    SB_LUT4 i1_3_lut_4_lut_adj_1034 (.I0(n27896), .I1(n48_adj_5077), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5231));
    defparam i1_3_lut_4_lut_adj_1034.LUT_INIT = 16'hefff;
    SB_LUT4 i48543_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5077), .I2(n27896), 
            .I3(GND_net), .O(n68038));   // verilog/uart_rx.v(119[33:55])
    defparam i48543_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48746_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n68241));
    defparam i48746_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i6245_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n24096));   // verilog/uart_rx.v(119[33:55])
    defparam i6245_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48791_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n68286));
    defparam i48791_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i45018_1_lut_2_lut (.I0(baudrate[12]), .I1(n64467), .I2(GND_net), 
            .I3(GND_net), .O(n61291));
    defparam i45018_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 equal_349_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(98[17:39])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45048_1_lut_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), 
            .I2(n64529), .I3(GND_net), .O(n61308));
    defparam i45048_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i49048_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n68543));
    defparam i49048_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45017_2_lut (.I0(baudrate[12]), .I1(n64467), .I2(GND_net), 
            .I3(GND_net), .O(n64503));
    defparam i45017_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8137[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1035 (.I0(n70227), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63145), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1035.LUT_INIT = 16'h7100;
    SB_LUT4 i51500_2_lut_4_lut (.I0(n70227), .I1(baudrate[16]), .I2(n2476), 
            .I3(n64323), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i51500_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8163[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50704_3_lut (.I0(n32_adj_5244), .I1(baudrate[5]), .I2(n39_adj_5242), 
            .I3(GND_net), .O(n70199));   // verilog/uart_rx.v(119[33:55])
    defparam i50704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50705_3_lut (.I0(n70199), .I1(baudrate[6]), .I2(n41_adj_5243), 
            .I3(GND_net), .O(n70200));   // verilog/uart_rx.v(119[33:55])
    defparam i50705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49337_4_lut (.I0(n41_adj_5243), .I1(n39_adj_5242), .I2(n37_adj_5241), 
            .I3(n67815), .O(n68832));
    defparam i49337_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49060_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n68555));
    defparam i49060_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i2314_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2314_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5230), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n59798), .O(n63237));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n63237), .O(n63243));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h0100;
    SB_LUT4 i50720_3_lut (.I0(n34_adj_5246), .I1(baudrate[4]), .I2(n37_adj_5241), 
            .I3(GND_net), .O(n70215));   // verilog/uart_rx.v(119[33:55])
    defparam i50720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(n63243), .I1(n6), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n31398));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'h0323;
    SB_LUT4 i1_3_lut_4_lut_adj_1039 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n63057));
    defparam i1_3_lut_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2307_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2307_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45046_1_lut_2_lut (.I0(baudrate[8]), .I1(n64529), .I2(GND_net), 
            .I3(GND_net), .O(n61304));
    defparam i45046_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i49257_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5230), .I3(n60086), .O(n67620));
    defparam i49257_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i49254_4_lut (.I0(n67620), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n67617));
    defparam i49254_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(r_SM_Main[1]), .I1(n67617), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n30080));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i49635_3_lut (.I0(n70200), .I1(baudrate[7]), .I2(n43_adj_5240), 
            .I3(GND_net), .O(n69130));   // verilog/uart_rx.v(119[33:55])
    defparam i49635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i41488_2_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n60927));
    defparam i41488_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51007_4_lut (.I0(n69130), .I1(n70215), .I2(n43_adj_5240), 
            .I3(n68832), .O(n70502));   // verilog/uart_rx.v(119[33:55])
    defparam i51007_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51008_3_lut (.I0(n70502), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n70503));   // verilog/uart_rx.v(119[33:55])
    defparam i51008_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1040 (.I0(n70523), .I1(baudrate[21]), .I2(n3046), 
            .I3(n63155), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1040.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_4_lut_adj_1041 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n63979));
    defparam i1_2_lut_4_lut_adj_1041.LUT_INIT = 16'hfffe;
    SB_LUT4 i51523_2_lut_4_lut (.I0(n70523), .I1(baudrate[21]), .I2(n3046), 
            .I3(n27999), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i51523_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_1042 (.I0(n59798), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main[1]), .O(n63257));
    defparam i1_3_lut_4_lut_adj_1042.LUT_INIT = 16'hfdfc;
    SB_LUT4 i51691_2_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[2]), .O(n30084));
    defparam i51691_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8293[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n63965));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n63967));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n63969));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n70503), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63961));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8007[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8033[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8059[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8085[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n63923));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8267[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8267[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8267[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8267[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i45045_2_lut (.I0(baudrate[8]), .I1(n64529), .I2(GND_net), 
            .I3(GND_net), .O(n64531));
    defparam i45045_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i45044_1_lut (.I0(n64529), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61300));
    defparam i45044_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8267[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8267[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n63921));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'heeee;
    SB_LUT4 i4036_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n24096), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n9625));   // verilog/uart_rx.v(119[33:55])
    defparam i4036_2_lut_3_lut_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8267[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8267[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8267[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(n63979), .I1(n63057), .I2(n63055), 
            .I3(n63969), .O(n27987));
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8267[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22890_rep_4_2_lut (.I0(n7981[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61294));   // verilog/uart_rx.v(119[33:55])
    defparam i22890_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49062_4_lut (.I0(n23_adj_5245), .I1(n21_adj_5104), .I2(n19_adj_5103), 
            .I3(n17_adj_5255), .O(n68557));
    defparam i49062_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49054_4_lut (.I0(n29_adj_5101), .I1(n27_adj_5100), .I2(n25_adj_5248), 
            .I3(n68557), .O(n68549));
    defparam i49054_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_adj_1050 (.I0(n70772), .I1(baudrate[17]), .I2(n2596), 
            .I3(n63147), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1050.LUT_INIT = 16'h7100;
    SB_LUT4 i50855_4_lut (.I0(n35_adj_5099), .I1(n33_adj_5098), .I2(n31_adj_5097), 
            .I3(n68549), .O(n70350));
    defparam i50855_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n61294), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50702_3_lut (.I0(n32_adj_5258), .I1(baudrate[6]), .I2(n39_adj_5197), 
            .I3(GND_net), .O(n70197));   // verilog/uart_rx.v(119[33:55])
    defparam i50702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50670_3_lut (.I0(n16_adj_5259), .I1(baudrate[13]), .I2(n39_adj_5096), 
            .I3(GND_net), .O(n70165));   // verilog/uart_rx.v(119[33:55])
    defparam i50670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8267[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50703_3_lut (.I0(n70197), .I1(baudrate[7]), .I2(n41_adj_5198), 
            .I3(GND_net), .O(n70198));   // verilog/uart_rx.v(119[33:55])
    defparam i50703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50211_4_lut (.I0(n41_adj_5198), .I1(n39_adj_5197), .I2(n37_adj_5199), 
            .I3(n68817), .O(n69706));
    defparam i50211_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50722_3_lut (.I0(n34_adj_5260), .I1(baudrate[5]), .I2(n37_adj_5199), 
            .I3(GND_net), .O(n70217));   // verilog/uart_rx.v(119[33:55])
    defparam i50722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8267[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51511_2_lut_4_lut (.I0(n70710), .I1(baudrate[18]), .I2(n2713), 
            .I3(n27990), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i51511_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1051 (.I0(n70710), .I1(baudrate[18]), .I2(n2713), 
            .I3(n63149), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1051.LUT_INIT = 16'h7100;
    SB_LUT4 i44991_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n64477));
    defparam i44991_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49289_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n68784));
    defparam i49289_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49638_3_lut (.I0(n70198), .I1(baudrate[8]), .I2(n43_adj_5253), 
            .I3(GND_net), .O(n69133));   // verilog/uart_rx.v(119[33:55])
    defparam i49638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i45001_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n64487));
    defparam i45001_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1052 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n63055));
    defparam i1_3_lut_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 i45043_2_lut_3_lut (.I0(n63899), .I1(n64503), .I2(baudrate[9]), 
            .I3(GND_net), .O(n64529));
    defparam i45043_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_adj_1053 (.I0(n63899), .I1(n64503), .I2(n7981[14]), 
            .I3(n48_adj_5249), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1053.LUT_INIT = 16'h0010;
    SB_LUT4 i51005_4_lut (.I0(n69133), .I1(n70217), .I2(n43_adj_5253), 
            .I3(n69706), .O(n70500));   // verilog/uart_rx.v(119[33:55])
    defparam i51005_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51006_3_lut (.I0(n70500), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n70501));   // verilog/uart_rx.v(119[33:55])
    defparam i51006_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50671_3_lut (.I0(n70165), .I1(baudrate[14]), .I2(n41_adj_5095), 
            .I3(GND_net), .O(n70166));   // verilog/uart_rx.v(119[33:55])
    defparam i50671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51480_2_lut_3_lut (.I0(n63899), .I1(n64503), .I2(n48_adj_5249), 
            .I3(GND_net), .O(n294[14]));
    defparam i51480_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i50001_4_lut (.I0(n41_adj_5095), .I1(n39_adj_5096), .I2(n27_adj_5100), 
            .I3(n68555), .O(n69496));
    defparam i50001_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50733_3_lut (.I0(n22_adj_5239), .I1(baudrate[7]), .I2(n27_adj_5100), 
            .I3(GND_net), .O(n70228));   // verilog/uart_rx.v(119[33:55])
    defparam i50733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n70501), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8267[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44993_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n64479));
    defparam i44993_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i49681_3_lut (.I0(n70166), .I1(baudrate[15]), .I2(n43_adj_5043), 
            .I3(GND_net), .O(n69176));   // verilog/uart_rx.v(119[33:55])
    defparam i49681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1054 (.I0(n63965), .I1(n63921), .I2(n63923), 
            .I3(baudrate[11]), .O(n63951));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1055 (.I0(n63951), .I1(n63953), .I2(n63941), 
            .I3(n63897), .O(n27966));
    defparam i1_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8267[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8267[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5238), .I1(baudrate[9]), 
            .I2(n31_adj_5097), .I3(GND_net), .O(n28_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49135_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n68630));
    defparam i49135_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8267[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1056 (.I0(n27966), .I1(n48_adj_5263), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1056.LUT_INIT = 16'hefef;
    SB_LUT4 i51153_4_lut (.I0(n28_adj_5265), .I1(n18_adj_5237), .I2(n31_adj_5097), 
            .I3(n68543), .O(n70648));   // verilog/uart_rx.v(119[33:55])
    defparam i51153_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51154_3_lut (.I0(n70648), .I1(baudrate[10]), .I2(n33_adj_5098), 
            .I3(GND_net), .O(n70649));   // verilog/uart_rx.v(119[33:55])
    defparam i51154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8319[19]), .I3(n294[1]), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8319[20]), .I3(n294[1]), .O(n41_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8319[16]), .I3(n294[1]), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8319[17]), .I3(n294[1]), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8319[18]), .I3(n294[1]), .O(n37_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8267[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8319[14]), .I3(n294[1]), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8319[15]), .I3(n294[1]), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8319[11]), .I3(n294[1]), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8319[12]), .I3(n294[1]), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8319[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8319[22]), .I3(n294[1]), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8319[21]), .I3(n294[1]), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8319[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8319[8]), .I3(n294[1]), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8319[9]), .I3(n294[1]), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8319[10]), .I3(n294[1]), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8319[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8319[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8319[7]), .I3(n294[1]), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8319[13]), .I3(n294[1]), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8033[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63141), .I3(n48_adj_5046), .O(n20_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i49140_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n68635));
    defparam i49140_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50986_3_lut (.I0(n70649), .I1(baudrate[11]), .I2(n35_adj_5099), 
            .I3(GND_net), .O(n70481));   // verilog/uart_rx.v(119[33:55])
    defparam i50986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50009_4_lut (.I0(n41_adj_5095), .I1(n39_adj_5096), .I2(n37), 
            .I3(n70350), .O(n69504));
    defparam i50009_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5223), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8267[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8267[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48757_4_lut (.I0(n31_adj_5269), .I1(n19_adj_5268), .I2(n17_adj_5267), 
            .I3(n15_adj_5266), .O(n68252));
    defparam i48757_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49815_4_lut (.I0(n13_adj_5271), .I1(n11_adj_5270), .I2(n3065), 
            .I3(baudrate[2]), .O(n69310));
    defparam i49815_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50413_4_lut (.I0(n19_adj_5268), .I1(n17_adj_5267), .I2(n15_adj_5266), 
            .I3(n69310), .O(n69908));
    defparam i50413_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(n63621), 
            .I3(GND_net), .O(n63605));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7903[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7929[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1057 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n63549), .I3(GND_net), .O(n63515));
    defparam i1_2_lut_3_lut_adj_1057.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7955[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50407_4_lut (.I0(n25_adj_5262), .I1(n23_adj_5261), .I2(n21_adj_5264), 
            .I3(n69908), .O(n69902));
    defparam i50407_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48759_4_lut (.I0(n31_adj_5269), .I1(n29_adj_5257), .I2(n27_adj_5256), 
            .I3(n69902), .O(n68254));
    defparam i48759_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7981[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49179_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n68674));
    defparam i49179_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8007[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50636_3_lut (.I0(n8_adj_5272), .I1(baudrate[13]), .I2(n31_adj_5269), 
            .I3(GND_net), .O(n70131));   // verilog/uart_rx.v(119[33:55])
    defparam i50636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8033[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50637_3_lut (.I0(n70131), .I1(baudrate[14]), .I2(n33_adj_5252), 
            .I3(GND_net), .O(n70132));   // verilog/uart_rx.v(119[33:55])
    defparam i50637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8059[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1058 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n63549), .I3(GND_net), .O(n63551));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1058.LUT_INIT = 16'hfbfb;
    SB_LUT4 i49187_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n68682));
    defparam i49187_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_adj_1059 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n63621), .I3(GND_net), .O(n63641));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1059.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1060 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n63549), .I3(GND_net), .O(n63587));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1060.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1061 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n63621), .I3(GND_net), .O(n63623));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1061.LUT_INIT = 16'hfdfd;
    SB_LUT4 i49247_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n68742));
    defparam i49247_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i22839_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n40931));
    defparam i22839_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5234), .I1(baudrate[17]), 
            .I2(n39_adj_5251), .I3(GND_net), .O(n34_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1062 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n63475));
    defparam i1_4_lut_adj_1062.LUT_INIT = 16'h0100;
    SB_LUT4 i48748_4_lut (.I0(n37_adj_5254), .I1(n35_adj_5250), .I2(n33_adj_5252), 
            .I3(n68252), .O(n68243));
    defparam i48748_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51173_4_lut (.I0(n34_adj_5273), .I1(n14_adj_5233), .I2(n39_adj_5251), 
            .I3(n68241), .O(n70668));   // verilog/uart_rx.v(119[33:55])
    defparam i51173_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49719_3_lut (.I0(n70132), .I1(baudrate[15]), .I2(n35_adj_5250), 
            .I3(GND_net), .O(n69214));   // verilog/uart_rx.v(119[33:55])
    defparam i49719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44995_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n64481));
    defparam i44995_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51599_2_lut_4_lut (.I0(n70774), .I1(baudrate[13]), .I2(n2098), 
            .I3(n27975), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i51599_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50638_3_lut (.I0(n10_adj_5232), .I1(baudrate[10]), .I2(n25_adj_5262), 
            .I3(GND_net), .O(n70133));   // verilog/uart_rx.v(119[33:55])
    defparam i50638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50639_3_lut (.I0(n70133), .I1(baudrate[11]), .I2(n27_adj_5256), 
            .I3(GND_net), .O(n70134));   // verilog/uart_rx.v(119[33:55])
    defparam i50639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49789_4_lut (.I0(n27_adj_5256), .I1(n25_adj_5262), .I2(n23_adj_5261), 
            .I3(n68286), .O(n69284));
    defparam i49789_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5235), .I1(baudrate[9]), 
            .I2(n23_adj_5261), .I3(GND_net), .O(n20_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49717_3_lut (.I0(n70134), .I1(baudrate[12]), .I2(n29_adj_5257), 
            .I3(GND_net), .O(n69212));   // verilog/uart_rx.v(119[33:55])
    defparam i49717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50777_4_lut (.I0(n37_adj_5254), .I1(n35_adj_5250), .I2(n33_adj_5252), 
            .I3(n68254), .O(n70272));
    defparam i50777_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51351_4_lut (.I0(n69214), .I1(n70668), .I2(n39_adj_5251), 
            .I3(n68243), .O(n70846));   // verilog/uart_rx.v(119[33:55])
    defparam i51351_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50361_4_lut (.I0(n69212), .I1(n20_adj_5274), .I2(n29_adj_5257), 
            .I3(n69284), .O(n69856));   // verilog/uart_rx.v(119[33:55])
    defparam i50361_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51420_4_lut (.I0(n69856), .I1(n70846), .I2(n39_adj_5251), 
            .I3(n70272), .O(n70915));   // verilog/uart_rx.v(119[33:55])
    defparam i51420_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1063 (.I0(n60980), .I1(n63475), .I2(n64063), 
            .I3(baudrate[16]), .O(n63503));
    defparam i1_4_lut_adj_1063.LUT_INIT = 16'h0004;
    SB_LUT4 i51421_3_lut (.I0(n70915), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n70916));   // verilog/uart_rx.v(119[33:55])
    defparam i51421_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51413_3_lut (.I0(n70916), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n70908));   // verilog/uart_rx.v(119[33:55])
    defparam i51413_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51028_3_lut (.I0(n70908), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n70523));   // verilog/uart_rx.v(119[33:55])
    defparam i51028_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i45071_4_lut (.I0(n64481), .I1(n64477), .I2(n64479), .I3(n64383), 
            .O(n64557));
    defparam i45071_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8241[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8241[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8241[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8241[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51439_4_lut (.I0(n64539), .I1(n68038), .I2(n64557), .I3(n63503), 
            .O(n70934));
    defparam i51439_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8241[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8241[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22841_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n40933));
    defparam i22841_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_i535_4_lut (.I0(n70934), .I1(n44_adj_5231), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8241[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1064 (.I0(n70835), .I1(baudrate[11]), .I2(n1831), 
            .I3(n63139), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1064.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51483_2_lut_4_lut (.I0(n70835), .I1(baudrate[11]), .I2(n1831), 
            .I3(n64503), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i51483_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8241[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8241[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8241[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6254_4_lut (.I0(n804), .I1(n40931), .I2(n24096), .I3(baudrate[2]), 
            .O(n24106));   // verilog/uart_rx.v(119[33:55])
    defparam i6254_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8241[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8241[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5230), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6268_4_lut (.I0(n960), .I1(n9789), .I2(n24122), .I3(baudrate[3]), 
            .O(n24124));   // verilog/uart_rx.v(119[33:55])
    defparam i6268_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8241[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8241[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8241[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8241[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5229), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i49101_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n68596));
    defparam i49101_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7903[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5286));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7929[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5287));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7955[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8215[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63143), .I3(n48_adj_5109), .O(n18_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8215[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8215[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8215[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5288));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8215[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5289));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8215[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49211_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n68706));
    defparam i49211_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49111_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n68606));
    defparam i49111_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7981[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51486_2_lut_4_lut (.I0(n70776), .I1(baudrate[12]), .I2(n1966), 
            .I3(n64467), .O(n294[11]));
    defparam i51486_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8007[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5290));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51596_2_lut_4_lut (.I0(n70501), .I1(baudrate[10]), .I2(n1693), 
            .I3(n27966), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i51596_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8215[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5291));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8033[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8215[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8215[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8215[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5292));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5293));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5294));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8215[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8215[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8059[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5295));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(baudrate[24]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n63925));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n63919));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_adj_1067 (.I0(n70509), .I1(baudrate[6]), .I2(n1111), 
            .I3(n63133), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1067.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5296));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8215[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8215[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51466_2_lut_4_lut (.I0(n70509), .I1(baudrate[6]), .I2(n1111), 
            .I3(n64533), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i51466_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8215[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5297));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5298));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5299));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8215[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49322_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n68817));   // verilog/uart_rx.v(119[33:55])
    defparam i49322_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8215[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5300));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n63819));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48320_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n67815));   // verilog/uart_rx.v(119[33:55])
    defparam i48320_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_3_lut_adj_1069 (.I0(n63819), .I1(n63979), .I2(n63941), 
            .I3(GND_net), .O(n27993));
    defparam i1_3_lut_adj_1069.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5301));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5302));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48902_4_lut (.I0(n35_adj_5302), .I1(n23_adj_5299), .I2(n21_adj_5298), 
            .I3(n19_adj_5297), .O(n68397));
    defparam i48902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48350_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n67845));   // verilog/uart_rx.v(119[33:55])
    defparam i48350_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i49931_4_lut (.I0(n17_adj_5296), .I1(n15_adj_5295), .I2(n2844), 
            .I3(baudrate[2]), .O(n69426));
    defparam i49931_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n63841));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'heeee;
    SB_LUT4 i50479_4_lut (.I0(n23_adj_5299), .I1(n21_adj_5298), .I2(n19_adj_5297), 
            .I3(n69426), .O(n69974));
    defparam i50479_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50477_4_lut (.I0(n29_adj_5294), .I1(n27_adj_5293), .I2(n25_adj_5292), 
            .I3(n69974), .O(n69972));
    defparam i50477_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48978_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n68473));
    defparam i48978_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48906_4_lut (.I0(n35_adj_5302), .I1(n33_adj_5301), .I2(n31_adj_5300), 
            .I3(n69972), .O(n68401));
    defparam i48906_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5303));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n67662), .I1(baudrate[2]), 
            .I2(n70934), .I3(n48_adj_5077), .O(n46_adj_5304));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5304), .I1(baudrate[3]), 
            .I2(n60961), .I3(GND_net), .O(n48_adj_5305));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n63841), .I1(n63901), .I2(n63903), 
            .I3(n63899), .O(n63853));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'hfffe;
    SB_LUT4 i41814_1_lut (.I0(n27993), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61262));
    defparam i41814_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50658_3_lut (.I0(n12_adj_5303), .I1(baudrate[13]), .I2(n35_adj_5302), 
            .I3(GND_net), .O(n70153));   // verilog/uart_rx.v(119[33:55])
    defparam i50658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(n63853), .I1(n27993), .I2(n63845), 
            .I3(n63981), .O(n27945));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1073 (.I0(n27945), .I1(n48_adj_5305), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1073.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5228), .I1(baudrate[17]), 
            .I2(n43_adj_5290), .I3(GND_net), .O(n38_adj_5306));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51586_2_lut_4_lut (.I0(n70405), .I1(baudrate[5]), .I2(n60967), 
            .I3(n27951), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i51586_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i51526_2_lut_4_lut (.I0(n70679), .I1(baudrate[22]), .I2(n3151), 
            .I3(n28002), .O(n294[1]));
    defparam i51526_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50659_3_lut (.I0(n70153), .I1(baudrate[14]), .I2(n37_adj_5289), 
            .I3(GND_net), .O(n70154));   // verilog/uart_rx.v(119[33:55])
    defparam i50659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i48549_2_lut (.I0(baudrate[1]), .I1(n294[20]), .I2(GND_net), 
            .I3(GND_net), .O(n68044));   // verilog/uart_rx.v(119[33:55])
    defparam i48549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49194_4_lut (.I0(n27896), .I1(n68044), .I2(n48_adj_5077), 
            .I3(baudrate[0]), .O(n804));
    defparam i49194_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i44839_1_lut_2_lut (.I0(baudrate[17]), .I1(n27987), .I2(GND_net), 
            .I3(GND_net), .O(n61274));
    defparam i44839_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i48890_4_lut (.I0(n41_adj_5291), .I1(n39_adj_5288), .I2(n37_adj_5289), 
            .I3(n68397), .O(n68385));
    defparam i48890_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48936_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n68431));
    defparam i48936_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n63711));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5307));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51009_3_lut (.I0(n42_adj_5307), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n70504));   // verilog/uart_rx.v(119[33:55])
    defparam i51009_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51131_4_lut (.I0(n38_adj_5306), .I1(n18_adj_5227), .I2(n43_adj_5290), 
            .I3(n68381), .O(n70626));   // verilog/uart_rx.v(119[33:55])
    defparam i51131_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51010_3_lut (.I0(n70504), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n70505));   // verilog/uart_rx.v(119[33:55])
    defparam i51010_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50709_3_lut (.I0(n70505), .I1(baudrate[4]), .I2(n60965), 
            .I3(GND_net), .O(n48_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam i50709_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i49701_3_lut (.I0(n70154), .I1(baudrate[15]), .I2(n39_adj_5288), 
            .I3(GND_net), .O(n69196));   // verilog/uart_rx.v(119[33:55])
    defparam i49701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48661_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n68156));
    defparam i48661_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5225), .I1(baudrate[9]), 
            .I2(n27_adj_5293), .I3(GND_net), .O(n24_adj_5308));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51159_4_lut (.I0(n24_adj_5308), .I1(n14_adj_5224), .I2(n27_adj_5293), 
            .I3(n68411), .O(n70654));   // verilog/uart_rx.v(119[33:55])
    defparam i51159_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51160_3_lut (.I0(n70654), .I1(baudrate[10]), .I2(n29_adj_5294), 
            .I3(GND_net), .O(n70655));   // verilog/uart_rx.v(119[33:55])
    defparam i51160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50976_3_lut (.I0(n70655), .I1(baudrate[11]), .I2(n31_adj_5300), 
            .I3(GND_net), .O(n70471));   // verilog/uart_rx.v(119[33:55])
    defparam i50976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50833_4_lut (.I0(n41_adj_5291), .I1(n39_adj_5288), .I2(n37_adj_5289), 
            .I3(n68401), .O(n70328));
    defparam i50833_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51337_4_lut (.I0(n69196), .I1(n70626), .I2(n43_adj_5290), 
            .I3(n68385), .O(n70832));   // verilog/uart_rx.v(119[33:55])
    defparam i51337_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49699_3_lut (.I0(n70471), .I1(baudrate[12]), .I2(n33_adj_5301), 
            .I3(GND_net), .O(n69194));   // verilog/uart_rx.v(119[33:55])
    defparam i49699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51402_4_lut (.I0(n69194), .I1(n70832), .I2(n43_adj_5290), 
            .I3(n70328), .O(n70897));   // verilog/uart_rx.v(119[33:55])
    defparam i51402_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51403_3_lut (.I0(n70897), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n70898));   // verilog/uart_rx.v(119[33:55])
    defparam i51403_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1075 (.I0(n70635), .I1(baudrate[7]), .I2(n1261), 
            .I3(n63135), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1075.LUT_INIT = 16'h7100;
    SB_LUT4 i51474_2_lut_4_lut (.I0(n70635), .I1(baudrate[7]), .I2(n1261), 
            .I3(n64531), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i51474_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51508_2_lut_4_lut (.I0(n70772), .I1(baudrate[17]), .I2(n2596), 
            .I3(n27987), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i51508_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51583_2_lut_4_lut (.I0(n46_adj_5304), .I1(baudrate[3]), .I2(n60961), 
            .I3(n27945), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i51583_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8215[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8241[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48691_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n68186));
    defparam i48691_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8241[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5309));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5310));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48836_4_lut (.I0(n33_adj_5287), .I1(n21_adj_5286), .I2(n19_adj_5285), 
            .I3(n17_adj_5284), .O(n68331));
    defparam i48836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49875_4_lut (.I0(n15_adj_5310), .I1(n13_adj_5309), .I2(n2956), 
            .I3(baudrate[2]), .O(n69370));
    defparam i49875_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i50451_4_lut (.I0(n21_adj_5286), .I1(n19_adj_5285), .I2(n17_adj_5284), 
            .I3(n69370), .O(n69946));
    defparam i50451_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50447_4_lut (.I0(n27_adj_5283), .I1(n25_adj_5282), .I2(n23_adj_5281), 
            .I3(n69946), .O(n69942));
    defparam i50447_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48840_4_lut (.I0(n33_adj_5287), .I1(n31_adj_5280), .I2(n29_adj_5279), 
            .I3(n69942), .O(n68335));
    defparam i48840_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_3_lut_adj_1076 (.I0(baudrate[26]), .I1(baudrate[30]), 
            .I2(baudrate[23]), .I3(GND_net), .O(n64069));
    defparam i1_2_lut_3_lut_adj_1076.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5311));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50652_3_lut (.I0(n10_adj_5311), .I1(baudrate[13]), .I2(n33_adj_5287), 
            .I3(GND_net), .O(n70147));   // verilog/uart_rx.v(119[33:55])
    defparam i50652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6267_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n24122));   // verilog/uart_rx.v(119[33:55])
    defparam i6267_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48342_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n67837));   // verilog/uart_rx.v(119[33:55])
    defparam i48342_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50653_3_lut (.I0(n70147), .I1(baudrate[14]), .I2(n35_adj_5277), 
            .I3(GND_net), .O(n70148));   // verilog/uart_rx.v(119[33:55])
    defparam i50653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_2_lut (.I0(n24122), .I1(n9789), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_5312));   // verilog/uart_rx.v(119[33:55])
    defparam i4202_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5226), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5312), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5222), .I1(baudrate[17]), 
            .I2(n41_adj_5276), .I3(GND_net), .O(n36_adj_5313));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48823_4_lut (.I0(n39_adj_5278), .I1(n37_adj_5275), .I2(n35_adj_5277), 
            .I3(n68331), .O(n68318));
    defparam i48823_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51169_4_lut (.I0(n36_adj_5313), .I1(n16_adj_5221), .I2(n41_adj_5276), 
            .I3(n68316), .O(n70664));   // verilog/uart_rx.v(119[33:55])
    defparam i51169_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49707_3_lut (.I0(n70148), .I1(baudrate[15]), .I2(n37_adj_5275), 
            .I3(GND_net), .O(n69202));   // verilog/uart_rx.v(119[33:55])
    defparam i49707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7903[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7929[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5220), .I1(baudrate[9]), 
            .I2(n25_adj_5282), .I3(GND_net), .O(n22_adj_5314));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51161_4_lut (.I0(n22_adj_5314), .I1(n12_adj_5219), .I2(n25_adj_5282), 
            .I3(n68351), .O(n70656));   // verilog/uart_rx.v(119[33:55])
    defparam i51161_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7955[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7981[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51162_3_lut (.I0(n70656), .I1(baudrate[10]), .I2(n27_adj_5283), 
            .I3(GND_net), .O(n70657));   // verilog/uart_rx.v(119[33:55])
    defparam i51162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1077 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n63845));
    defparam i1_2_lut_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 i50974_3_lut (.I0(n70657), .I1(baudrate[11]), .I2(n29_adj_5279), 
            .I3(GND_net), .O(n70469));   // verilog/uart_rx.v(119[33:55])
    defparam i50974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50821_4_lut (.I0(n39_adj_5278), .I1(n37_adj_5275), .I2(n35_adj_5277), 
            .I3(n68335), .O(n70316));
    defparam i50821_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8007[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8033[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8059[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51349_4_lut (.I0(n69202), .I1(n70664), .I2(n41_adj_5276), 
            .I3(n68318), .O(n70844));   // verilog/uart_rx.v(119[33:55])
    defparam i51349_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49705_3_lut (.I0(n70469), .I1(baudrate[12]), .I2(n31_adj_5280), 
            .I3(GND_net), .O(n69200));   // verilog/uart_rx.v(119[33:55])
    defparam i49705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51418_4_lut (.I0(n69200), .I1(n70844), .I2(n41_adj_5276), 
            .I3(n70316), .O(n70913));   // verilog/uart_rx.v(119[33:55])
    defparam i51418_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51419_3_lut (.I0(n70913), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n70914));   // verilog/uart_rx.v(119[33:55])
    defparam i51419_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51415_3_lut (.I0(n70914), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n70910));   // verilog/uart_rx.v(119[33:55])
    defparam i51415_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8241[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n63901));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n63903));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n63873));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n64065));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'heeee;
    SB_LUT4 i41802_1_lut_4_lut (.I0(n64067), .I1(n64069), .I2(n63921), 
            .I3(n64065), .O(n61250));
    defparam i41802_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1082 (.I0(n63973), .I1(n63969), .I2(n63971), 
            .I3(n63967), .O(n63953));
    defparam i1_4_lut_adj_1082.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8267[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44843_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n27987), .I3(baudrate[15]), .O(n61282));
    defparam i44843_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8293[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1083 (.I0(n64065), .I1(n63883), .I2(n63965), 
            .I3(n63873), .O(n27999));
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'hfffe;
    SB_LUT4 i51492_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n27987), .I3(n48_adj_5109), .O(n294[8]));
    defparam i51492_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i44841_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n27987), .I3(GND_net), .O(n61278));
    defparam i44841_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i22851_rep_5_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n61311));   // verilog/uart_rx.v(119[33:55])
    defparam i22851_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48560_4_lut (.I0(n27_c), .I1(n15), .I2(n13), .I3(n11), 
            .O(n68055));
    defparam i48560_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8189[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8189[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51276_4_lut (.I0(n69174), .I1(n70478), .I2(n43_adj_5043), 
            .I3(n69504), .O(n70771));   // verilog/uart_rx.v(119[33:55])
    defparam i51276_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n61311), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (clk16MHz, GND_net, \state_7__N_3918[0] , ID, baudrate, 
            n31874, n31873, n31872, n31871, n31870, n31869, n31868, 
            n31867, data_ready, data, n30137, scl_enable, VCC_net, 
            scl, sda_enable, n32663, n32651, n32650, n32649, n32645, 
            n32644, n32640, n6720, n32250, n8, \state[0] , \state_7__N_4126[3] , 
            n4, n4_adj_4, n40902, sda_out, n10, n10_adj_5, n27930, 
            n27881, n67782) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    input GND_net;
    input \state_7__N_3918[0] ;
    output [7:0]ID;
    output [31:0]baudrate;
    input n31874;
    input n31873;
    input n31872;
    input n31871;
    input n31870;
    input n31869;
    input n31868;
    input n31867;
    output data_ready;
    output [7:0]data;
    output n30137;
    output scl_enable;
    input VCC_net;
    output scl;
    output sda_enable;
    input n32663;
    input n32651;
    input n32650;
    input n32649;
    input n32645;
    input n32644;
    input n32640;
    output n6720;
    input n32250;
    input n8;
    output \state[0] ;
    input \state_7__N_4126[3] ;
    output n4;
    output n4_adj_4;
    output n40902;
    output sda_out;
    output n10;
    output n10_adj_5;
    output n27930;
    output n27881;
    output n67782;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire enable_slow_N_4213, ready_prev;
    wire [0:0]n5940;
    
    wire enable;
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    wire [7:0]state_7__N_3885;
    
    wire n62647;
    wire [15:0]delay_counter_15__N_3956;
    
    wire n30054;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n50787, n6945, n6947, n6948, n50765, n6949, n6950, n6951, 
        n3;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n40765, n4_c, n5, n27757;
    wire [7:0]state_adj_5042;   // verilog/i2c_controller.v(33[12:17])
    
    wire n67803;
    wire [2:0]n17;
    
    wire n30244, n31664, n31905, n31904, n31903, n31902, n31901, 
        n31900, n31899, n31898, n31897, n31896, n31895, n31894, 
        n31893, n31892, n31891, n31890, n31889, n31888, n31887, 
        n59507, n59503, n59509, n59505, n31882, n31881, n31880, 
        n31879, n31878, n31877, n31876, n31875, n54952;
    wire [15:0]n5406;
    
    wire n52977, n52976, n52975, n52974, n52973, n52972, n50768, 
        n52971, n52970, n52969, n52968, n52967, n52966, n52965, 
        n52964, n52963, n32664, n59501, n59335, rw, n31698, n31697, 
        n28, n26, n27, n25, n54341, n4_adj_5036, n30060, n10_c, 
        n6, n12, n67802;
    wire [7:0]state_7__N_4110;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n41157, n59747, n15, n23973, n50795, n64279;
    
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5940[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n62647), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n30054), 
            .D(delay_counter_15__N_3956[1]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n30054), 
            .D(delay_counter_15__N_3956[2]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n30054), 
            .D(delay_counter_15__N_3956[3]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n30054), 
            .D(n6945), .S(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n30054), 
            .D(delay_counter_15__N_3956[5]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n30054), 
            .D(n6947), .S(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n30054), 
            .D(n6948), .S(n50765));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n30054), 
            .D(n6949), .S(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n30054), 
            .D(n6950), .S(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n30054), .D(n6951), .S(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n30054), .D(delay_counter_15__N_3956[11]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n30054), .D(delay_counter_15__N_3956[12]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n30054), .D(delay_counter_15__N_3956[13]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n30054), .D(delay_counter_15__N_3956[14]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n30054), .D(delay_counter_15__N_3956[15]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(state[0]), .I2(n3), .I3(state[2]), 
            .O(n50787));
    defparam i1_4_lut.LUT_INIT = 16'h0144;
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n3));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i22673_2_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n40765));
    defparam i22673_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_976 (.I0(state[2]), .I1(state[1]), .I2(\state_7__N_3918[0] ), 
            .I3(state[0]), .O(n4_c));
    defparam i1_4_lut_adj_976.LUT_INIT = 16'hbbba;
    SB_LUT4 i49295_4_lut (.I0(n5), .I1(n27757), .I2(state[1]), .I3(state_adj_5042[3]), 
            .O(n67803));
    defparam i49295_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n67803), .I1(n4_c), .I2(n40765), .I3(state[0]), 
            .O(n62647));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_DFFESR byte_counter_2047__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n30244), .D(n17[2]), .R(n31664));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n30244), .D(n17[1]), .R(n31664));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n31905));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n31904));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n31903));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n31902));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n31901));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n31900));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n31899));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n31898));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n31897));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n31896));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n31895));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n31894));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n31893));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n31892));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n31891));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n31890));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n31889));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n31888));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n31887));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n59507));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n59503));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n59509));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n59505));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n31882));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n31881));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n31880));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n31879));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n31878));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n31877));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n31876));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n31875));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n31874));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n31873));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n31872));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n31871));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n31870));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n31869));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n31868));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n31867));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_4_lut_adj_977 (.I0(n3), .I1(state[0]), .I2(state[2]), .I3(state[1]), 
            .O(state_7__N_3885[1]));
    defparam i1_4_lut_adj_977.LUT_INIT = 16'hf31c;
    SB_DFFESR byte_counter_2047__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n30244), .D(n54952), .R(n31664));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n30054), 
            .D(delay_counter_15__N_3956[0]), .R(n50787));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1198_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5406[9]), 
            .I3(n52977), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1198_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5406[9]), 
            .I3(n52976), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_16 (.CI(n52976), .I0(delay_counter[14]), .I1(n5406[9]), 
            .CO(n52977));
    SB_LUT4 add_1198_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5406[9]), 
            .I3(n52975), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_15 (.CI(n52975), .I0(delay_counter[13]), .I1(n5406[9]), 
            .CO(n52976));
    SB_LUT4 add_1198_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5406[9]), 
            .I3(n52974), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_14 (.CI(n52974), .I0(delay_counter[12]), .I1(n5406[9]), 
            .CO(n52975));
    SB_LUT4 add_1198_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5406[9]), 
            .I3(n52973), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_13 (.CI(n52973), .I0(delay_counter[11]), .I1(n5406[9]), 
            .CO(n52974));
    SB_LUT4 add_1198_12_lut (.I0(n50768), .I1(delay_counter[10]), .I2(n5406[9]), 
            .I3(n52972), .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_12 (.CI(n52972), .I0(delay_counter[10]), .I1(n5406[9]), 
            .CO(n52973));
    SB_LUT4 add_1198_11_lut (.I0(n50768), .I1(delay_counter[9]), .I2(n5406[9]), 
            .I3(n52971), .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_11 (.CI(n52971), .I0(delay_counter[9]), .I1(n5406[9]), 
            .CO(n52972));
    SB_LUT4 add_1198_10_lut (.I0(n50768), .I1(delay_counter[8]), .I2(n5406[9]), 
            .I3(n52970), .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_10 (.CI(n52970), .I0(delay_counter[8]), .I1(n5406[9]), 
            .CO(n52971));
    SB_LUT4 add_1198_9_lut (.I0(n50768), .I1(delay_counter[7]), .I2(n5406[9]), 
            .I3(n52969), .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_9 (.CI(n52969), .I0(delay_counter[7]), .I1(n5406[9]), 
            .CO(n52970));
    SB_LUT4 add_1198_8_lut (.I0(n50768), .I1(delay_counter[6]), .I2(n5406[9]), 
            .I3(n52968), .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_8 (.CI(n52968), .I0(delay_counter[6]), .I1(n5406[9]), 
            .CO(n52969));
    SB_LUT4 add_1198_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5406[9]), 
            .I3(n52967), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_7 (.CI(n52967), .I0(delay_counter[5]), .I1(n5406[9]), 
            .CO(n52968));
    SB_LUT4 add_1198_6_lut (.I0(n50768), .I1(delay_counter[4]), .I2(n5406[9]), 
            .I3(n52966), .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_6 (.CI(n52966), .I0(delay_counter[4]), .I1(n5406[9]), 
            .CO(n52967));
    SB_LUT4 add_1198_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5406[9]), 
            .I3(n52965), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_5 (.CI(n52965), .I0(delay_counter[3]), .I1(n5406[9]), 
            .CO(n52966));
    SB_LUT4 add_1198_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5406[9]), 
            .I3(n52964), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_4 (.CI(n52964), .I0(delay_counter[2]), .I1(n5406[9]), 
            .CO(n52965));
    SB_LUT4 add_1198_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5406[9]), 
            .I3(n52963), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_3 (.CI(n52963), .I0(delay_counter[1]), .I1(n5406[9]), 
            .CO(n52964));
    SB_LUT4 add_1198_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5406[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5406[9]), 
            .CO(n52963));
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n32664));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n59501));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n59335));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n31698));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n31697));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n27757));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n27757), .I1(state[0]), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n54341));
    defparam i2_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut (.I0(state[2]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_5036));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i14_4_lut (.I0(n30060), .I1(state[1]), .I2(data_ready), .I3(n4_adj_5036), 
            .O(n31698));   // verilog/eeprom.v(27[11:16])
    defparam i14_4_lut.LUT_INIT = 16'h5072;
    SB_LUT4 i1_4_lut_adj_978 (.I0(state[1]), .I1(rw), .I2(n54341), .I3(state[2]), 
            .O(n10_c));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_978.LUT_INIT = 16'h888a;
    SB_LUT4 i1_4_lut_adj_979 (.I0(n10_c), .I1(rw), .I2(state[0]), .I3(state[2]), 
            .O(n59335));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_979.LUT_INIT = 16'heeae;
    SB_LUT4 i30_4_lut (.I0(\state_7__N_3918[0] ), .I1(n5), .I2(state[1]), 
            .I3(n6), .O(n12));
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12), .I1(n67802), .I2(state[0]), .I3(state[2]), 
            .O(n59501));
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i1_4_lut_adj_980 (.I0(state_7__N_4110[0]), .I1(saved_addr[0]), 
            .I2(rw), .I3(n41157), .O(n59747));   // verilog/i2c_controller.v(34[12:22])
    defparam i1_4_lut_adj_980.LUT_INIT = 16'hcce4;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n54952));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i32717_4_lut_4_lut (.I0(state[1]), .I1(n3), .I2(state[2]), 
            .I3(state[0]), .O(n50765));
    defparam i32717_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i25_4_lut_4_lut (.I0(state[1]), .I1(n3), .I2(state[0]), .I3(state[2]), 
            .O(n30054));
    defparam i25_4_lut_4_lut.LUT_INIT = 16'h015a;
    SB_LUT4 i1_4_lut_adj_981 (.I0(state[1]), .I1(state[0]), .I2(n40765), 
            .I3(state[2]), .O(n32664));
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hee08;
    SB_LUT4 i34489_2_lut_3_lut_4_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i34489_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 i1_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n3), .O(n30060));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(\state_7__N_3918[0] ), 
            .I3(state[2]), .O(n31664));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i34496_3_lut_4_lut (.I0(n40765), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i34496_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i13506_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(ID[0]), .O(n31697));
    defparam i13506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13708_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(ID[7]), .O(n31899));
    defparam i13708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13709_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(ID[6]), .O(n31900));
    defparam i13709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13710_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(ID[5]), .O(n31901));
    defparam i13710_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_2_lut (.I0(state[2]), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n50768));
    defparam i13_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i51505_2_lut (.I0(n27757), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5406[9]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i51505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13711_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(ID[4]), .O(n31902));
    defparam i13711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13712_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(ID[3]), .O(n31903));
    defparam i13712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13713_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(ID[2]), .O(n31904));
    defparam i13713_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13714_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(ID[1]), .O(n31905));
    defparam i13714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(byte_counter[1]), .I1(n23973), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n30137));
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_3_lut_adj_983 (.I0(byte_counter[1]), .I1(n23973), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n15));
    defparam i1_2_lut_3_lut_adj_983.LUT_INIT = 16'hfefe;
    SB_LUT4 i13707_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(baudrate[0]), .O(n31898));   // verilog/eeprom.v(68[25:39])
    defparam i13707_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13706_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(baudrate[1]), .O(n31897));   // verilog/eeprom.v(68[25:39])
    defparam i13706_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13705_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(baudrate[2]), .O(n31896));   // verilog/eeprom.v(68[25:39])
    defparam i13705_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13704_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(baudrate[3]), .O(n31895));   // verilog/eeprom.v(68[25:39])
    defparam i13704_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13703_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(baudrate[4]), .O(n31894));   // verilog/eeprom.v(68[25:39])
    defparam i13703_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13702_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(baudrate[5]), .O(n31893));   // verilog/eeprom.v(68[25:39])
    defparam i13702_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13701_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(baudrate[6]), .O(n31892));   // verilog/eeprom.v(68[25:39])
    defparam i13701_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13700_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(baudrate[7]), .O(n31891));   // verilog/eeprom.v(68[25:39])
    defparam i13700_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13697_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[2]), 
            .I3(baudrate[10]), .O(n31888));   // verilog/eeprom.v(68[25:39])
    defparam i13697_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[5]), 
            .I3(baudrate[13]), .O(n59503));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13699_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[0]), 
            .I3(baudrate[8]), .O(n31890));   // verilog/eeprom.v(68[25:39])
    defparam i13699_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13696_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[3]), 
            .I3(baudrate[11]), .O(n31887));   // verilog/eeprom.v(68[25:39])
    defparam i13696_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_984 (.I0(byte_counter[0]), .I1(n50795), 
            .I2(data[4]), .I3(baudrate[12]), .O(n59507));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_984.LUT_INIT = 16'hfb40;
    SB_LUT4 i13698_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[1]), 
            .I3(baudrate[9]), .O(n31889));   // verilog/eeprom.v(68[25:39])
    defparam i13698_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_985 (.I0(byte_counter[0]), .I1(n50795), 
            .I2(data[6]), .I3(baudrate[14]), .O(n59509));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_985.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_986 (.I0(byte_counter[0]), .I1(n50795), 
            .I2(data[7]), .I3(baudrate[15]), .O(n59505));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_986.LUT_INIT = 16'hfb40;
    SB_LUT4 i13691_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[0]), 
            .I3(baudrate[16]), .O(n31882));   // verilog/eeprom.v(68[25:39])
    defparam i13691_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13690_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[1]), 
            .I3(baudrate[17]), .O(n31881));   // verilog/eeprom.v(68[25:39])
    defparam i13690_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13689_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[2]), 
            .I3(baudrate[18]), .O(n31880));   // verilog/eeprom.v(68[25:39])
    defparam i13689_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13688_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[3]), 
            .I3(baudrate[19]), .O(n31879));   // verilog/eeprom.v(68[25:39])
    defparam i13688_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13687_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[4]), 
            .I3(baudrate[20]), .O(n31878));   // verilog/eeprom.v(68[25:39])
    defparam i13687_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13686_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[5]), 
            .I3(baudrate[21]), .O(n31877));   // verilog/eeprom.v(68[25:39])
    defparam i13686_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13685_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[6]), 
            .I3(baudrate[22]), .O(n31876));   // verilog/eeprom.v(68[25:39])
    defparam i13685_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13684_3_lut_4_lut (.I0(byte_counter[0]), .I1(n50795), .I2(data[7]), 
            .I3(baudrate[23]), .O(n31875));   // verilog/eeprom.v(68[25:39])
    defparam i13684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i49294_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(state[1]), .I3(GND_net), .O(n67802));
    defparam i49294_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i2_3_lut_adj_987 (.I0(n23973), .I1(byte_counter[1]), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n50795));
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h0404;
    SB_LUT4 i44800_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n64279));
    defparam i44800_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(state[2]), .I1(ready_prev), .I2(n41157), .I3(n64279), 
            .O(n23973));
    defparam i4_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mux_1515_Mux_0_i3_3_lut_4_lut (.I0(state[0]), .I1(n27757), .I2(enable_slow_N_4213), 
            .I3(state[1]), .O(n5940[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1515_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h10aa;
    SB_LUT4 i1_4_lut_adj_988 (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(\state_7__N_3918[0] ), .O(n30244));
    defparam i1_4_lut_adj_988.LUT_INIT = 16'h4140;
    i2c_controller i2c (.clk16MHz(clk16MHz), .scl_enable(scl_enable), .GND_net(GND_net), 
            .VCC_net(VCC_net), .\state_7__N_4110[0] (state_7__N_4110[0]), 
            .scl(scl), .sda_enable(sda_enable), .n32663(n32663), .data({data}), 
            .n32651(n32651), .n32650(n32650), .n32649(n32649), .n32645(n32645), 
            .n32644(n32644), .n32640(n32640), .n59747(n59747), .\saved_addr[0] (saved_addr[0]), 
            .n6720(n6720), .\state[3] (state_adj_5042[3]), .n32250(n32250), 
            .n8(n8), .\state[0] (\state[0] ), .enable_slow_N_4213(enable_slow_N_4213), 
            .\state_7__N_4126[3] (\state_7__N_4126[3] ), .enable(enable), 
            .n27757(n27757), .n6(n6), .n5(n5), .n4(n4), .n4_adj_2(n4_adj_4), 
            .n40902(n40902), .sda_out(sda_out), .n10(n10), .n10_adj_3(n10_adj_5), 
            .n27930(n27930), .n27881(n27881), .n67782(n67782), .n41157(n41157)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (clk16MHz, scl_enable, GND_net, VCC_net, \state_7__N_4110[0] , 
            scl, sda_enable, n32663, data, n32651, n32650, n32649, 
            n32645, n32644, n32640, n59747, \saved_addr[0] , n6720, 
            \state[3] , n32250, n8, \state[0] , enable_slow_N_4213, 
            \state_7__N_4126[3] , enable, n27757, n6, n5, n4, n4_adj_2, 
            n40902, sda_out, n10, n10_adj_3, n27930, n27881, n67782, 
            n41157) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input clk16MHz;
    output scl_enable;
    input GND_net;
    input VCC_net;
    output \state_7__N_4110[0] ;
    output scl;
    output sda_enable;
    input n32663;
    output [7:0]data;
    input n32651;
    input n32650;
    input n32649;
    input n32645;
    input n32644;
    input n32640;
    input n59747;
    output \saved_addr[0] ;
    output n6720;
    output \state[3] ;
    input n32250;
    input n8;
    output \state[0] ;
    output enable_slow_N_4213;
    input \state_7__N_4126[3] ;
    input enable;
    input n27757;
    output n6;
    output n5;
    output n4;
    output n4_adj_2;
    output n40902;
    output sda_out;
    output n10;
    output n10_adj_3;
    output n27930;
    output n27881;
    output n67782;
    output n41157;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire i2c_clk_N_4199, scl_enable_N_4200;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n31419;
    wire [5:0]n29;
    
    wire n53685, n53684, n53683, n53682, n53681, enable_slow_N_4212, 
        n30114, n62545, n30108, n59387, n62193, n30106, sda_out_adj_5026;
    wire [7:0]n119;
    
    wire n30163;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n31351, n52984, n52983, n52982, n52981, n52980, n52979, 
        n52978, n5_c;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n40979, n41037, n41214, n62913, n62860, n11, n11_adj_5027, 
        n4_c, n29985, n6713, n11_adj_5028, n40727, n11_adj_5029, 
        n67765, n9, n12, n61130, n28, n70936, n61032;
    wire [1:0]n6789;
    
    wire n11_adj_5035, n15;
    
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n31419));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n31419), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4199));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 counter2_2057_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n53685), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2057_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n53684), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_6 (.CI(n53684), .I0(GND_net), .I1(counter2[4]), 
            .CO(n53685));
    SB_LUT4 counter2_2057_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n53683), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_5 (.CI(n53683), .I0(GND_net), .I1(counter2[3]), 
            .CO(n53684));
    SB_LUT4 counter2_2057_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n53682), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_4 (.CI(n53682), .I0(GND_net), .I1(counter2[2]), 
            .CO(n53683));
    SB_LUT4 counter2_2057_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n53681), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_3 (.CI(n53681), .I0(GND_net), .I1(counter2[1]), 
            .CO(n53682));
    SB_LUT4 counter2_2057_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n53681));
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n30114), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFSR counter2_2057_2058__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i22700_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i22700_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n30108), 
            .D(n62545), .S(n59387));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_5026), .C(i2c_clk), .E(n30106), 
            .D(n62193), .S(n59387));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n30163), .D(n119[0]), 
            .S(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n52984), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n52983), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n52983), .I0(counter[6]), .I1(VCC_net), 
            .CO(n52984));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n52982), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n52982), .I0(counter[5]), .I1(VCC_net), 
            .CO(n52983));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n52981), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n52981), .I0(counter[4]), .I1(VCC_net), 
            .CO(n52982));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n52980), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n52980), .I0(counter[3]), .I1(VCC_net), 
            .CO(n52981));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n52979), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n52979), .I0(counter[2]), .I1(VCC_net), 
            .CO(n52980));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n52978), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n52978), .I0(counter[1]), .I1(VCC_net), 
            .CO(n52979));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n52978));
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n32663));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n32651));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n32650));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n32649));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n32645));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n32644));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n32640));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n59747));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n30163), .D(n119[1]), 
            .S(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n30163), .D(n119[2]), 
            .S(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n30163), .D(n119[3]), 
            .R(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n30163), .D(n119[4]), 
            .R(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n30163), .D(n119[5]), 
            .R(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n30163), .D(n119[6]), 
            .R(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n30163), .D(n119[7]), 
            .R(n31351));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n6720), .D(n5_c), 
            .S(n40979));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(state[2]), .C(i2c_clk), .E(n6720), .D(n41037), 
            .S(n41214));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6720), .D(n62913), 
            .S(n62860));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n32250));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n31419));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i51673_2_lut (.I0(enable_slow_N_4213), .I1(\state_7__N_4110[0] ), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));
    defparam i51673_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut (.I0(\state_7__N_4126[3] ), .I1(n11), .I2(n11_adj_5027), 
            .I3(enable), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'h2a2f;
    SB_LUT4 i51615_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n41037));
    defparam i51615_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i51457_4_lut (.I0(n29985), .I1(n6713), .I2(n11_adj_5028), 
            .I3(n40727), .O(n6720));
    defparam i51457_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n11_adj_5029), .I1(n11), .I2(\state_7__N_4126[3] ), 
            .I3(\saved_addr[0] ), .O(n5_c));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h5755;
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n27757), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(state[1]), .O(n11_adj_5028));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i22778_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(state[2]), 
            .I3(\state[3] ), .O(scl_enable_N_4200));   // verilog/i2c_controller.v(44[32:47])
    defparam i22778_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[2]), .I3(\state[3] ), .O(n11_adj_5029));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i49227_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(n6713), 
            .I3(GND_net), .O(n67765));
    defparam i49227_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 equal_1562_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(state[2]), .I3(\state[3] ), .O(n11_adj_5027));
    defparam equal_1562_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(\state[0] ), 
            .I3(GND_net), .O(n5));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[3] ), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[2]), .O(n62545));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1110;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i22810_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n40902));
    defparam i22810_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2555_2_lut (.I0(sda_out_adj_5026), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_964 (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut_adj_964.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[6]), 
            .I3(counter[5]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[4]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6713));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i41682_3_lut (.I0(state[2]), .I1(\state_7__N_4126[3] ), .I2(state[1]), 
            .I3(GND_net), .O(n61130));
    defparam i41682_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_965 (.I0(\state[3] ), .I1(n67765), .I2(n61130), 
            .I3(\state[0] ), .O(n30163));
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h0544;
    SB_LUT4 i1_4_lut_adj_966 (.I0(\state[3] ), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[2]), .O(n28));
    defparam i1_4_lut_adj_966.LUT_INIT = 16'h5110;
    SB_LUT4 i51441_2_lut (.I0(\state[3] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n70936));
    defparam i51441_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_967 (.I0(n11_adj_5027), .I1(n70936), .I2(n28), 
            .I3(n61032), .O(n30106));
    defparam i1_4_lut_adj_967.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1830_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6789[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1830_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 state_7__I_0_144_i10_2_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i41586_2_lut (.I0(\state[0] ), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n61032));
    defparam i41586_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n11_adj_5027), .I1(n61032), .I2(\state[3] ), 
            .I3(state[1]), .O(n59387));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_968 (.I0(n11_adj_5027), .I1(state[1]), .I2(\state[3] ), 
            .I3(n61032), .O(n30108));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), .I2(state[2]), 
            .I3(\state[3] ), .O(n29985));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(\state[3] ), .I3(state[2]), .O(n11));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i23055_2_lut_3_lut (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n40727));
    defparam i23055_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i51580_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), .I2(state[1]), 
            .I3(n6720), .O(n62860));
    defparam i51580_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_969 (.I0(enable), .I1(enable_slow_N_4213), 
            .I2(\state_7__N_4110[0] ), .I3(GND_net), .O(n30114));
    defparam i1_2_lut_3_lut_adj_969.LUT_INIT = 16'hbaba;
    SB_LUT4 i51588_3_lut_4_lut (.I0(n9), .I1(n10_adj_3), .I2(n11_adj_5035), 
            .I3(n6720), .O(n41214));   // verilog/i2c_controller.v(151[5:14])
    defparam i51588_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut_adj_970 (.I0(n9), .I1(n10_adj_3), .I2(counter[0]), 
            .I3(GND_net), .O(n27930));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_970.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_971 (.I0(n9), .I1(n10_adj_3), .I2(counter[0]), 
            .I3(GND_net), .O(n27881));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_971.LUT_INIT = 16'hefef;
    SB_LUT4 i48756_3_lut_4_lut (.I0(n11_adj_5028), .I1(n11_adj_5035), .I2(enable_slow_N_4213), 
            .I3(\state_7__N_4110[0] ), .O(n67782));
    defparam i48756_3_lut_4_lut.LUT_INIT = 16'h0888;
    SB_LUT4 i51590_3_lut_4_lut (.I0(n11_adj_5028), .I1(n11_adj_5035), .I2(n15), 
            .I3(n6720), .O(n40979));
    defparam i51590_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(state[1]), .I3(\state[0] ), .O(n11_adj_5035));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_972 (.I0(state[2]), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9), .O(n62913));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_972.LUT_INIT = 16'hf0f4;
    SB_LUT4 i51670_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[3] ), 
            .I3(state[2]), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i51670_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_4_lut_adj_973 (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(state[1]), .O(n41157));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_973.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_276_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(\state[3] ), 
            .I2(state[1]), .I3(\state[0] ), .O(n15));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam equal_276_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_974 (.I0(state[2]), .I1(\state[3] ), .I2(n6789[1]), 
            .I3(state[1]), .O(n62193));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_974.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(state[2]), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(n30163), .O(n31351));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'h1000;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_setpoint, GND_net, n2887, pwm_out, clk32MHz, VCC_net, 
            reset) /* synthesis syn_module_defined=1 */ ;
    input [23:0]pwm_setpoint;
    input GND_net;
    input n2887;
    output pwm_out;
    input clk32MHz;
    input VCC_net;
    input reset;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n41, n39, n45, n43, n37, n23, n25, n29, n31, n35, 
        n33, n9, n17, n19, n21, n11, n15, n27, n13, n68322, 
        n68298, n12, n30, n68450, n69442, n69360, n70564, n69912, 
        n70717, n6, n70306, n70307, n16, n24, n68227, n8, n68209, 
        n69772, n68957, n4, n69914, n69915, n68269, n10, n68260, 
        n70674, n68955, n70855, n70856, n70758, n68229, n70432, 
        n70118, n70684, pwm_out_N_577, n4_adj_5022, n62406, n62108, 
        n16_adj_5023, n15_adj_5024, n17_adj_5025, n48, n58445, n53539, 
        n58487, n53538, n58519, n53537, n58559, n53536, n58599, 
        n53535, n58639, n53534, n58673, n53533, n58719, n53532, 
        n58759, n53531, n58797, n53530, n58829, n53529, n58867, 
        n53528, n58905, n53527, n58947, n53526, n58995, n53525, 
        n59039, n53524, n59091, n53523, n59169, n53522, n59311, 
        n53521, n59475, n53520, n59589, n53519, n59587, n53518, 
        n59585, n53517, n59577;
    
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48827_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n68322));
    defparam i48827_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48803_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n68298));
    defparam i48803_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49947_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n68450), 
            .O(n69442));
    defparam i49947_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49865_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n69442), 
            .O(n69360));
    defparam i49865_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51069_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n69360), 
            .O(n70564));
    defparam i51069_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50417_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n70564), 
            .O(n69912));
    defparam i50417_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51222_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69912), 
            .O(n70717));
    defparam i51222_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50811_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n70306));   // verilog/pwm.v(21[8:24])
    defparam i50811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50812_3_lut (.I0(n70306), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n70307));   // verilog/pwm.v(21[8:24])
    defparam i50812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48732_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n68322), 
            .O(n68227));
    defparam i48732_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50277_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n68209), 
            .O(n69772));   // verilog/pwm.v(21[8:24])
    defparam i50277_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49462_3_lut (.I0(n70307), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n68957));   // verilog/pwm.v(21[8:24])
    defparam i49462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50419_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n69914));   // verilog/pwm.v(21[8:24])
    defparam i50419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50420_3_lut (.I0(n69914), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n69915));   // verilog/pwm.v(21[8:24])
    defparam i50420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48774_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n68298), 
            .O(n68269));
    defparam i48774_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51179_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n68260), 
            .O(n70674));   // verilog/pwm.v(21[8:24])
    defparam i51179_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49460_3_lut (.I0(n69915), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n68955));   // verilog/pwm.v(21[8:24])
    defparam i49460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51360_4_lut (.I0(n68955), .I1(n70674), .I2(n35), .I3(n68269), 
            .O(n70855));   // verilog/pwm.v(21[8:24])
    defparam i51360_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51361_3_lut (.I0(n70855), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n70856));   // verilog/pwm.v(21[8:24])
    defparam i51361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51263_3_lut (.I0(n70856), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n70758));   // verilog/pwm.v(21[8:24])
    defparam i51263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48734_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n70717), 
            .O(n68229));
    defparam i48734_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50937_4_lut (.I0(n68957), .I1(n69772), .I2(n45), .I3(n68227), 
            .O(n70432));   // verilog/pwm.v(21[8:24])
    defparam i50937_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50623_3_lut (.I0(n70758), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n70118));   // verilog/pwm.v(21[8:24])
    defparam i50623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51189_4_lut (.I0(n70118), .I1(n70432), .I2(n45), .I3(n68229), 
            .O(n70684));   // verilog/pwm.v(21[8:24])
    defparam i51189_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51190_3_lut (.I0(n70684), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i51190_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2887), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i1_2_lut (.I0(pwm_counter[8]), .I1(pwm_counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5022));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(pwm_counter[11]), .I1(pwm_counter[16]), .I2(pwm_counter[18]), 
            .I3(pwm_counter[19]), .O(n62406));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(pwm_counter[6]), .I1(pwm_counter[10]), .I2(n4_adj_5022), 
            .I3(pwm_counter[9]), .O(n62108));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[21]), .I1(n62108), .I2(n62406), 
            .I3(pwm_counter[12]), .O(n16_adj_5023));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(pwm_counter[17]), .I1(pwm_counter[13]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5024));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[20]), .I2(pwm_counter[15]), 
            .I3(pwm_counter[14]), .O(n17_adj_5025));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n17_adj_5025), .I2(n15_adj_5024), 
            .I3(n16_adj_5023), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_counter_2040_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n53539), .O(n58445)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2040_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n53538), .O(n58487)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_24 (.CI(n53538), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n53539));
    SB_LUT4 pwm_counter_2040_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n53537), .O(n58519)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_23 (.CI(n53537), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n53538));
    SB_LUT4 pwm_counter_2040_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n53536), .O(n58559)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_22 (.CI(n53536), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n53537));
    SB_LUT4 pwm_counter_2040_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n53535), .O(n58599)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_21 (.CI(n53535), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n53536));
    SB_LUT4 pwm_counter_2040_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n53534), .O(n58639)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_20 (.CI(n53534), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n53535));
    SB_LUT4 pwm_counter_2040_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n53533), .O(n58673)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_19 (.CI(n53533), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n53534));
    SB_LUT4 pwm_counter_2040_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n53532), .O(n58719)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_18 (.CI(n53532), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n53533));
    SB_LUT4 pwm_counter_2040_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n53531), .O(n58759)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_17 (.CI(n53531), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n53532));
    SB_LUT4 pwm_counter_2040_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n53530), .O(n58797)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_16 (.CI(n53530), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n53531));
    SB_LUT4 pwm_counter_2040_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n53529), .O(n58829)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_15 (.CI(n53529), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n53530));
    SB_LUT4 pwm_counter_2040_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n53528), .O(n58867)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_14 (.CI(n53528), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n53529));
    SB_LUT4 pwm_counter_2040_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n53527), .O(n58905)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_13 (.CI(n53527), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n53528));
    SB_LUT4 pwm_counter_2040_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n53526), .O(n58947)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_12 (.CI(n53526), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n53527));
    SB_LUT4 pwm_counter_2040_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n53525), .O(n58995)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_11 (.CI(n53525), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n53526));
    SB_LUT4 pwm_counter_2040_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n53524), .O(n59039)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_10 (.CI(n53524), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n53525));
    SB_LUT4 pwm_counter_2040_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n53523), .O(n59091)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_9 (.CI(n53523), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n53524));
    SB_LUT4 pwm_counter_2040_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n53522), .O(n59169)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_8 (.CI(n53522), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n53523));
    SB_LUT4 pwm_counter_2040_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n53521), .O(n59311)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_7 (.CI(n53521), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n53522));
    SB_LUT4 pwm_counter_2040_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n53520), .O(n59475)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_6 (.CI(n53520), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n53521));
    SB_LUT4 pwm_counter_2040_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n53519), .O(n59589)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_5 (.CI(n53519), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n53520));
    SB_LUT4 pwm_counter_2040_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n53518), .O(n59587)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_4 (.CI(n53518), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n53519));
    SB_LUT4 pwm_counter_2040_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n53517), .O(n59585)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_3 (.CI(n53517), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n53518));
    SB_LUT4 pwm_counter_2040_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n59577)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n53517));
    SB_DFFR pwm_counter_2040__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n59577), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n59585), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n59587), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n59589), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n59475), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n59311), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n59169), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n59091), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n59039), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n58995), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n58947), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n58905), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n58867), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n58829), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n58797), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n58759), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n58719), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n58673), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n58639), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n58599), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n58559), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n58519), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n58487), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n58445), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i48955_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n68450));   // verilog/pwm.v(21[8:24])
    defparam i48955_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48714_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n68209));
    defparam i48714_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48765_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n68260));
    defparam i48765_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[4] , n335, GND_net, \Ki[5] , \Ki[6] , \Ki[7] , 
            setpoint, motor_state, IntegralLimit, \Ki[9] , \Kp[8] , 
            \Ki[10] , \Ki[11] , \Ki[8] , \Kp[9] , \Kp[10] , \Ki[1] , 
            \Ki[0] , \Ki[2] , \Ki[3] , \Kp[11] , \Kp[12] , \Kp[13] , 
            \Kp[1] , \Kp[0] , \Ki[12] , \Kp[2] , \Ki[13] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , control_update, duty, clk16MHz, 
            reset, \Kp[7] , \Ki[14] , \Ki[15] , VCC_net, \Kp[14] , 
            \PID_CONTROLLER.integral , n32594, n32593, n32592, n32591, 
            n32590, n32589, n32588, n32587, n32586, n32585, n32584, 
            n32583, n32582, n32581, n32580, n32579, n32578, n32577, 
            n32576, n32575, n32574, n32573, n32570, n31682, \motor_state[23] , 
            \motor_state[22] , \motor_state[21] , \encoder1_position_scaled[0] , 
            n15, n67541, n15_adj_1, \motor_state[20] , \motor_state[19] , 
            \motor_state[18] , \motor_state[17] , \motor_state[16] , \motor_state[15] , 
            \motor_state[14] , \motor_state[13] , \motor_state[12] , \motor_state[11] , 
            \Kp[15] , deadband, PWMLimit, n41195, \control_mode[0] , 
            \control_mode[7] , \control_mode[6] , n62692, \control_mode[1] , 
            n43) /* synthesis syn_module_defined=1 */ ;
    input \Ki[4] ;
    output [23:0]n335;
    input GND_net;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input [23:0]IntegralLimit;
    input \Ki[9] ;
    input \Kp[8] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[12] ;
    input \Kp[2] ;
    input \Ki[13] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input \Kp[7] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input VCC_net;
    input \Kp[14] ;
    output [23:0]\PID_CONTROLLER.integral ;
    input n32594;
    input n32593;
    input n32592;
    input n32591;
    input n32590;
    input n32589;
    input n32588;
    input n32587;
    input n32586;
    input n32585;
    input n32584;
    input n32583;
    input n32582;
    input n32581;
    input n32580;
    input n32579;
    input n32578;
    input n32577;
    input n32576;
    input n32575;
    input n32574;
    input n32573;
    input n32570;
    input n31682;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \encoder1_position_scaled[0] ;
    input n15;
    input n67541;
    input n15_adj_1;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \Kp[15] ;
    input [23:0]deadband;
    input [23:0]PWMLimit;
    output n41195;
    input \control_mode[0] ;
    input \control_mode[7] ;
    input \control_mode[6] ;
    input n62692;
    input \control_mode[1] ;
    input n43;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n314, n53769;
    wire [16:0]n18318;
    
    wire n1111, n53770, n387, n53123;
    wire [16:0]n17992;
    
    wire n673, n53124, n460, n533, n52744, n52745;
    wire [17:0]n17230;
    
    wire n1038, n53768;
    wire [23:0]n207;
    
    wire n52743;
    wire [17:0]n16847;
    
    wire n600, n53122, n52742, n965, n53767, n527, n53121, n52741, 
        n892, n53766;
    wire [23:0]n233;
    
    wire n68528, n6, n819, n53765, n454, n53120, n746, n53764, 
        n676, n673_adj_4430, n53763, n381, n53119, n600_adj_4431, 
        n53762, n527_adj_4432, n53761, n454_adj_4433, n53760, n381_adj_4434, 
        n53759, n615, n749, n822, n606, n688, n761;
    wire [23:0]n285;
    
    wire n284;
    wire [23:0]n310;
    
    wire n258, n104, n35, n177, n250, n679, n752, n308, n53758, 
        n235, n53757, n162, n53756, n20, n89;
    wire [15:0]n19272;
    
    wire n53755, n53754, n1114, n53753, n1041, n53752, n968, n53751, 
        n895, n53750, n822_adj_4435, n53749, n749_adj_4436, n53748, 
        n676_adj_4437, n53747, n603, n53746, n530, n53745, n457, 
        n53744, n384, n53743, n311, n53742, n238, n53741, n165, 
        n53740, n23, n92;
    wire [14:0]n20100;
    
    wire n53739, n1117, n53738, n1044, n53737, n971, n53736, n898, 
        n53735, n825, n53734, n752_adj_4438, n53733, n679_adj_4439, 
        n53732, n606_adj_4440, n53731, n533_adj_4441, n53730, n460_adj_4442, 
        n53729, n308_adj_4443, n53118, n387_adj_4444, n53728, n834, 
        n907, n314_adj_4445, n53727, n980, n235_adj_4446, n53117, 
        n9977, n67775, n4749, n71661, n241, n53726;
    wire [23:0]n535;
    wire [23:0]n455;
    
    wire n71664, n101, n32, n895_adj_4447, n174, n968_adj_4448, 
        n247, n320, n825_adj_4449, n393, n466, n107, n38, n168, 
        n53725, n26, n95;
    wire [13:0]n20810;
    
    wire n1120, n53724, n1047, n53723, n974, n53722, n901, n53721, 
        n828, n53720, n162_adj_4450, n53116, n755, n53719, n682, 
        n53718, n609, n53717, n536_adj_4451, n53716, n463, n53715, 
        n71406, counter_31__N_3714, n390, n53714, n20_adj_4452, n89_adj_4453;
    wire [15:0]n19000;
    
    wire n53115, n317, n53713, n53114, n244, n53712, n67717, n71421, 
        n171, n53711, n29, n98;
    wire [12:0]n21408;
    
    wire n1050, n53710, n977, n53709, n904, n53708, n539, n71424, 
        n1114_adj_4454, n53113, n831, n53707, n67716, n71415, n758, 
        n53706, n685, n53705, n1041_adj_4455, n53112, n612, n53704, 
        n53703, n53702, n180, n53701, n253, n326, n53700, n53699, 
        n53111, n53698, n53110, n399;
    wire [11:0]n21901;
    
    wire n53697, n53696, n472, n53695, n53694, n53693, n53109, 
        n53108, n53692, n71418, n53107, n545, n542, n53691, n469, 
        n53690, n396, n53689, n323_adj_4456, n53688, n603_adj_4457, 
        n53106, n250_adj_4458, n53687, n618, n177_adj_4459, n53686, 
        n530_adj_4460, n53105, n457_adj_4461, n53104, n52740, n67715, 
        n71409, n35_adj_4462, n104_adj_4463, n384_adj_4464, n53103, 
        n691, n764, n837, n910, n122, n323_adj_4466, n53, n195, 
        n268, n396_adj_4467, n125, n341, n414, n487, n56, n311_adj_4469, 
        n53102, n52739, n560, n469_adj_4470, n542_adj_4471, n238_adj_4472, 
        n53101, n615_adj_4473, n198, n898_adj_4474, n165_adj_4475, 
        n53100, n23_adj_4476, n92_adj_4477, n688_adj_4478, n271, n71412;
    wire [8:0]n22816;
    wire [7:0]n22995;
    
    wire n700, n53099, n627, n53098, n761_adj_4479, n52738, n834_adj_4480, 
        n907_adj_4481, n980_adj_4482, n554, n53097, n67714, n71403, 
        n52737;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n53621, n53620, n53619, n344, n53618, n481, n53096, n119, 
        n53617, n50, n53616, n53615, n52736, n192, n53614, n417, 
        n53613;
    wire [3:0]n23323;
    
    wire n6_adj_4483;
    wire [4:0]n23266;
    
    wire n53612, n53611, n971_adj_4484, n53610, n408, n53095, n52735, 
        n53609, n335_c, n53094, n204;
    wire [23:0]motor_state_c;   // verilog/TinyFPGA_B.v(282[22:33])
    wire [5:0]n23217;
    
    wire n62834, n490, n54080;
    wire [4:0]n23287;
    
    wire n417_adj_4485, n54079, n344_adj_4486, n54078, n271_adj_4487, 
        n54077, n262, n53093, n198_adj_4488, n54076, n56_adj_4489, 
        n125_adj_4490;
    wire [8:0]n22739;
    wire [7:0]n22935;
    
    wire n700_adj_4491, n54075, n627_adj_4492, n54074, n554_adj_4493, 
        n54073, n189, n53092, n481_adj_4494, n54072, n408_adj_4495, 
        n54071, n335_adj_4496, n54070, n262_adj_4497, n54069, n189_adj_4498, 
        n54068, n47, n116;
    wire [6:0]n23076;
    
    wire n630, n54067, n1044_adj_4499, n557_adj_4500, n54066, n484, 
        n54065, n411, n54064, n338, n54063, n265, n54062, n192_adj_4501, 
        n54061, n50_adj_4502, n119_adj_4503, n47_adj_4504, n116_adj_4505;
    wire [1:0]n23381;
    
    wire n52428;
    wire [2:0]n23360;
    wire [14:0]n19879;
    
    wire n53091, n131, n62_adj_4506, n1117_adj_4507, n53090, n53089, 
        n53088, n53087;
    wire [5:0]n23185;
    
    wire n53973, n53972, n53971, n53970, n53969, n53968;
    wire [10:0]n22294;
    
    wire n53506, n53505, n53504, n53503, n53502, n53501, n53500, 
        n53499, n53498, n53497, n53496, n53086, n53085, n53084, 
        n53083, n53082, n53081, n53080, n53079, n241_adj_4513, n53078, 
        n490_adj_4514, n64007, n168_adj_4515, n53077, n26_adj_4516, 
        n95_adj_4517;
    wire [13:0]n20618;
    
    wire n1120_adj_4518, n53076, n1047_adj_4519, n53075, n974_adj_4520, 
        n53074, n901_adj_4521, n53073, n828_adj_4522, n53072, n755_adj_4523, 
        n53071, n682_adj_4524, n53070, n609_adj_4525, n53069, n536_adj_4526, 
        n53068, n463_adj_4527, n53067, n390_adj_4528, n53066, n317_adj_4529, 
        n53065, n244_adj_4530, n53064, n171_adj_4531, n53063, n64011, 
        n29_adj_4532, n98_adj_4533;
    wire [12:0]n21243;
    
    wire n1050_adj_4534, n53062, n977_adj_4535, n53061, n904_adj_4536, 
        n53060, n831_adj_4537, n53059, n758_adj_4538, n53058, n685_adj_4539, 
        n53057, n64009, n612_adj_4540, n53056, n539_adj_4541, n53055, 
        n466_adj_4542, n53054, n393_adj_4543, n53053, n320_adj_4544, 
        n53052, n247_adj_4545, n53051, n52398, n64017, n4, n174_adj_4547, 
        n53050, n32_adj_4548, n101_adj_4549, n8;
    wire [6:0]n23121;
    
    wire n630_adj_4550, n53049, n67737, n71547, n6_adj_4552, n62888, 
        n557_adj_4553, n53048, n484_adj_4554, n53047, n71550, n411_adj_4556, 
        n53046, n338_adj_4557, n53045, n265_adj_4558, n53044, n53918, 
        n53917, n53043, n53916;
    wire [11:0]n21761;
    
    wire n53042, n53041, n53040, n53039, n53915, n53038, n53914, 
        n53037, n53036, n53035, n53034, n53033, n53032, n53031;
    wire [0:0]n10676;
    wire [21:0]n11135;
    
    wire n53913;
    wire [43:0]n360;
    
    wire n53912;
    wire [10:0]n22177;
    
    wire n910_adj_4559, n53030, n837_adj_4560, n53029, n764_adj_4561, 
        n53028, n53911, n691_adj_4562, n53027, n53910, n618_adj_4564, 
        n53026;
    wire [9:0]n22597;
    
    wire n840, n53290, n53909, n767, n53289, n545_adj_4565, n53025, 
        n472_adj_4566, n53024, n694, n53288, n399_adj_4567, n53023, 
        n326_adj_4568, n53022, n53908, n621, n53287, n253_adj_4569, 
        n53021, n53907, n180_adj_4571, n53020, n53906, n548, n53286, 
        n38_adj_4572, n107_adj_4573, n560_adj_4574, n53019, n487_adj_4575, 
        n53018, n475, n53285, n414_adj_4576, n53017, n402, n53284, 
        n341_adj_4577, n53016, n1096, n53905, n1023, n53904, n67735, 
        n71541, n329, n53283, n268_adj_4579, n53015, n195_adj_4580, 
        n53014, n950, n53903, n53_adj_4581, n122_adj_4582, n256, 
        n53282, n877, n53902;
    wire [9:0]n22501;
    
    wire n840_adj_4583, n53013, n767_adj_4584, n53012, n694_adj_4585, 
        n53011, n804, n53901, n183, n53281, n41, n110, n621_adj_4587, 
        n53010, n548_adj_4588, n53009, n475_adj_4589, n53008, n731, 
        n53900, n71544, n402_adj_4590, n53007, n329_adj_4591, n53006, 
        n256_adj_4592, n53005, n658, n53899, n183_adj_4593, n53004, 
        n585, n53898, n41_adj_4595, n110_adj_4596, n770, n53003, 
        n512, n53897, n697, n53002, n624, n53001, n551, n53000, 
        n439, n53896, n478_adj_4597, n52999, n405, n52998, n366, 
        n53895, n332, n52997, n293_adj_4599, n53894, n259, n52996, 
        n186, n52995, n44, n113, n220, n53893, n41_adj_4600, n147, 
        n53892, n5, n74_adj_4602, n39;
    wire [0:0]n10017;
    
    wire n52803;
    wire [47:0]n28;
    
    wire n52802, n52801, n71532, n71520, n71514, n71508, n71502, 
        n71496, n71490, n71484, n71478, n71472, n71466, n71460, 
        n71454, n71448, n71442, n71436, n71430, n52800, n52799, 
        n52798, n52797, n52796, n52795, n52794, n52793, n52792, 
        n52791, n52790, n52789, n25, n67734, n71529, n17, n19, 
        n67733, n71517, n23_adj_4609, n67732, n71511, n21, n67731, 
        n71505, n67730, n71499, n43_c, n67729, n71493, n770_adj_4612, 
        n53241;
    wire [20:0]n13103;
    
    wire n53870, n53869, n697_adj_4613, n53240, n53868, n624_adj_4614, 
        n53239, n551_adj_4615, n53238, n478_adj_4616, n53237, n53867, 
        n405_adj_4617, n53236, n332_adj_4618, n53235, n53866, n259_adj_4619, 
        n53234, n186_adj_4620, n53233, n53865, n44_adj_4621, n113_adj_4622, 
        n53864, n1099, n53863, n1026, n53862;
    wire [21:0]n10524;
    
    wire n53232, n53231, n53230, n953, n53861, n53229, n53228, 
        n880, n53860, n53227, n53226, n807, n53859, n53225, n734, 
        n53858, n1096_adj_4623, n53224, n661, n53857, n1023_adj_4624, 
        n53223, n950_adj_4625, n53222, n588, n53856, n877_adj_4626, 
        n53221, n804_adj_4627, n53220, n27, n515, n53855, n442_adj_4629, 
        n53854, n731_adj_4630, n53219, n658_adj_4631, n53218, n52788, 
        n369, n53853, n585_adj_4632, n53217, n512_adj_4633, n53216, 
        n296, n53852, n439_adj_4634, n53215, n52787, n29_adj_4636, 
        n52786, n366_adj_4637, n53214, n293_adj_4638, n53213, n223_adj_4639, 
        n53851, n220_adj_4640, n53212, n147_adj_4641, n53211, n31, 
        n150, n53850, n5_adj_4642, n74_adj_4643, n8_adj_4644, n77;
    wire [20:0]n12531;
    
    wire n53210, n53209;
    wire [23:0]n1_adj_5019;
    
    wire n52949, n52948, n52785;
    wire [19:0]n14630;
    
    wire n53849, n53208, n52947, n52946, n53848, n53207, n52945, 
        n52784, n52944, n53206, n52943, n45, n52783, n52942, n53847, 
        n53846, n52941, n52782, n53205, n52940, n52781, n53845, 
        n52458, n64059, n52939, n53844, n53204, n52938, n52780, 
        n52779;
    wire [3:0]n23335;
    
    wire n4_adj_4652, n347, n6_adj_4653, n60165, n64055, n68_adj_4654, 
        n52937, n1099_adj_4656, n53203, n1026_adj_4657, n53202, n52778, 
        n1102, n53843, n67728, n71487, n953_adj_4658, n53201, n52936, 
        n52935, n52777, n880_adj_4659, n53200, n52934, n52776, n1029, 
        n53842, n52933, n52775, n807_adj_4662, n53199, n52932, n52774, 
        n956, n53841, n734_adj_4664, n53198, n52931, n52773, n52772, 
        n883, n53840, n52930, n52453, n54083, n810, n53839, n661_adj_4668, 
        n53197, n52929, n52771, n52928, n588_adj_4670, n53196, n52927, 
        n737, n53838, n515_adj_4672, n53195, n47_adj_4673;
    wire [23:0]n1_adj_5020;
    
    wire n52926, n64045, n664, n53837, n71973, n64049, n8_adj_4675, 
        n442_adj_4676, n53194;
    wire [23:0]n34;
    
    wire n52925, n6_adj_4678, n591, n53836, n52924, n369_adj_4681, 
        n53193, n52770, n52923, n518, n53835, n33, n52922, n445_adj_4684, 
        n53834, n296_adj_4685, n53192, n52921, n52769, n372, n53833, 
        n52920, n223_adj_4689, n53191, n52919, n299_adj_4691, n53832, 
        n52918, n150_adj_4694, n53190, n52917, n226_adj_4696, n53831, 
        n8_adj_4697, n77_adj_4698, n52916, n52915, n52768, n153, 
        n53830;
    wire [19:0]n14124;
    
    wire n53189, n52914, n53188, n52913, n53187, n52912, n52767, 
        n11_adj_4704, n80, n52766, n52911, n52910, n52765, n53186, 
        n52909, n52764, n52908, n53185, n52763, n52907;
    wire [18:0]n16003;
    
    wire n53829, n53828, n52762, n53827, n53184, n52906, n52761, 
        n53826, n52905, n52760, n1102_adj_4715, n53183, n52904, 
        n52759, n67585, n41203, n52758, n53825, n1029_adj_4719, 
        n53182;
    wire [23:0]n1_adj_5021;
    
    wire n52903, n52902, n52901, n52757, n52756, n1105, n53824, 
        n956_adj_4723, n53181, n52900, n52755, n1032, n53823, n52899, 
        n52754, n959, n53822, n883_adj_4728, n53180, n810_adj_4729, 
        n53179, n886, n53821, n737_adj_4730, n53178, n664_adj_4731, 
        n53177, n813, n53820, n591_adj_4732, n53176, n518_adj_4733, 
        n53175, n740, n53819, n445_adj_4734, n53174, n667, n53818, 
        n594, n53817, n372_adj_4735, n53173, n52898, n52753, n521, 
        n53816, n299_adj_4737, n53172, n448_adj_4738, n53815, n226_adj_4739, 
        n53171, n153_adj_4740, n53170, n375, n53814, n11_adj_4741, 
        n80_adj_4742, n302, n53813;
    wire [18:0]n15560;
    
    wire n53169, n52897, n229, n53812, n53168, n53167, n156, n53811, 
        n53166, n53165, n52896, n14_adj_4745, n83, n1105_adj_4746, 
        n53164, n1032_adj_4747, n53163, n53810, n959_adj_4748, n53162, 
        n53809, n886_adj_4749, n53161, n52895, n53808, n813_adj_4751, 
        n53160, n740_adj_4752, n53159, n53807, n667_adj_4753, n53158, 
        n594_adj_4754, n53157, n1108, n53806, n521_adj_4755, n53156, 
        n1035, n53805, n448_adj_4756, n53155, n375_adj_4757, n53154, 
        n962, n53804, n302_adj_4758, n53153, n229_adj_4759, n53152, 
        n889, n53803, n156_adj_4760, n53151, n52894, n816, n53802, 
        n14_adj_4762, n83_adj_4763, n53150, n53149, n743, n53801, 
        n53148, n670, n53800, n53147, n52893, n1108_adj_4766, n53146, 
        n52892, n597, n53799, n52891, n1035_adj_4769, n53145, n524, 
        n53798, n52890, n962_adj_4771, n53144, n52889, n52888, n451_adj_4774, 
        n53797, n889_adj_4775, n53143, n52887, n52886, n52752, n816_adj_4779, 
        n53142, n52885, n52884, n378, n53796, n743_adj_4782, n53141, 
        n52883, n305_adj_4784, n53795, n232, n53794, n670_adj_4785, 
        n53140, n159, n53793, n52882, n52881, n597_adj_4789, n53139, 
        n17_adj_4790, n86, n524_adj_4792, n53138, n451_adj_4793, n53137, 
        n52751, n378_adj_4794, n53136, n305_adj_4795, n53135, n52750, 
        n52749, n232_adj_4796, n53134, n159_adj_4797, n53133, n52748, 
        n52747, n17_adj_4798, n86_adj_4799, n52746, n53132, n53131, 
        n53130, n35_adj_4800, n1111_adj_4801, n53129, n1038_adj_4802, 
        n53128, n965_adj_4803, n53127, n892_adj_4804, n53126, n819_adj_4805, 
        n53125, n746_adj_4806, n64310, n23_adj_4807, n53772, n53771, 
        n22_adj_4808, n26_adj_4809, n37, n67727, n71481, n9_adj_4810, 
        n68510, n15_adj_4811, n13_adj_4812, n11_adj_4813, n68489, 
        n12_adj_4814, n9_adj_4815, n11_adj_4816, n13_adj_4817, n15_adj_4818, 
        n10_adj_4819, n30, n69514, n41_adj_4820, n39_adj_4821, n45_adj_4822, 
        n43_adj_4823, n69508, n29_adj_4824, n31_adj_4825, n37_adj_4826, 
        n23_adj_4827, n25_adj_4828, n35_adj_4829, n33_adj_4830, n11_adj_4831, 
        n13_adj_4832, n15_adj_4833, n27_adj_4834, n9_adj_4835, n17_adj_4836, 
        n19_adj_4837, n21_adj_4838, n68588, n68576, n12_adj_4839, 
        n10_adj_4840, n30_adj_4841, n68608, n69580, n69572, n70604, 
        n70032, n70737, n16_adj_4842, n6_adj_4843, n70294, n70295, 
        n70596, n8_adj_4844, n24_adj_4845, n68537, n68530, n69794, 
        n70000, n68999, n4_adj_4846, n70290, n70291, n68553, n68551, 
        n70610, n69001, n70818, n68369, n70819, n70805, n68539, 
        n70446, n69007, n70688, n68387, n131_adj_4847, n41_adj_4848, 
        n39_adj_4849, n45_adj_4850, n37_adj_4851, n21_adj_4852, n23_adj_4853, 
        n25_adj_4854, n17_adj_4855, n19_adj_4856, n9_adj_4857, n35_adj_4858, 
        n43_adj_4859, n29_adj_4860, n31_adj_4861, n11_adj_4863, n13_adj_4864, 
        n27_adj_4865, n15_adj_4866, n33_adj_4867, n39_adj_4868, n41_adj_4869, 
        n45_adj_4870, n29_adj_4871, n31_adj_4872, n67878, n43_adj_4873, 
        n37_adj_4874, n23_adj_4875, n25_adj_4876, n35_adj_4877, n33_adj_4878, 
        n9_adj_4879, n17_adj_4880, n67942, n19_adj_4881, n21_adj_4882, 
        n11_adj_4883, n13_adj_4884, n15_adj_4885, n27_adj_4886, n41_adj_4887, 
        n39_adj_4888, n45_adj_4889, n37_adj_4890, n43_adj_4891, n70729, 
        n23_adj_4892, n25_adj_4893, n29_adj_4894, n67726, n71475, 
        n31_adj_4895, n35_adj_4896, n33_adj_4897, n9_adj_4898, n17_adj_4899, 
        n19_adj_4900, n21_adj_4901, n11_adj_4902, n13_adj_4903, n15_adj_4904, 
        n27_adj_4905, n68256, n68235, n12_adj_4906, n10_adj_4907, 
        n30_adj_4908, n68277, n69286, n69278, n8_adj_4909, n70546, 
        n68610, n69884, n70711, n16_adj_4910, n6_adj_4911, n70262, 
        n70263, n8_adj_4912, n24_adj_4913, n68154, n68148, n69802, 
        n16_adj_4914, n69039, n4_adj_4915, n16_adj_4916, n69880, n69881, 
        n68225, n67725, n71469, n68220, n70538, n69041, n70786, 
        n70787, n70714, n10_adj_4917, n68158, n68663, n70454, n69047, 
        n70696, n506, n12_adj_4918, n68343, n68329, n12_adj_4919, 
        n10_adj_4920, n30_adj_4921, n68441, n68365, n69366, n69356, 
        n70570, n69932, n70719, n16_adj_4922, n6_adj_4923, n70268, 
        n70269, n8_adj_4924, n24_adj_4925, n68284, n68279, n69800, 
        n69029, n4_adj_4926, n70266, n68011, n70267, n68320, n68314, 
        n70616, n69031, n70826, n70827, n68040, n70797, n68292, 
        n70452, n69037, n70694, n480, n41_adj_4927, n39_adj_4928, 
        n45_adj_4929, n29_adj_4930, n31_adj_4931, n43_adj_4932, n37_adj_4933, 
        n68435, n6_adj_4934, n23_adj_4935, n25_adj_4936, n35_adj_4937, 
        n33_adj_4938, n11_adj_4939, n13_adj_4940, n15_adj_4941, n70286, 
        n27_adj_4942, n4_adj_4943, n9_adj_4944, n17_adj_4945, n19_adj_4946, 
        n21_adj_4947, n68110, n68088, n12_adj_4949, n10_adj_4950, 
        n30_adj_4951, n68146, n69108, n69102, n70490, n69822, n70702, 
        n16_adj_4952, n6_adj_4953, n69872, n69873, n8_adj_4954, n67724, 
        n71463, n24_adj_4955, n68013, n69804, n69049, n4_adj_4956, 
        n69870, n70287, n69871, n68046, n52562, n70848, n69051, 
        n70903, n70904, n70886, n68017, n70456, n40, n70458, n41_adj_4957, 
        n39_adj_4958, n45_adj_4959, n29_adj_4960, n31_adj_4961, n23_adj_4962, 
        n25_adj_4963, n37_adj_4964, n35_adj_4965, n11_adj_4966, n13_adj_4967, 
        n15_adj_4968, n8_adj_4969, n27_adj_4970, n33_adj_4971, n10_adj_4972, 
        n59791, n67723, n71457, n24_adj_4973, n9_adj_4974, n68444, 
        n69796, n17_adj_4975, n69009, n19_adj_4976, n4_adj_4977, n21_adj_4978, 
        n68712, n70284, n68687, n30_adj_4980, n70285, n68829, n69700, 
        n67722, n71451, n69664, n68475, n70662, n68467, n70612, 
        n69011, n70820, n70821, n70803, n70074, n70749, n6_adj_4981, 
        n70302, n70303, n24_adj_4982, n68620, n69792, n68989, n68448, 
        n4_adj_4984, n70298, n70299, n68676, n70448, n69017, n70608, 
        n68991, n70816, n70817, n70807, n70690, n68624, n70444, 
        n68997, n70686, n105, n7067, n7069, n27766, n62775, n67968, 
        n12_adj_4985, n10_adj_4986, n30_adj_4987, n68003, n68972, 
        n68966, n70438, n27800, n4_adj_4988, n69766, n70682, n6_adj_4989, 
        n70410, n70411, n16_adj_4990, n27764, n8_adj_4991, n24_adj_4992, 
        n4_adj_4993, n67986, n67888, n69806, n70140, n4_adj_4994, 
        n70376, n70377, n67948, n70735, n70142, n70889, n41_adj_4995, 
        n70890, n70843, n67892, n70145, n40_adj_4996, n70462, n62767, 
        n39_adj_4997, n29_adj_4998, n31_adj_4999, n27_adj_5000, n25_adj_5001, 
        n17_adj_5002, n45_adj_5003, n19_adj_5004, n43_adj_5005, n23_adj_5006, 
        n33_adj_5007, n67721, n71445, n35_adj_5008, n37_adj_5009, 
        n21_adj_5010, n68407, n68395, n12_adj_5011, n67718, n67719, 
        n10_adj_5012, n30_adj_5013, n67720, n69432, n69424, n70580, 
        n69964, n70725, n16_adj_5014, n70280, n70281, n8_adj_5015, 
        n24_adj_5016, n68373, n69798, n69019, n4_adj_5017, n70278, 
        n70279, n68391, n70614, n71439, n69021, n70824, n70825, 
        n70799, n68377, n70450, n69027, n70692, n71433, n71427;
    
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_16 (.CI(n53769), .I0(n18318[13]), .I1(n1111), .CO(n53770));
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5140_10 (.CI(n53123), .I0(n17992[7]), .I1(n673), .CO(n53124));
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_12 (.CI(n52744), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n52745));
    SB_LUT4 add_5159_15_lut (.I0(GND_net), .I1(n18318[12]), .I2(n1038), 
            .I3(n53768), .O(n17230[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_15 (.CI(n53768), .I0(n18318[12]), .I1(n1038), .CO(n53769));
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n52743), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_9_lut (.I0(GND_net), .I1(n17992[6]), .I2(n600), .I3(n53122), 
            .O(n16847[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_9 (.CI(n53122), .I0(n17992[6]), .I1(n600), .CO(n53123));
    SB_CARRY sub_15_add_2_11 (.CI(n52743), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n52744));
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n52742), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_10 (.CI(n52742), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n52743));
    SB_LUT4 add_5159_14_lut (.I0(GND_net), .I1(n18318[11]), .I2(n965), 
            .I3(n53767), .O(n17230[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_8_lut (.I0(GND_net), .I1(n17992[5]), .I2(n527), .I3(n53121), 
            .O(n16847[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_8 (.CI(n53121), .I0(n17992[5]), .I1(n527), .CO(n53122));
    SB_CARRY add_5159_14 (.CI(n53767), .I0(n18318[11]), .I1(n965), .CO(n53768));
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n52741), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_13_lut (.I0(GND_net), .I1(n18318[10]), .I2(n892), 
            .I3(n53766), .O(n17230[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49033_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n68528));   // verilog/motorControl.v(56[14:36])
    defparam i49033_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_5159_13 (.CI(n53766), .I0(n18318[10]), .I1(n892), .CO(n53767));
    SB_LUT4 add_5159_12_lut (.I0(GND_net), .I1(n18318[9]), .I2(n819), 
            .I3(n53765), .O(n17230[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_12 (.CI(n53765), .I0(n18318[9]), .I1(n819), .CO(n53766));
    SB_LUT4 add_5140_7_lut (.I0(GND_net), .I1(n17992[4]), .I2(n454), .I3(n53120), 
            .O(n16847[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_11_lut (.I0(GND_net), .I1(n18318[8]), .I2(n746), 
            .I3(n53764), .O(n17230[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_11 (.CI(n53764), .I0(n18318[8]), .I1(n746), .CO(n53765));
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5140_7 (.CI(n53120), .I0(n17992[4]), .I1(n454), .CO(n53121));
    SB_LUT4 add_5159_10_lut (.I0(GND_net), .I1(n18318[7]), .I2(n673_adj_4430), 
            .I3(n53763), .O(n17230[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_10 (.CI(n53763), .I0(n18318[7]), .I1(n673_adj_4430), 
            .CO(n53764));
    SB_LUT4 add_5140_6_lut (.I0(GND_net), .I1(n17992[3]), .I2(n381), .I3(n53119), 
            .O(n16847[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_9_lut (.I0(GND_net), .I1(n18318[6]), .I2(n600_adj_4431), 
            .I3(n53762), .O(n17230[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_9 (.CI(n53762), .I0(n18318[6]), .I1(n600_adj_4431), 
            .CO(n53763));
    SB_LUT4 add_5159_8_lut (.I0(GND_net), .I1(n18318[5]), .I2(n527_adj_4432), 
            .I3(n53761), .O(n17230[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_8 (.CI(n53761), .I0(n18318[5]), .I1(n527_adj_4432), 
            .CO(n53762));
    SB_LUT4 add_5159_7_lut (.I0(GND_net), .I1(n18318[4]), .I2(n454_adj_4433), 
            .I3(n53760), .O(n17230[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_6 (.CI(n53119), .I0(n17992[3]), .I1(n381), .CO(n53120));
    SB_CARRY add_5159_7 (.CI(n53760), .I0(n18318[4]), .I1(n454_adj_4433), 
            .CO(n53761));
    SB_LUT4 add_5159_6_lut (.I0(GND_net), .I1(n18318[3]), .I2(n381_adj_4434), 
            .I3(n53759), .O(n17230[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n335[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_6 (.CI(n53759), .I0(n18318[3]), .I1(n381_adj_4434), 
            .CO(n53760));
    SB_LUT4 add_5159_5_lut (.I0(GND_net), .I1(n18318[2]), .I2(n308), .I3(n53758), 
            .O(n17230[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_5 (.CI(n53758), .I0(n18318[2]), .I1(n308), .CO(n53759));
    SB_LUT4 add_5159_4_lut (.I0(GND_net), .I1(n18318[1]), .I2(n235), .I3(n53757), 
            .O(n17230[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_4 (.CI(n53757), .I0(n18318[1]), .I1(n235), .CO(n53758));
    SB_LUT4 add_5159_3_lut (.I0(GND_net), .I1(n18318[0]), .I2(n162), .I3(n53756), 
            .O(n17230[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_3 (.CI(n53756), .I0(n18318[0]), .I1(n162), .CO(n53757));
    SB_LUT4 add_5159_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n17230[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n53756));
    SB_LUT4 add_5211_18_lut (.I0(GND_net), .I1(n19272[15]), .I2(GND_net), 
            .I3(n53755), .O(n18318[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5211_17_lut (.I0(GND_net), .I1(n19272[14]), .I2(GND_net), 
            .I3(n53754), .O(n18318[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_17 (.CI(n53754), .I0(n19272[14]), .I1(GND_net), 
            .CO(n53755));
    SB_LUT4 add_5211_16_lut (.I0(GND_net), .I1(n19272[13]), .I2(n1114), 
            .I3(n53753), .O(n18318[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_16 (.CI(n53753), .I0(n19272[13]), .I1(n1114), .CO(n53754));
    SB_LUT4 add_5211_15_lut (.I0(GND_net), .I1(n19272[12]), .I2(n1041), 
            .I3(n53752), .O(n18318[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_15 (.CI(n53752), .I0(n19272[12]), .I1(n1041), .CO(n53753));
    SB_LUT4 add_5211_14_lut (.I0(GND_net), .I1(n19272[11]), .I2(n968), 
            .I3(n53751), .O(n18318[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_14 (.CI(n53751), .I0(n19272[11]), .I1(n968), .CO(n53752));
    SB_LUT4 add_5211_13_lut (.I0(GND_net), .I1(n19272[10]), .I2(n895), 
            .I3(n53750), .O(n18318[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_13 (.CI(n53750), .I0(n19272[10]), .I1(n895), .CO(n53751));
    SB_LUT4 add_5211_12_lut (.I0(GND_net), .I1(n19272[9]), .I2(n822_adj_4435), 
            .I3(n53749), .O(n18318[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_12 (.CI(n53749), .I0(n19272[9]), .I1(n822_adj_4435), 
            .CO(n53750));
    SB_LUT4 add_5211_11_lut (.I0(GND_net), .I1(n19272[8]), .I2(n749_adj_4436), 
            .I3(n53748), .O(n18318[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_11 (.CI(n53748), .I0(n19272[8]), .I1(n749_adj_4436), 
            .CO(n53749));
    SB_LUT4 add_5211_10_lut (.I0(GND_net), .I1(n19272[7]), .I2(n676_adj_4437), 
            .I3(n53747), .O(n18318[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_10 (.CI(n53747), .I0(n19272[7]), .I1(n676_adj_4437), 
            .CO(n53748));
    SB_LUT4 add_5211_9_lut (.I0(GND_net), .I1(n19272[6]), .I2(n603), .I3(n53746), 
            .O(n18318[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_9 (.CI(n53746), .I0(n19272[6]), .I1(n603), .CO(n53747));
    SB_LUT4 add_5211_8_lut (.I0(GND_net), .I1(n19272[5]), .I2(n530), .I3(n53745), 
            .O(n18318[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_8 (.CI(n53745), .I0(n19272[5]), .I1(n530), .CO(n53746));
    SB_LUT4 add_5211_7_lut (.I0(GND_net), .I1(n19272[4]), .I2(n457), .I3(n53744), 
            .O(n18318[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_7 (.CI(n53744), .I0(n19272[4]), .I1(n457), .CO(n53745));
    SB_LUT4 add_5211_6_lut (.I0(GND_net), .I1(n19272[3]), .I2(n384), .I3(n53743), 
            .O(n18318[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_6 (.CI(n53743), .I0(n19272[3]), .I1(n384), .CO(n53744));
    SB_LUT4 add_5211_5_lut (.I0(GND_net), .I1(n19272[2]), .I2(n311), .I3(n53742), 
            .O(n18318[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_5 (.CI(n53742), .I0(n19272[2]), .I1(n311), .CO(n53743));
    SB_LUT4 add_5211_4_lut (.I0(GND_net), .I1(n19272[1]), .I2(n238), .I3(n53741), 
            .O(n18318[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_4 (.CI(n53741), .I0(n19272[1]), .I1(n238), .CO(n53742));
    SB_LUT4 add_5211_3_lut (.I0(GND_net), .I1(n19272[0]), .I2(n165), .I3(n53740), 
            .O(n18318[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_3 (.CI(n53740), .I0(n19272[0]), .I1(n165), .CO(n53741));
    SB_LUT4 add_5211_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n18318[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n53740));
    SB_LUT4 add_5258_17_lut (.I0(GND_net), .I1(n20100[14]), .I2(GND_net), 
            .I3(n53739), .O(n19272[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5258_16_lut (.I0(GND_net), .I1(n20100[13]), .I2(n1117), 
            .I3(n53738), .O(n19272[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_16 (.CI(n53738), .I0(n20100[13]), .I1(n1117), .CO(n53739));
    SB_LUT4 add_5258_15_lut (.I0(GND_net), .I1(n20100[12]), .I2(n1044), 
            .I3(n53737), .O(n19272[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_15 (.CI(n53737), .I0(n20100[12]), .I1(n1044), .CO(n53738));
    SB_LUT4 add_5258_14_lut (.I0(GND_net), .I1(n20100[11]), .I2(n971), 
            .I3(n53736), .O(n19272[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_14 (.CI(n53736), .I0(n20100[11]), .I1(n971), .CO(n53737));
    SB_LUT4 add_5258_13_lut (.I0(GND_net), .I1(n20100[10]), .I2(n898), 
            .I3(n53735), .O(n19272[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_13 (.CI(n53735), .I0(n20100[10]), .I1(n898), .CO(n53736));
    SB_LUT4 add_5258_12_lut (.I0(GND_net), .I1(n20100[9]), .I2(n825), 
            .I3(n53734), .O(n19272[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_12 (.CI(n53734), .I0(n20100[9]), .I1(n825), .CO(n53735));
    SB_LUT4 add_5258_11_lut (.I0(GND_net), .I1(n20100[8]), .I2(n752_adj_4438), 
            .I3(n53733), .O(n19272[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_11 (.CI(n53733), .I0(n20100[8]), .I1(n752_adj_4438), 
            .CO(n53734));
    SB_LUT4 add_5258_10_lut (.I0(GND_net), .I1(n20100[7]), .I2(n679_adj_4439), 
            .I3(n53732), .O(n19272[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_10 (.CI(n53732), .I0(n20100[7]), .I1(n679_adj_4439), 
            .CO(n53733));
    SB_LUT4 add_5258_9_lut (.I0(GND_net), .I1(n20100[6]), .I2(n606_adj_4440), 
            .I3(n53731), .O(n19272[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_9 (.CI(n53731), .I0(n20100[6]), .I1(n606_adj_4440), 
            .CO(n53732));
    SB_LUT4 add_5258_8_lut (.I0(GND_net), .I1(n20100[5]), .I2(n533_adj_4441), 
            .I3(n53730), .O(n19272[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_8 (.CI(n53730), .I0(n20100[5]), .I1(n533_adj_4441), 
            .CO(n53731));
    SB_LUT4 add_5258_7_lut (.I0(GND_net), .I1(n20100[4]), .I2(n460_adj_4442), 
            .I3(n53729), .O(n19272[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_5_lut (.I0(GND_net), .I1(n17992[2]), .I2(n308_adj_4443), 
            .I3(n53118), .O(n16847[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_7 (.CI(n53729), .I0(n20100[4]), .I1(n460_adj_4442), 
            .CO(n53730));
    SB_LUT4 add_5258_6_lut (.I0(GND_net), .I1(n20100[3]), .I2(n387_adj_4444), 
            .I3(n53728), .O(n19272[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5258_6 (.CI(n53728), .I0(n20100[3]), .I1(n387_adj_4444), 
            .CO(n53729));
    SB_CARRY add_5140_5 (.CI(n53118), .I0(n17992[2]), .I1(n308_adj_4443), 
            .CO(n53119));
    SB_LUT4 add_5258_5_lut (.I0(GND_net), .I1(n20100[2]), .I2(n314_adj_4445), 
            .I3(n53727), .O(n19272[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5140_4_lut (.I0(GND_net), .I1(n17992[1]), .I2(n235_adj_4446), 
            .I3(n53117), .O(n16847[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_5 (.CI(n53727), .I0(n20100[2]), .I1(n314_adj_4445), 
            .CO(n53728));
    SB_LUT4 n9977_bdd_4_lut (.I0(n9977), .I1(n67775), .I2(setpoint[23]), 
            .I3(n4749), .O(n71661));
    defparam n9977_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5258_4_lut (.I0(GND_net), .I1(n20100[1]), .I2(n241), .I3(n53726), 
            .O(n19272[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71661_bdd_4_lut (.I0(n71661), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4749), .O(n71664));
    defparam n71661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4447));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5258_4 (.CI(n53726), .I0(n20100[1]), .I1(n241), .CO(n53727));
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4448));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4449));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5258_3_lut (.I0(GND_net), .I1(n20100[0]), .I2(n168), .I3(n53725), 
            .O(n19272[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_3 (.CI(n53725), .I0(n20100[0]), .I1(n168), .CO(n53726));
    SB_CARRY add_5140_4 (.CI(n53117), .I0(n17992[1]), .I1(n235_adj_4446), 
            .CO(n53118));
    SB_LUT4 add_5258_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n19272[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5258_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5258_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n53725));
    SB_LUT4 add_5302_16_lut (.I0(GND_net), .I1(n20810[13]), .I2(n1120), 
            .I3(n53724), .O(n20100[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5302_15_lut (.I0(GND_net), .I1(n20810[12]), .I2(n1047), 
            .I3(n53723), .O(n20100[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_15 (.CI(n53723), .I0(n20810[12]), .I1(n1047), .CO(n53724));
    SB_LUT4 add_5302_14_lut (.I0(GND_net), .I1(n20810[11]), .I2(n974), 
            .I3(n53722), .O(n20100[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_14 (.CI(n53722), .I0(n20810[11]), .I1(n974), .CO(n53723));
    SB_LUT4 add_5302_13_lut (.I0(GND_net), .I1(n20810[10]), .I2(n901), 
            .I3(n53721), .O(n20100[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_13 (.CI(n53721), .I0(n20810[10]), .I1(n901), .CO(n53722));
    SB_LUT4 add_5302_12_lut (.I0(GND_net), .I1(n20810[9]), .I2(n828), 
            .I3(n53720), .O(n20100[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_3_lut (.I0(GND_net), .I1(n17992[0]), .I2(n162_adj_4450), 
            .I3(n53116), .O(n16847[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_12 (.CI(n53720), .I0(n20810[9]), .I1(n828), .CO(n53721));
    SB_LUT4 add_5302_11_lut (.I0(GND_net), .I1(n20810[8]), .I2(n755), 
            .I3(n53719), .O(n20100[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_11 (.CI(n53719), .I0(n20810[8]), .I1(n755), .CO(n53720));
    SB_LUT4 add_5302_10_lut (.I0(GND_net), .I1(n20810[7]), .I2(n682), 
            .I3(n53718), .O(n20100[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_10 (.CI(n53718), .I0(n20810[7]), .I1(n682), .CO(n53719));
    SB_LUT4 add_5302_9_lut (.I0(GND_net), .I1(n20810[6]), .I2(n609), .I3(n53717), 
            .O(n20100[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_9 (.CI(n53717), .I0(n20810[6]), .I1(n609), .CO(n53718));
    SB_LUT4 add_5302_8_lut (.I0(GND_net), .I1(n20810[5]), .I2(n536_adj_4451), 
            .I3(n53716), .O(n20100[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_3 (.CI(n53116), .I0(n17992[0]), .I1(n162_adj_4450), 
            .CO(n53117));
    SB_CARRY add_5302_8 (.CI(n53716), .I0(n20810[5]), .I1(n536_adj_4451), 
            .CO(n53717));
    SB_LUT4 add_5302_7_lut (.I0(GND_net), .I1(n20810[4]), .I2(n463), .I3(n53715), 
            .O(n20100[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n71406), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_CARRY add_5302_7 (.CI(n53715), .I0(n20810[4]), .I1(n463), .CO(n53716));
    SB_LUT4 add_5302_6_lut (.I0(GND_net), .I1(n20810[3]), .I2(n390), .I3(n53714), 
            .O(n20100[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_2_lut (.I0(GND_net), .I1(n20_adj_4452), .I2(n89_adj_4453), 
            .I3(GND_net), .O(n16847[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_2 (.CI(GND_net), .I0(n20_adj_4452), .I1(n89_adj_4453), 
            .CO(n53116));
    SB_CARRY add_5302_6 (.CI(n53714), .I0(n20810[3]), .I1(n390), .CO(n53715));
    SB_LUT4 add_5194_18_lut (.I0(GND_net), .I1(n19000[15]), .I2(GND_net), 
            .I3(n53115), .O(n17992[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5302_5_lut (.I0(GND_net), .I1(n20810[2]), .I2(n317), .I3(n53713), 
            .O(n20100[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_5 (.CI(n53713), .I0(n20810[2]), .I1(n317), .CO(n53714));
    SB_LUT4 add_5194_17_lut (.I0(GND_net), .I1(n19000[14]), .I2(GND_net), 
            .I3(n53114), .O(n17992[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5302_4_lut (.I0(GND_net), .I1(n20810[1]), .I2(n244), .I3(n53712), 
            .O(n20100[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_4 (.CI(n53712), .I0(n20810[1]), .I1(n244), .CO(n53713));
    SB_LUT4 n9977_bdd_4_lut_51889 (.I0(n9977), .I1(n67717), .I2(setpoint[3]), 
            .I3(n4749), .O(n71421));
    defparam n9977_bdd_4_lut_51889.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5302_3_lut (.I0(GND_net), .I1(n20810[0]), .I2(n171), .I3(n53711), 
            .O(n20100[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_3 (.CI(n53711), .I0(n20810[0]), .I1(n171), .CO(n53712));
    SB_LUT4 add_5302_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n20100[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5302_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n53711));
    SB_LUT4 add_5341_15_lut (.I0(GND_net), .I1(n21408[12]), .I2(n1050), 
            .I3(n53710), .O(n20810[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_14_lut (.I0(GND_net), .I1(n21408[11]), .I2(n977), 
            .I3(n53709), .O(n20810[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_17 (.CI(n53114), .I0(n19000[14]), .I1(GND_net), 
            .CO(n53115));
    SB_CARRY add_5341_14 (.CI(n53709), .I0(n21408[11]), .I1(n977), .CO(n53710));
    SB_LUT4 add_5341_13_lut (.I0(GND_net), .I1(n21408[10]), .I2(n904), 
            .I3(n53708), .O(n20810[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71421_bdd_4_lut (.I0(n71421), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4749), .O(n71424));
    defparam n71421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_5341_13 (.CI(n53708), .I0(n21408[10]), .I1(n904), .CO(n53709));
    SB_LUT4 add_5194_16_lut (.I0(GND_net), .I1(n19000[13]), .I2(n1114_adj_4454), 
            .I3(n53113), .O(n17992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_12_lut (.I0(GND_net), .I1(n21408[9]), .I2(n831), 
            .I3(n53707), .O(n20810[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9977_bdd_4_lut_51884 (.I0(n9977), .I1(n67716), .I2(setpoint[2]), 
            .I3(n4749), .O(n71415));
    defparam n9977_bdd_4_lut_51884.LUT_INIT = 16'he4aa;
    SB_CARRY add_5341_12 (.CI(n53707), .I0(n21408[9]), .I1(n831), .CO(n53708));
    SB_LUT4 add_5341_11_lut (.I0(GND_net), .I1(n21408[8]), .I2(n758), 
            .I3(n53706), .O(n20810[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_11 (.CI(n53706), .I0(n21408[8]), .I1(n758), .CO(n53707));
    SB_LUT4 add_5341_10_lut (.I0(GND_net), .I1(n21408[7]), .I2(n685), 
            .I3(n53705), .O(n20810[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_16 (.CI(n53113), .I0(n19000[13]), .I1(n1114_adj_4454), 
            .CO(n53114));
    SB_CARRY add_5341_10 (.CI(n53705), .I0(n21408[7]), .I1(n685), .CO(n53706));
    SB_LUT4 add_5194_15_lut (.I0(GND_net), .I1(n19000[12]), .I2(n1041_adj_4455), 
            .I3(n53112), .O(n17992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_9_lut (.I0(GND_net), .I1(n21408[6]), .I2(n612), .I3(n53704), 
            .O(n20810[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_9 (.CI(n53704), .I0(n21408[6]), .I1(n612), .CO(n53705));
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5341_8_lut (.I0(GND_net), .I1(n21408[5]), .I2(n539), .I3(n53703), 
            .O(n20810[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4455));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5341_8 (.CI(n53703), .I0(n21408[5]), .I1(n539), .CO(n53704));
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5341_7_lut (.I0(GND_net), .I1(n21408[4]), .I2(n466), .I3(n53702), 
            .O(n20810[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_7 (.CI(n53702), .I0(n21408[4]), .I1(n466), .CO(n53703));
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5341_6_lut (.I0(GND_net), .I1(n21408[3]), .I2(n393), .I3(n53701), 
            .O(n20810[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_6 (.CI(n53701), .I0(n21408[3]), .I1(n393), .CO(n53702));
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5341_5_lut (.I0(GND_net), .I1(n21408[2]), .I2(n320), .I3(n53700), 
            .O(n20810[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_5 (.CI(n53700), .I0(n21408[2]), .I1(n320), .CO(n53701));
    SB_LUT4 add_5341_4_lut (.I0(GND_net), .I1(n21408[1]), .I2(n247), .I3(n53699), 
            .O(n20810[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_4 (.CI(n53699), .I0(n21408[1]), .I1(n247), .CO(n53700));
    SB_CARRY add_5194_15 (.CI(n53112), .I0(n19000[12]), .I1(n1041_adj_4455), 
            .CO(n53113));
    SB_LUT4 add_5194_14_lut (.I0(GND_net), .I1(n19000[11]), .I2(n968_adj_4448), 
            .I3(n53111), .O(n17992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5341_3_lut (.I0(GND_net), .I1(n21408[0]), .I2(n174), .I3(n53698), 
            .O(n20810[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_14 (.CI(n53111), .I0(n19000[11]), .I1(n968_adj_4448), 
            .CO(n53112));
    SB_LUT4 add_5194_13_lut (.I0(GND_net), .I1(n19000[10]), .I2(n895_adj_4447), 
            .I3(n53110), .O(n17992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5341_3 (.CI(n53698), .I0(n21408[0]), .I1(n174), .CO(n53699));
    SB_LUT4 add_5341_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n20810[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5341_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5341_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n53698));
    SB_LUT4 add_5377_14_lut (.I0(GND_net), .I1(n21901[11]), .I2(n980), 
            .I3(n53697), .O(n21408[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_13_lut (.I0(GND_net), .I1(n21901[10]), .I2(n907), 
            .I3(n53696), .O(n21408[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_13 (.CI(n53696), .I0(n21901[10]), .I1(n907), .CO(n53697));
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5377_12_lut (.I0(GND_net), .I1(n21901[9]), .I2(n834), 
            .I3(n53695), .O(n21408[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_12 (.CI(n53695), .I0(n21901[9]), .I1(n834), .CO(n53696));
    SB_LUT4 add_5377_11_lut (.I0(GND_net), .I1(n21901[8]), .I2(n761), 
            .I3(n53694), .O(n21408[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_11 (.CI(n53694), .I0(n21901[8]), .I1(n761), .CO(n53695));
    SB_CARRY add_5194_13 (.CI(n53110), .I0(n19000[10]), .I1(n895_adj_4447), 
            .CO(n53111));
    SB_LUT4 add_5377_10_lut (.I0(GND_net), .I1(n21901[7]), .I2(n688), 
            .I3(n53693), .O(n21408[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5194_12_lut (.I0(GND_net), .I1(n19000[9]), .I2(n822), 
            .I3(n53109), .O(n17992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_12 (.CI(n53109), .I0(n19000[9]), .I1(n822), .CO(n53110));
    SB_LUT4 add_5194_11_lut (.I0(GND_net), .I1(n19000[8]), .I2(n749), 
            .I3(n53108), .O(n17992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_10 (.CI(n53693), .I0(n21901[7]), .I1(n688), .CO(n53694));
    SB_CARRY add_5194_11 (.CI(n53108), .I0(n19000[8]), .I1(n749), .CO(n53109));
    SB_LUT4 add_5377_9_lut (.I0(GND_net), .I1(n21901[6]), .I2(n615), .I3(n53692), 
            .O(n21408[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71415_bdd_4_lut (.I0(n71415), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4749), .O(n71418));
    defparam n71415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5194_10_lut (.I0(GND_net), .I1(n19000[7]), .I2(n676), 
            .I3(n53107), .O(n17992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_9 (.CI(n53692), .I0(n21901[6]), .I1(n615), .CO(n53693));
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5377_8_lut (.I0(GND_net), .I1(n21901[5]), .I2(n542), .I3(n53691), 
            .O(n21408[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_8 (.CI(n53691), .I0(n21901[5]), .I1(n542), .CO(n53692));
    SB_LUT4 add_5377_7_lut (.I0(GND_net), .I1(n21901[4]), .I2(n469), .I3(n53690), 
            .O(n21408[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_7 (.CI(n53690), .I0(n21901[4]), .I1(n469), .CO(n53691));
    SB_LUT4 add_5377_6_lut (.I0(GND_net), .I1(n21901[3]), .I2(n396), .I3(n53689), 
            .O(n21408[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_6 (.CI(n53689), .I0(n21901[3]), .I1(n396), .CO(n53690));
    SB_CARRY add_5194_10 (.CI(n53107), .I0(n19000[7]), .I1(n676), .CO(n53108));
    SB_LUT4 add_5377_5_lut (.I0(GND_net), .I1(n21901[2]), .I2(n323_adj_4456), 
            .I3(n53688), .O(n21408[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_5 (.CI(n53688), .I0(n21901[2]), .I1(n323_adj_4456), 
            .CO(n53689));
    SB_LUT4 add_5194_9_lut (.I0(GND_net), .I1(n19000[6]), .I2(n603_adj_4457), 
            .I3(n53106), .O(n17992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5377_4_lut (.I0(GND_net), .I1(n21901[1]), .I2(n250_adj_4458), 
            .I3(n53687), .O(n21408[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_4 (.CI(n53687), .I0(n21901[1]), .I1(n250_adj_4458), 
            .CO(n53688));
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5377_3_lut (.I0(GND_net), .I1(n21901[0]), .I2(n177_adj_4459), 
            .I3(n53686), .O(n21408[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_9 (.CI(n53106), .I0(n19000[6]), .I1(n603_adj_4457), 
            .CO(n53107));
    SB_LUT4 add_5194_8_lut (.I0(GND_net), .I1(n19000[5]), .I2(n530_adj_4460), 
            .I3(n53105), .O(n17992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_8 (.CI(n53105), .I0(n19000[5]), .I1(n530_adj_4460), 
            .CO(n53106));
    SB_LUT4 add_5194_7_lut (.I0(GND_net), .I1(n19000[4]), .I2(n457_adj_4461), 
            .I3(n53104), .O(n17992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n52741), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n52742));
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n52740), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_8 (.CI(n52740), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n52741));
    SB_LUT4 n9977_bdd_4_lut_51879 (.I0(n9977), .I1(n67715), .I2(setpoint[1]), 
            .I3(n4749), .O(n71409));
    defparam n9977_bdd_4_lut_51879.LUT_INIT = 16'he4aa;
    SB_CARRY add_5377_3 (.CI(n53686), .I0(n21901[0]), .I1(n177_adj_4459), 
            .CO(n53687));
    SB_CARRY add_5194_7 (.CI(n53104), .I0(n19000[4]), .I1(n457_adj_4461), 
            .CO(n53105));
    SB_LUT4 add_5377_2_lut (.I0(GND_net), .I1(n35_adj_4462), .I2(n104_adj_4463), 
            .I3(GND_net), .O(n21408[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5377_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5377_2 (.CI(GND_net), .I0(n35_adj_4462), .I1(n104_adj_4463), 
            .CO(n53686));
    SB_LUT4 add_5194_6_lut (.I0(GND_net), .I1(n19000[3]), .I2(n384_adj_4464), 
            .I3(n53103), .O(n17992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5194_6 (.CI(n53103), .I0(n19000[3]), .I1(n384_adj_4464), 
            .CO(n53104));
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n335[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4466));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4467));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i38_2_lut (.I0(\Ki[0] ), .I1(n335[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5194_5_lut (.I0(GND_net), .I1(n19000[2]), .I2(n311_adj_4469), 
            .I3(n53102), .O(n17992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n52739), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5194_5 (.CI(n53102), .I0(n19000[2]), .I1(n311_adj_4469), 
            .CO(n53103));
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4470));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4471));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5194_4_lut (.I0(GND_net), .I1(n19000[1]), .I2(n238_adj_4472), 
            .I3(n53101), .O(n17992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4473));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5194_4 (.CI(n53101), .I0(n19000[1]), .I1(n238_adj_4472), 
            .CO(n53102));
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4474));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5194_3_lut (.I0(GND_net), .I1(n19000[0]), .I2(n165_adj_4475), 
            .I3(n53100), .O(n17992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_3 (.CI(n53100), .I0(n19000[0]), .I1(n165_adj_4475), 
            .CO(n53101));
    SB_LUT4 add_5194_2_lut (.I0(GND_net), .I1(n23_adj_4476), .I2(n92_adj_4477), 
            .I3(GND_net), .O(n17992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5194_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5194_2 (.CI(GND_net), .I0(n23_adj_4476), .I1(n92_adj_4477), 
            .CO(n53100));
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4478));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71409_bdd_4_lut (.I0(n71409), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4749), .O(n71412));
    defparam n71409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY sub_15_add_2_7 (.CI(n52739), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n52740));
    SB_LUT4 add_5479_10_lut (.I0(GND_net), .I1(n22995[7]), .I2(n700), 
            .I3(n53099), .O(n22816[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5479_9_lut (.I0(GND_net), .I1(n22995[6]), .I2(n627), .I3(n53098), 
            .O(n22816[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4479));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n52738), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4480));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5479_9 (.CI(n53098), .I0(n22995[6]), .I1(n627), .CO(n53099));
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4482));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5479_8_lut (.I0(GND_net), .I1(n22995[5]), .I2(n554), .I3(n53097), 
            .O(n22816[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_6 (.CI(n52738), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n52739));
    SB_LUT4 n9977_bdd_4_lut_51874 (.I0(n9977), .I1(n67714), .I2(setpoint[0]), 
            .I3(n4749), .O(n71403));
    defparam n9977_bdd_4_lut_51874.LUT_INIT = 16'he4aa;
    SB_CARRY sub_15_add_2_5 (.CI(n52737), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n52738));
    SB_LUT4 n71403_bdd_4_lut (.I0(n71403), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4749), .O(n71406));
    defparam n71403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 counter_2045_2046_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n53621), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n53620), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_14 (.CI(n53620), .I0(GND_net), .I1(counter[12]), 
            .CO(n53621));
    SB_LUT4 counter_2045_2046_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n53619), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_13 (.CI(n53619), .I0(GND_net), .I1(counter[11]), 
            .CO(n53620));
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n53618), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_12 (.CI(n53618), .I0(GND_net), .I1(counter[10]), 
            .CO(n53619));
    SB_CARRY add_5479_8 (.CI(n53097), .I0(n22995[5]), .I1(n554), .CO(n53098));
    SB_LUT4 add_5479_7_lut (.I0(GND_net), .I1(n22995[4]), .I2(n481), .I3(n53096), 
            .O(n22816[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n53617), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_11 (.CI(n53617), .I0(GND_net), .I1(counter[9]), 
            .CO(n53618));
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n53616), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_10 (.CI(n53616), .I0(GND_net), .I1(counter[8]), 
            .CO(n53617));
    SB_LUT4 counter_2045_2046_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n53615), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_9 (.CI(n53615), .I0(GND_net), .I1(counter[7]), 
            .CO(n53616));
    SB_CARRY sub_15_add_2_4 (.CI(n52736), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n52737));
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n53614), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_8 (.CI(n53614), .I0(GND_net), .I1(counter[6]), 
            .CO(n53615));
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n53613), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(n23323[2]), .I1(n6_adj_4483), .I2(\Ki[4] ), 
            .I3(n335[18]), .O(n23266[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_CARRY counter_2045_2046_add_4_7 (.CI(n53613), .I0(GND_net), .I1(counter[5]), 
            .CO(n53614));
    SB_LUT4 counter_2045_2046_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n53612), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_6 (.CI(n53612), .I0(GND_net), .I1(counter[4]), 
            .CO(n53613));
    SB_LUT4 counter_2045_2046_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n53611), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_5 (.CI(n53611), .I0(GND_net), .I1(counter[3]), 
            .CO(n53612));
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4484));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n53610), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5479_7 (.CI(n53096), .I0(n22995[4]), .I1(n481), .CO(n53097));
    SB_LUT4 add_5479_6_lut (.I0(GND_net), .I1(n22995[3]), .I2(n408), .I3(n53095), 
            .O(n22816[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_3 (.CI(n52735), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n52736));
    SB_CARRY counter_2045_2046_add_4_4 (.CI(n53610), .I0(GND_net), .I1(counter[2]), 
            .CO(n53611));
    SB_CARRY add_5479_6 (.CI(n53095), .I0(n22995[3]), .I1(n408), .CO(n53096));
    SB_LUT4 counter_2045_2046_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n53609), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5479_5_lut (.I0(GND_net), .I1(n22995[2]), .I2(n335_c), 
            .I3(n53094), .O(n22816[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i138_2_lut (.I0(\Ki[2] ), .I1(n335[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_3 (.CI(n53609), .I0(GND_net), .I1(counter[1]), 
            .CO(n53610));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n52744), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state_c[0]), 
            .CO(n52735));
    SB_LUT4 add_5521_7_lut (.I0(GND_net), .I1(n62834), .I2(n490), .I3(n54080), 
            .O(n23217[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n53609));
    SB_LUT4 add_5521_6_lut (.I0(GND_net), .I1(n23287[3]), .I2(n417_adj_4485), 
            .I3(n54079), .O(n23217[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_6 (.CI(n54079), .I0(n23287[3]), .I1(n417_adj_4485), 
            .CO(n54080));
    SB_LUT4 add_5521_5_lut (.I0(GND_net), .I1(n23287[2]), .I2(n344_adj_4486), 
            .I3(n54078), .O(n23217[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5479_5 (.CI(n53094), .I0(n22995[2]), .I1(n335_c), .CO(n53095));
    SB_CARRY add_5521_5 (.CI(n54078), .I0(n23287[2]), .I1(n344_adj_4486), 
            .CO(n54079));
    SB_LUT4 add_5521_4_lut (.I0(GND_net), .I1(n23287[1]), .I2(n271_adj_4487), 
            .I3(n54077), .O(n23217[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5479_4_lut (.I0(GND_net), .I1(n22995[1]), .I2(n262), .I3(n53093), 
            .O(n22816[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_4 (.CI(n54077), .I0(n23287[1]), .I1(n271_adj_4487), 
            .CO(n54078));
    SB_LUT4 add_5521_3_lut (.I0(GND_net), .I1(n23287[0]), .I2(n198_adj_4488), 
            .I3(n54076), .O(n23217[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_3 (.CI(n54076), .I0(n23287[0]), .I1(n198_adj_4488), 
            .CO(n54077));
    SB_LUT4 add_5521_2_lut (.I0(GND_net), .I1(n56_adj_4489), .I2(n125_adj_4490), 
            .I3(GND_net), .O(n23217[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5521_2 (.CI(GND_net), .I0(n56_adj_4489), .I1(n125_adj_4490), 
            .CO(n54076));
    SB_LUT4 add_5472_10_lut (.I0(GND_net), .I1(n22935[7]), .I2(n700_adj_4491), 
            .I3(n54075), .O(n22739[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5472_9_lut (.I0(GND_net), .I1(n22935[6]), .I2(n627_adj_4492), 
            .I3(n54074), .O(n22739[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_9 (.CI(n54074), .I0(n22935[6]), .I1(n627_adj_4492), 
            .CO(n54075));
    SB_LUT4 add_5472_8_lut (.I0(GND_net), .I1(n22935[5]), .I2(n554_adj_4493), 
            .I3(n54073), .O(n22739[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5479_4 (.CI(n53093), .I0(n22995[1]), .I1(n262), .CO(n53094));
    SB_LUT4 add_5479_3_lut (.I0(GND_net), .I1(n22995[0]), .I2(n189), .I3(n53092), 
            .O(n22816[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_8 (.CI(n54073), .I0(n22935[5]), .I1(n554_adj_4493), 
            .CO(n54074));
    SB_LUT4 add_5472_7_lut (.I0(GND_net), .I1(n22935[4]), .I2(n481_adj_4494), 
            .I3(n54072), .O(n22739[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_7 (.CI(n54072), .I0(n22935[4]), .I1(n481_adj_4494), 
            .CO(n54073));
    SB_LUT4 add_5472_6_lut (.I0(GND_net), .I1(n22935[3]), .I2(n408_adj_4495), 
            .I3(n54071), .O(n22739[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_6 (.CI(n54071), .I0(n22935[3]), .I1(n408_adj_4495), 
            .CO(n54072));
    SB_LUT4 add_5472_5_lut (.I0(GND_net), .I1(n22935[2]), .I2(n335_adj_4496), 
            .I3(n54070), .O(n22739[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_5 (.CI(n54070), .I0(n22935[2]), .I1(n335_adj_4496), 
            .CO(n54071));
    SB_LUT4 add_5472_4_lut (.I0(GND_net), .I1(n22935[1]), .I2(n262_adj_4497), 
            .I3(n54069), .O(n22739[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_4 (.CI(n54069), .I0(n22935[1]), .I1(n262_adj_4497), 
            .CO(n54070));
    SB_LUT4 add_5472_3_lut (.I0(GND_net), .I1(n22935[0]), .I2(n189_adj_4498), 
            .I3(n54068), .O(n22739[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_3 (.CI(n54068), .I0(n22935[0]), .I1(n189_adj_4498), 
            .CO(n54069));
    SB_LUT4 add_5472_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n22739[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5472_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5472_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n54068));
    SB_LUT4 add_5489_9_lut (.I0(GND_net), .I1(n23076[6]), .I2(n630), .I3(n54067), 
            .O(n22935[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4499));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5489_8_lut (.I0(GND_net), .I1(n23076[5]), .I2(n557_adj_4500), 
            .I3(n54066), .O(n22935[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_8 (.CI(n54066), .I0(n23076[5]), .I1(n557_adj_4500), 
            .CO(n54067));
    SB_CARRY add_5479_3 (.CI(n53092), .I0(n22995[0]), .I1(n189), .CO(n53093));
    SB_LUT4 add_5489_7_lut (.I0(GND_net), .I1(n23076[4]), .I2(n484), .I3(n54065), 
            .O(n22935[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_7 (.CI(n54065), .I0(n23076[4]), .I1(n484), .CO(n54066));
    SB_LUT4 add_5489_6_lut (.I0(GND_net), .I1(n23076[3]), .I2(n411), .I3(n54064), 
            .O(n22935[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_6 (.CI(n54064), .I0(n23076[3]), .I1(n411), .CO(n54065));
    SB_LUT4 add_5489_5_lut (.I0(GND_net), .I1(n23076[2]), .I2(n338), .I3(n54063), 
            .O(n22935[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_5 (.CI(n54063), .I0(n23076[2]), .I1(n338), .CO(n54064));
    SB_LUT4 add_5489_4_lut (.I0(GND_net), .I1(n23076[1]), .I2(n265), .I3(n54062), 
            .O(n22935[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_4 (.CI(n54062), .I0(n23076[1]), .I1(n265), .CO(n54063));
    SB_LUT4 add_5489_3_lut (.I0(GND_net), .I1(n23076[0]), .I2(n192_adj_4501), 
            .I3(n54061), .O(n22935[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_3 (.CI(n54061), .I0(n23076[0]), .I1(n192_adj_4501), 
            .CO(n54062));
    SB_LUT4 add_5489_2_lut (.I0(GND_net), .I1(n50_adj_4502), .I2(n119_adj_4503), 
            .I3(GND_net), .O(n22935[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5489_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5489_2 (.CI(GND_net), .I0(n50_adj_4502), .I1(n119_adj_4503), 
            .CO(n54061));
    SB_LUT4 add_5479_2_lut (.I0(GND_net), .I1(n47_adj_4504), .I2(n116_adj_4505), 
            .I3(GND_net), .O(n22816[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5479_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5479_2 (.CI(GND_net), .I0(n47_adj_4504), .I1(n116_adj_4505), 
            .CO(n53092));
    SB_LUT4 i1_4_lut_adj_944 (.I0(n23381[0]), .I1(n52428), .I2(\Ki[2] ), 
            .I3(n335[20]), .O(n23360[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_944.LUT_INIT = 16'h9666;
    SB_LUT4 add_5243_17_lut (.I0(GND_net), .I1(n19879[14]), .I2(GND_net), 
            .I3(n53091), .O(n19000[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i89_2_lut (.I0(\Ki[1] ), .I1(n335[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i42_2_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4506));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5243_16_lut (.I0(GND_net), .I1(n19879[13]), .I2(n1117_adj_4507), 
            .I3(n53090), .O(n19000[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_16 (.CI(n53090), .I0(n19879[13]), .I1(n1117_adj_4507), 
            .CO(n53091));
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4507));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5243_15_lut (.I0(GND_net), .I1(n19879[12]), .I2(n1044_adj_4499), 
            .I3(n53089), .O(n19000[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5243_15 (.CI(n53089), .I0(n19879[12]), .I1(n1044_adj_4499), 
            .CO(n53090));
    SB_LUT4 add_5243_14_lut (.I0(GND_net), .I1(n19879[11]), .I2(n971_adj_4484), 
            .I3(n53088), .O(n19000[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_14 (.CI(n53088), .I0(n19879[11]), .I1(n971_adj_4484), 
            .CO(n53089));
    SB_LUT4 add_5243_13_lut (.I0(GND_net), .I1(n19879[10]), .I2(n898_adj_4474), 
            .I3(n53087), .O(n19000[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_13 (.CI(n53087), .I0(n19879[10]), .I1(n898_adj_4474), 
            .CO(n53088));
    SB_LUT4 add_5504_8_lut (.I0(GND_net), .I1(n23185[5]), .I2(n560), .I3(n53973), 
            .O(n23076[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5504_7_lut (.I0(GND_net), .I1(n23185[4]), .I2(n487), .I3(n53972), 
            .O(n23076[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_7 (.CI(n53972), .I0(n23185[4]), .I1(n487), .CO(n53973));
    SB_LUT4 add_5504_6_lut (.I0(GND_net), .I1(n23185[3]), .I2(n414), .I3(n53971), 
            .O(n23076[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_6 (.CI(n53971), .I0(n23185[3]), .I1(n414), .CO(n53972));
    SB_LUT4 add_5504_5_lut (.I0(GND_net), .I1(n23185[2]), .I2(n341), .I3(n53970), 
            .O(n23076[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_5 (.CI(n53970), .I0(n23185[2]), .I1(n341), .CO(n53971));
    SB_LUT4 add_5504_4_lut (.I0(GND_net), .I1(n23185[1]), .I2(n268), .I3(n53969), 
            .O(n23076[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_4 (.CI(n53969), .I0(n23185[1]), .I1(n268), .CO(n53970));
    SB_LUT4 add_5504_3_lut (.I0(GND_net), .I1(n23185[0]), .I2(n195), .I3(n53968), 
            .O(n23076[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_3 (.CI(n53968), .I0(n23185[0]), .I1(n195), .CO(n53969));
    SB_LUT4 add_5504_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n23076[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5504_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5504_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n53968));
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5409_13_lut (.I0(GND_net), .I1(n22294[10]), .I2(n910), 
            .I3(n53506), .O(n21901[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5409_12_lut (.I0(GND_net), .I1(n22294[9]), .I2(n837), 
            .I3(n53505), .O(n21901[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_12 (.CI(n53505), .I0(n22294[9]), .I1(n837), .CO(n53506));
    SB_LUT4 add_5409_11_lut (.I0(GND_net), .I1(n22294[8]), .I2(n764), 
            .I3(n53504), .O(n21901[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_11 (.CI(n53504), .I0(n22294[8]), .I1(n764), .CO(n53505));
    SB_LUT4 add_5409_10_lut (.I0(GND_net), .I1(n22294[7]), .I2(n691), 
            .I3(n53503), .O(n21901[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_10 (.CI(n53503), .I0(n22294[7]), .I1(n691), .CO(n53504));
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n335[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n310[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5409_9_lut (.I0(GND_net), .I1(n22294[6]), .I2(n618), .I3(n53502), 
            .O(n21901[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i22_3_lut (.I0(n310[21]), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n335[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5409_9 (.CI(n53502), .I0(n22294[6]), .I1(n618), .CO(n53503));
    SB_LUT4 add_5409_8_lut (.I0(GND_net), .I1(n22294[5]), .I2(n545), .I3(n53501), 
            .O(n21901[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_8 (.CI(n53501), .I0(n22294[5]), .I1(n545), .CO(n53502));
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4505));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4504));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n335[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5409_7_lut (.I0(GND_net), .I1(n22294[4]), .I2(n472), .I3(n53500), 
            .O(n21901[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_7 (.CI(n53500), .I0(n22294[4]), .I1(n472), .CO(n53501));
    SB_LUT4 add_5409_6_lut (.I0(GND_net), .I1(n22294[3]), .I2(n399), .I3(n53499), 
            .O(n21901[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_6 (.CI(n53499), .I0(n22294[3]), .I1(n399), .CO(n53500));
    SB_LUT4 add_5409_5_lut (.I0(GND_net), .I1(n22294[2]), .I2(n326), .I3(n53498), 
            .O(n21901[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_5 (.CI(n53498), .I0(n22294[2]), .I1(n326), .CO(n53499));
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n335[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5409_4_lut (.I0(GND_net), .I1(n22294[1]), .I2(n253), .I3(n53497), 
            .O(n21901[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_4 (.CI(n53497), .I0(n22294[1]), .I1(n253), .CO(n53498));
    SB_LUT4 add_5409_3_lut (.I0(GND_net), .I1(n22294[0]), .I2(n180), .I3(n53496), 
            .O(n21901[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_3 (.CI(n53496), .I0(n22294[0]), .I1(n180), .CO(n53497));
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n335[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5409_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n21901[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5409_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5409_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n53496));
    SB_LUT4 add_5243_12_lut (.I0(GND_net), .I1(n19879[9]), .I2(n825_adj_4449), 
            .I3(n53086), .O(n19000[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_12 (.CI(n53086), .I0(n19879[9]), .I1(n825_adj_4449), 
            .CO(n53087));
    SB_LUT4 add_5243_11_lut (.I0(GND_net), .I1(n19879[8]), .I2(n752), 
            .I3(n53085), .O(n19000[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_11 (.CI(n53085), .I0(n19879[8]), .I1(n752), .CO(n53086));
    SB_LUT4 add_5243_10_lut (.I0(GND_net), .I1(n19879[7]), .I2(n679), 
            .I3(n53084), .O(n19000[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i19_3_lut (.I0(n233[18]), .I1(n285[18]), .I2(n284), 
            .I3(GND_net), .O(n310[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5243_10 (.CI(n53084), .I0(n19879[7]), .I1(n679), .CO(n53085));
    SB_LUT4 add_5243_9_lut (.I0(GND_net), .I1(n19879[6]), .I2(n606), .I3(n53083), 
            .O(n19000[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_9 (.CI(n53083), .I0(n19879[6]), .I1(n606), .CO(n53084));
    SB_LUT4 add_5243_8_lut (.I0(GND_net), .I1(n19879[5]), .I2(n533), .I3(n53082), 
            .O(n19000[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_8 (.CI(n53082), .I0(n19879[5]), .I1(n533), .CO(n53083));
    SB_LUT4 mux_22_i19_3_lut (.I0(n310[18]), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n335[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5243_7_lut (.I0(GND_net), .I1(n19879[4]), .I2(n460), .I3(n53081), 
            .O(n19000[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_7 (.CI(n53081), .I0(n19879[4]), .I1(n460), .CO(n53082));
    SB_LUT4 add_5243_6_lut (.I0(GND_net), .I1(n19879[3]), .I2(n387), .I3(n53080), 
            .O(n19000[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_6 (.CI(n53080), .I0(n19879[3]), .I1(n387), .CO(n53081));
    SB_LUT4 add_5243_5_lut (.I0(GND_net), .I1(n19879[2]), .I2(n314), .I3(n53079), 
            .O(n19000[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_5 (.CI(n53079), .I0(n19879[2]), .I1(n314), .CO(n53080));
    SB_LUT4 add_5243_4_lut (.I0(GND_net), .I1(n19879[1]), .I2(n241_adj_4513), 
            .I3(n53078), .O(n19000[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4514));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_945 (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(n335[23]), 
            .I3(n335[22]), .O(n64007));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h9c50;
    SB_CARRY add_5243_4 (.CI(n53078), .I0(n19879[1]), .I1(n241_adj_4513), 
            .CO(n53079));
    SB_LUT4 add_5243_3_lut (.I0(GND_net), .I1(n19879[0]), .I2(n168_adj_4515), 
            .I3(n53077), .O(n19000[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_3 (.CI(n53077), .I0(n19879[0]), .I1(n168_adj_4515), 
            .CO(n53078));
    SB_LUT4 add_5243_2_lut (.I0(GND_net), .I1(n26_adj_4516), .I2(n95_adj_4517), 
            .I3(GND_net), .O(n19000[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5243_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5243_2 (.CI(GND_net), .I0(n26_adj_4516), .I1(n95_adj_4517), 
            .CO(n53077));
    SB_LUT4 add_5289_16_lut (.I0(GND_net), .I1(n20618[13]), .I2(n1120_adj_4518), 
            .I3(n53076), .O(n19879[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5289_15_lut (.I0(GND_net), .I1(n20618[12]), .I2(n1047_adj_4519), 
            .I3(n53075), .O(n19879[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_15 (.CI(n53075), .I0(n20618[12]), .I1(n1047_adj_4519), 
            .CO(n53076));
    SB_LUT4 add_5289_14_lut (.I0(GND_net), .I1(n20618[11]), .I2(n974_adj_4520), 
            .I3(n53074), .O(n19879[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_14 (.CI(n53074), .I0(n20618[11]), .I1(n974_adj_4520), 
            .CO(n53075));
    SB_LUT4 add_5289_13_lut (.I0(GND_net), .I1(n20618[10]), .I2(n901_adj_4521), 
            .I3(n53073), .O(n19879[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_13 (.CI(n53073), .I0(n20618[10]), .I1(n901_adj_4521), 
            .CO(n53074));
    SB_LUT4 add_5289_12_lut (.I0(GND_net), .I1(n20618[9]), .I2(n828_adj_4522), 
            .I3(n53072), .O(n19879[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_12 (.CI(n53072), .I0(n20618[9]), .I1(n828_adj_4522), 
            .CO(n53073));
    SB_LUT4 add_5289_11_lut (.I0(GND_net), .I1(n20618[8]), .I2(n755_adj_4523), 
            .I3(n53071), .O(n19879[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_11 (.CI(n53071), .I0(n20618[8]), .I1(n755_adj_4523), 
            .CO(n53072));
    SB_LUT4 add_5289_10_lut (.I0(GND_net), .I1(n20618[7]), .I2(n682_adj_4524), 
            .I3(n53070), .O(n19879[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_10 (.CI(n53070), .I0(n20618[7]), .I1(n682_adj_4524), 
            .CO(n53071));
    SB_LUT4 add_5289_9_lut (.I0(GND_net), .I1(n20618[6]), .I2(n609_adj_4525), 
            .I3(n53069), .O(n19879[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_9 (.CI(n53069), .I0(n20618[6]), .I1(n609_adj_4525), 
            .CO(n53070));
    SB_LUT4 add_5289_8_lut (.I0(GND_net), .I1(n20618[5]), .I2(n536_adj_4526), 
            .I3(n53068), .O(n19879[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_8 (.CI(n53068), .I0(n20618[5]), .I1(n536_adj_4526), 
            .CO(n53069));
    SB_LUT4 add_5289_7_lut (.I0(GND_net), .I1(n20618[4]), .I2(n463_adj_4527), 
            .I3(n53067), .O(n19879[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_7 (.CI(n53067), .I0(n20618[4]), .I1(n463_adj_4527), 
            .CO(n53068));
    SB_LUT4 add_5289_6_lut (.I0(GND_net), .I1(n20618[3]), .I2(n390_adj_4528), 
            .I3(n53066), .O(n19879[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_6 (.CI(n53066), .I0(n20618[3]), .I1(n390_adj_4528), 
            .CO(n53067));
    SB_LUT4 add_5289_5_lut (.I0(GND_net), .I1(n20618[2]), .I2(n317_adj_4529), 
            .I3(n53065), .O(n19879[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_5 (.CI(n53065), .I0(n20618[2]), .I1(n317_adj_4529), 
            .CO(n53066));
    SB_LUT4 add_5289_4_lut (.I0(GND_net), .I1(n20618[1]), .I2(n244_adj_4530), 
            .I3(n53064), .O(n19879[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_4 (.CI(n53064), .I0(n20618[1]), .I1(n244_adj_4530), 
            .CO(n53065));
    SB_LUT4 add_5289_3_lut (.I0(GND_net), .I1(n20618[0]), .I2(n171_adj_4531), 
            .I3(n53063), .O(n19879[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(n335[18]), 
            .I3(n335[19]), .O(n64011));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h6ca0;
    SB_CARRY add_5289_3 (.CI(n53063), .I0(n20618[0]), .I1(n171_adj_4531), 
            .CO(n53064));
    SB_LUT4 add_5289_2_lut (.I0(GND_net), .I1(n29_adj_4532), .I2(n98_adj_4533), 
            .I3(GND_net), .O(n19879[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5289_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5289_2 (.CI(GND_net), .I0(n29_adj_4532), .I1(n98_adj_4533), 
            .CO(n53063));
    SB_LUT4 add_5329_15_lut (.I0(GND_net), .I1(n21243[12]), .I2(n1050_adj_4534), 
            .I3(n53062), .O(n20618[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5329_14_lut (.I0(GND_net), .I1(n21243[11]), .I2(n977_adj_4535), 
            .I3(n53061), .O(n20618[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_14 (.CI(n53061), .I0(n21243[11]), .I1(n977_adj_4535), 
            .CO(n53062));
    SB_LUT4 add_5329_13_lut (.I0(GND_net), .I1(n21243[10]), .I2(n904_adj_4536), 
            .I3(n53060), .O(n20618[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_13 (.CI(n53060), .I0(n21243[10]), .I1(n904_adj_4536), 
            .CO(n53061));
    SB_LUT4 add_5329_12_lut (.I0(GND_net), .I1(n21243[9]), .I2(n831_adj_4537), 
            .I3(n53059), .O(n20618[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_12 (.CI(n53059), .I0(n21243[9]), .I1(n831_adj_4537), 
            .CO(n53060));
    SB_LUT4 add_5329_11_lut (.I0(GND_net), .I1(n21243[8]), .I2(n758_adj_4538), 
            .I3(n53058), .O(n20618[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_11 (.CI(n53058), .I0(n21243[8]), .I1(n758_adj_4538), 
            .CO(n53059));
    SB_LUT4 add_5329_10_lut (.I0(GND_net), .I1(n21243[7]), .I2(n685_adj_4539), 
            .I3(n53057), .O(n20618[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_10 (.CI(n53057), .I0(n21243[7]), .I1(n685_adj_4539), 
            .CO(n53058));
    SB_LUT4 i1_4_lut_adj_947 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(n335[20]), 
            .I3(n335[21]), .O(n64009));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_5329_9_lut (.I0(GND_net), .I1(n21243[6]), .I2(n612_adj_4540), 
            .I3(n53056), .O(n20618[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_9 (.CI(n53056), .I0(n21243[6]), .I1(n612_adj_4540), 
            .CO(n53057));
    SB_LUT4 add_5329_8_lut (.I0(GND_net), .I1(n21243[5]), .I2(n539_adj_4541), 
            .I3(n53055), .O(n20618[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_8 (.CI(n53055), .I0(n21243[5]), .I1(n539_adj_4541), 
            .CO(n53056));
    SB_LUT4 add_5329_7_lut (.I0(GND_net), .I1(n21243[4]), .I2(n466_adj_4542), 
            .I3(n53054), .O(n20618[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_7 (.CI(n53054), .I0(n21243[4]), .I1(n466_adj_4542), 
            .CO(n53055));
    SB_LUT4 add_5329_6_lut (.I0(GND_net), .I1(n21243[3]), .I2(n393_adj_4543), 
            .I3(n53053), .O(n20618[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_6 (.CI(n53053), .I0(n21243[3]), .I1(n393_adj_4543), 
            .CO(n53054));
    SB_LUT4 add_5329_5_lut (.I0(GND_net), .I1(n21243[2]), .I2(n320_adj_4544), 
            .I3(n53052), .O(n20618[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_5 (.CI(n53052), .I0(n21243[2]), .I1(n320_adj_4544), 
            .CO(n53053));
    SB_LUT4 add_5329_4_lut (.I0(GND_net), .I1(n21243[1]), .I2(n247_adj_4545), 
            .I3(n53051), .O(n20618[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n64009), .I1(n52398), .I2(n64011), .I3(n64007), 
            .O(n64017));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i34409_4_lut (.I0(n23381[0]), .I1(\Ki[2] ), .I2(n52428), .I3(n335[20]), 
            .O(n4));   // verilog/motorControl.v(61[29:40])
    defparam i34409_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5329_4 (.CI(n53051), .I0(n21243[1]), .I1(n247_adj_4545), 
            .CO(n53052));
    SB_LUT4 add_5329_3_lut (.I0(GND_net), .I1(n21243[0]), .I2(n174_adj_4547), 
            .I3(n53050), .O(n20618[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5329_3 (.CI(n53050), .I0(n21243[0]), .I1(n174_adj_4547), 
            .CO(n53051));
    SB_LUT4 add_5329_2_lut (.I0(GND_net), .I1(n32_adj_4548), .I2(n101_adj_4549), 
            .I3(GND_net), .O(n20618[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5329_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34547_4_lut (.I0(n23323[2]), .I1(\Ki[4] ), .I2(n6_adj_4483), 
            .I3(n335[18]), .O(n8));   // verilog/motorControl.v(61[29:40])
    defparam i34547_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n335[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5329_2 (.CI(GND_net), .I0(n32_adj_4548), .I1(n101_adj_4549), 
            .CO(n53050));
    SB_LUT4 add_5495_9_lut (.I0(GND_net), .I1(n23121[6]), .I2(n630_adj_4550), 
            .I3(n53049), .O(n22995[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4503));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4502));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9977_bdd_4_lut_52082 (.I0(n9977), .I1(n67737), .I2(setpoint[22]), 
            .I3(n4749), .O(n71547));
    defparam n9977_bdd_4_lut_52082.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n6_adj_4552), .I1(n8), .I2(n4), .I3(n64017), 
            .O(n62888));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 add_5495_8_lut (.I0(GND_net), .I1(n23121[5]), .I2(n557_adj_4553), 
            .I3(n53048), .O(n22995[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_8 (.CI(n53048), .I0(n23121[5]), .I1(n557_adj_4553), 
            .CO(n53049));
    SB_LUT4 add_5495_7_lut (.I0(GND_net), .I1(n23121[4]), .I2(n484_adj_4554), 
            .I3(n53047), .O(n22995[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_7 (.CI(n53047), .I0(n23121[4]), .I1(n484_adj_4554), 
            .CO(n53048));
    SB_LUT4 n71547_bdd_4_lut (.I0(n71547), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4749), .O(n71550));
    defparam n71547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5495_6_lut (.I0(GND_net), .I1(n23121[3]), .I2(n411_adj_4556), 
            .I3(n53046), .O(n22995[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_6 (.CI(n53046), .I0(n23121[3]), .I1(n411_adj_4556), 
            .CO(n53047));
    SB_LUT4 add_5495_5_lut (.I0(GND_net), .I1(n23121[2]), .I2(n338_adj_4557), 
            .I3(n53045), .O(n22995[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_5 (.CI(n53045), .I0(n23121[2]), .I1(n338_adj_4557), 
            .CO(n53046));
    SB_LUT4 add_5495_4_lut (.I0(GND_net), .I1(n23121[1]), .I2(n265_adj_4558), 
            .I3(n53044), .O(n22995[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5517_7_lut (.I0(GND_net), .I1(n62888), .I2(n490_adj_4514), 
            .I3(n53918), .O(n23185[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_4 (.CI(n53044), .I0(n23121[1]), .I1(n265_adj_4558), 
            .CO(n53045));
    SB_LUT4 add_5517_6_lut (.I0(GND_net), .I1(n23266[3]), .I2(n417), .I3(n53917), 
            .O(n23185[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5495_3_lut (.I0(GND_net), .I1(n23121[0]), .I2(n192), .I3(n53043), 
            .O(n22995[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_6 (.CI(n53917), .I0(n23266[3]), .I1(n417), .CO(n53918));
    SB_CARRY add_5495_3 (.CI(n53043), .I0(n23121[0]), .I1(n192), .CO(n53044));
    SB_LUT4 add_5495_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n22995[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5495_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5517_5_lut (.I0(GND_net), .I1(n23266[2]), .I2(n344), .I3(n53916), 
            .O(n23185[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5495_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n53043));
    SB_LUT4 add_5366_14_lut (.I0(GND_net), .I1(n21761[11]), .I2(n980_adj_4482), 
            .I3(n53042), .O(n21243[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5366_13_lut (.I0(GND_net), .I1(n21761[10]), .I2(n907_adj_4481), 
            .I3(n53041), .O(n21243[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_5 (.CI(n53916), .I0(n23266[2]), .I1(n344), .CO(n53917));
    SB_CARRY add_5366_13 (.CI(n53041), .I0(n21761[10]), .I1(n907_adj_4481), 
            .CO(n53042));
    SB_LUT4 add_5366_12_lut (.I0(GND_net), .I1(n21761[9]), .I2(n834_adj_4480), 
            .I3(n53040), .O(n21243[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_12 (.CI(n53040), .I0(n21761[9]), .I1(n834_adj_4480), 
            .CO(n53041));
    SB_LUT4 add_5366_11_lut (.I0(GND_net), .I1(n21761[8]), .I2(n761_adj_4479), 
            .I3(n53039), .O(n21243[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_11 (.CI(n53039), .I0(n21761[8]), .I1(n761_adj_4479), 
            .CO(n53040));
    SB_LUT4 add_5517_4_lut (.I0(GND_net), .I1(n23266[1]), .I2(n271), .I3(n53915), 
            .O(n23185[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5366_10_lut (.I0(GND_net), .I1(n21761[7]), .I2(n688_adj_4478), 
            .I3(n53038), .O(n21243[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_4 (.CI(n53915), .I0(n23266[1]), .I1(n271), .CO(n53916));
    SB_CARRY add_5366_10 (.CI(n53038), .I0(n21761[7]), .I1(n688_adj_4478), 
            .CO(n53039));
    SB_LUT4 add_5517_3_lut (.I0(GND_net), .I1(n23266[0]), .I2(n198), .I3(n53914), 
            .O(n23185[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5366_9_lut (.I0(GND_net), .I1(n21761[6]), .I2(n615_adj_4473), 
            .I3(n53037), .O(n21243[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_9 (.CI(n53037), .I0(n21761[6]), .I1(n615_adj_4473), 
            .CO(n53038));
    SB_LUT4 add_5366_8_lut (.I0(GND_net), .I1(n21761[5]), .I2(n542_adj_4471), 
            .I3(n53036), .O(n21243[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5517_3 (.CI(n53914), .I0(n23266[0]), .I1(n198), .CO(n53915));
    SB_CARRY add_5366_8 (.CI(n53036), .I0(n21761[5]), .I1(n542_adj_4471), 
            .CO(n53037));
    SB_LUT4 add_5366_7_lut (.I0(GND_net), .I1(n21761[4]), .I2(n469_adj_4470), 
            .I3(n53035), .O(n21243[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_7 (.CI(n53035), .I0(n21761[4]), .I1(n469_adj_4470), 
            .CO(n53036));
    SB_LUT4 add_5517_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n23185[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5517_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5366_6_lut (.I0(GND_net), .I1(n21761[3]), .I2(n396_adj_4467), 
            .I3(n53034), .O(n21243[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_6 (.CI(n53034), .I0(n21761[3]), .I1(n396_adj_4467), 
            .CO(n53035));
    SB_LUT4 add_5366_5_lut (.I0(GND_net), .I1(n21761[2]), .I2(n323_adj_4466), 
            .I3(n53033), .O(n21243[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_5 (.CI(n53033), .I0(n21761[2]), .I1(n323_adj_4466), 
            .CO(n53034));
    SB_LUT4 add_5366_4_lut (.I0(GND_net), .I1(n21761[1]), .I2(n250), .I3(n53032), 
            .O(n21243[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_4 (.CI(n53032), .I0(n21761[1]), .I1(n250), .CO(n53033));
    SB_CARRY add_5517_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n53914));
    SB_LUT4 add_5366_3_lut (.I0(GND_net), .I1(n21761[0]), .I2(n177), .I3(n53031), 
            .O(n21243[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_3 (.CI(n53031), .I0(n21761[0]), .I1(n177), .CO(n53032));
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n11135[21]), .I2(GND_net), 
            .I3(n53913), .O(n10676[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n11135[20]), .I2(GND_net), 
            .I3(n53912), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5366_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n21243[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5366_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5366_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n53031));
    SB_LUT4 add_5399_13_lut (.I0(GND_net), .I1(n22177[10]), .I2(n910_adj_4559), 
            .I3(n53030), .O(n21761[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n53912), .I0(n11135[20]), .I1(GND_net), 
            .CO(n53913));
    SB_LUT4 add_5399_12_lut (.I0(GND_net), .I1(n22177[9]), .I2(n837_adj_4560), 
            .I3(n53029), .O(n21761[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_12 (.CI(n53029), .I0(n22177[9]), .I1(n837_adj_4560), 
            .CO(n53030));
    SB_LUT4 add_5399_11_lut (.I0(GND_net), .I1(n22177[8]), .I2(n764_adj_4561), 
            .I3(n53028), .O(n21761[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n11135[19]), .I2(GND_net), 
            .I3(n53911), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_11 (.CI(n53028), .I0(n22177[8]), .I1(n764_adj_4561), 
            .CO(n53029));
    SB_LUT4 add_5399_10_lut (.I0(GND_net), .I1(n22177[7]), .I2(n691_adj_4562), 
            .I3(n53027), .O(n21761[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_22 (.CI(n53911), .I0(n11135[19]), .I1(GND_net), 
            .CO(n53912));
    SB_CARRY add_5399_10 (.CI(n53027), .I0(n22177[7]), .I1(n691_adj_4562), 
            .CO(n53028));
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n11135[18]), .I2(GND_net), 
            .I3(n53910), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n53910), .I0(n11135[18]), .I1(GND_net), 
            .CO(n53911));
    SB_LUT4 add_5399_9_lut (.I0(GND_net), .I1(n22177[6]), .I2(n618_adj_4564), 
            .I3(n53026), .O(n21761[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5436_12_lut (.I0(GND_net), .I1(n22597[9]), .I2(n840), 
            .I3(n53290), .O(n22294[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_9 (.CI(n53026), .I0(n22177[6]), .I1(n618_adj_4564), 
            .CO(n53027));
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n11135[17]), .I2(GND_net), 
            .I3(n53909), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5436_11_lut (.I0(GND_net), .I1(n22597[8]), .I2(n767), 
            .I3(n53289), .O(n22294[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5399_8_lut (.I0(GND_net), .I1(n22177[5]), .I2(n545_adj_4565), 
            .I3(n53025), .O(n21761[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_8 (.CI(n53025), .I0(n22177[5]), .I1(n545_adj_4565), 
            .CO(n53026));
    SB_CARRY add_5436_11 (.CI(n53289), .I0(n22597[8]), .I1(n767), .CO(n53290));
    SB_LUT4 add_5399_7_lut (.I0(GND_net), .I1(n22177[4]), .I2(n472_adj_4566), 
            .I3(n53024), .O(n21761[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_7 (.CI(n53024), .I0(n22177[4]), .I1(n472_adj_4566), 
            .CO(n53025));
    SB_CARRY mult_23_add_1221_20 (.CI(n53909), .I0(n11135[17]), .I1(GND_net), 
            .CO(n53910));
    SB_LUT4 add_5436_10_lut (.I0(GND_net), .I1(n22597[7]), .I2(n694), 
            .I3(n53288), .O(n22294[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5399_6_lut (.I0(GND_net), .I1(n22177[3]), .I2(n399_adj_4567), 
            .I3(n53023), .O(n21761[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_6 (.CI(n53023), .I0(n22177[3]), .I1(n399_adj_4567), 
            .CO(n53024));
    SB_CARRY add_5436_10 (.CI(n53288), .I0(n22597[7]), .I1(n694), .CO(n53289));
    SB_LUT4 add_5399_5_lut (.I0(GND_net), .I1(n22177[2]), .I2(n326_adj_4568), 
            .I3(n53022), .O(n21761[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_5 (.CI(n53022), .I0(n22177[2]), .I1(n326_adj_4568), 
            .CO(n53023));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n11135[16]), .I2(GND_net), 
            .I3(n53908), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n53908), .I0(n11135[16]), .I1(GND_net), 
            .CO(n53909));
    SB_LUT4 add_5436_9_lut (.I0(GND_net), .I1(n22597[6]), .I2(n621), .I3(n53287), 
            .O(n22294[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5399_4_lut (.I0(GND_net), .I1(n22177[1]), .I2(n253_adj_4569), 
            .I3(n53021), .O(n21761[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_4 (.CI(n53021), .I0(n22177[1]), .I1(n253_adj_4569), 
            .CO(n53022));
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n11135[15]), .I2(GND_net), 
            .I3(n53907), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_18 (.CI(n53907), .I0(n11135[15]), .I1(GND_net), 
            .CO(n53908));
    SB_CARRY add_5436_9 (.CI(n53287), .I0(n22597[6]), .I1(n621), .CO(n53288));
    SB_LUT4 add_5399_3_lut (.I0(GND_net), .I1(n22177[0]), .I2(n180_adj_4571), 
            .I3(n53020), .O(n21761[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_3 (.CI(n53020), .I0(n22177[0]), .I1(n180_adj_4571), 
            .CO(n53021));
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n11135[14]), .I2(GND_net), 
            .I3(n53906), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5436_8_lut (.I0(GND_net), .I1(n22597[5]), .I2(n548), .I3(n53286), 
            .O(n22294[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5399_2_lut (.I0(GND_net), .I1(n38_adj_4572), .I2(n107_adj_4573), 
            .I3(GND_net), .O(n21761[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5399_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5399_2 (.CI(GND_net), .I0(n38_adj_4572), .I1(n107_adj_4573), 
            .CO(n53020));
    SB_CARRY add_5436_8 (.CI(n53286), .I0(n22597[5]), .I1(n548), .CO(n53287));
    SB_LUT4 add_5509_8_lut (.I0(GND_net), .I1(n23217[5]), .I2(n560_adj_4574), 
            .I3(n53019), .O(n23121[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4558));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5509_7_lut (.I0(GND_net), .I1(n23217[4]), .I2(n487_adj_4575), 
            .I3(n53018), .O(n23121[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5436_7_lut (.I0(GND_net), .I1(n22597[4]), .I2(n475), .I3(n53285), 
            .O(n22294[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5509_7 (.CI(n53018), .I0(n23217[4]), .I1(n487_adj_4575), 
            .CO(n53019));
    SB_CARRY mult_23_add_1221_17 (.CI(n53906), .I0(n11135[14]), .I1(GND_net), 
            .CO(n53907));
    SB_CARRY add_5436_7 (.CI(n53285), .I0(n22597[4]), .I1(n475), .CO(n53286));
    SB_LUT4 add_5509_6_lut (.I0(GND_net), .I1(n23217[3]), .I2(n414_adj_4576), 
            .I3(n53017), .O(n23121[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5509_6 (.CI(n53017), .I0(n23217[3]), .I1(n414_adj_4576), 
            .CO(n53018));
    SB_LUT4 add_5436_6_lut (.I0(GND_net), .I1(n22597[3]), .I2(n402), .I3(n53284), 
            .O(n22294[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5509_5_lut (.I0(GND_net), .I1(n23217[2]), .I2(n341_adj_4577), 
            .I3(n53016), .O(n23121[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5509_5 (.CI(n53016), .I0(n23217[2]), .I1(n341_adj_4577), 
            .CO(n53017));
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n11135[13]), .I2(n1096), 
            .I3(n53905), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n53905), .I0(n11135[13]), .I1(n1096), 
            .CO(n53906));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n11135[12]), .I2(n1023), 
            .I3(n53904), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5436_6 (.CI(n53284), .I0(n22597[3]), .I1(n402), .CO(n53285));
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4557));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9977_bdd_4_lut_51988 (.I0(n9977), .I1(n67735), .I2(setpoint[21]), 
            .I3(n4749), .O(n71541));
    defparam n9977_bdd_4_lut_51988.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5436_5_lut (.I0(GND_net), .I1(n22597[2]), .I2(n329), .I3(n53283), 
            .O(n22294[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5509_4_lut (.I0(GND_net), .I1(n23217[1]), .I2(n268_adj_4579), 
            .I3(n53015), .O(n23121[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4556));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5509_4 (.CI(n53015), .I0(n23217[1]), .I1(n268_adj_4579), 
            .CO(n53016));
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4554));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4553));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5509_3_lut (.I0(GND_net), .I1(n23217[0]), .I2(n195_adj_4580), 
            .I3(n53014), .O(n23121[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_2045_2046__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n71664), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY mult_23_add_1221_15 (.CI(n53904), .I0(n11135[12]), .I1(n1023), 
            .CO(n53905));
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n11135[11]), .I2(n950), 
            .I3(n53903), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5436_5 (.CI(n53283), .I0(n22597[2]), .I1(n329), .CO(n53284));
    SB_CARRY add_5509_3 (.CI(n53014), .I0(n23217[0]), .I1(n195_adj_4580), 
            .CO(n53015));
    SB_LUT4 add_5509_2_lut (.I0(GND_net), .I1(n53_adj_4581), .I2(n122_adj_4582), 
            .I3(GND_net), .O(n23121[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5509_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_14 (.CI(n53903), .I0(n11135[11]), .I1(n950), 
            .CO(n53904));
    SB_LUT4 add_5436_4_lut (.I0(GND_net), .I1(n22597[1]), .I2(n256), .I3(n53282), 
            .O(n22294[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5509_2 (.CI(GND_net), .I0(n53_adj_4581), .I1(n122_adj_4582), 
            .CO(n53014));
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n11135[10]), .I2(n877), 
            .I3(n53902), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5427_12_lut (.I0(GND_net), .I1(n22501[9]), .I2(n840_adj_4583), 
            .I3(n53013), .O(n22177[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5436_4 (.CI(n53282), .I0(n22597[1]), .I1(n256), .CO(n53283));
    SB_LUT4 add_5427_11_lut (.I0(GND_net), .I1(n22501[8]), .I2(n767_adj_4584), 
            .I3(n53012), .O(n22177[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_11 (.CI(n53012), .I0(n22501[8]), .I1(n767_adj_4584), 
            .CO(n53013));
    SB_LUT4 add_5427_10_lut (.I0(GND_net), .I1(n22501[7]), .I2(n694_adj_4585), 
            .I3(n53011), .O(n22177[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_13 (.CI(n53902), .I0(n11135[10]), .I1(n877), 
            .CO(n53903));
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n11135[9]), .I2(n804), 
            .I3(n53901), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5436_3_lut (.I0(GND_net), .I1(n22597[0]), .I2(n183), .I3(n53281), 
            .O(n22294[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5436_3 (.CI(n53281), .I0(n22597[0]), .I1(n183), .CO(n53282));
    SB_LUT4 add_5436_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n22294[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_10 (.CI(n53011), .I0(n22501[7]), .I1(n694_adj_4585), 
            .CO(n53012));
    SB_LUT4 add_5427_9_lut (.I0(GND_net), .I1(n22501[6]), .I2(n621_adj_4587), 
            .I3(n53010), .O(n22177[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5436_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n53281));
    SB_CARRY add_5427_9 (.CI(n53010), .I0(n22501[6]), .I1(n621_adj_4587), 
            .CO(n53011));
    SB_LUT4 add_5427_8_lut (.I0(GND_net), .I1(n22501[5]), .I2(n548_adj_4588), 
            .I3(n53009), .O(n22177[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_12 (.CI(n53901), .I0(n11135[9]), .I1(n804), 
            .CO(n53902));
    SB_CARRY add_5427_8 (.CI(n53009), .I0(n22501[5]), .I1(n548_adj_4588), 
            .CO(n53010));
    SB_LUT4 add_5427_7_lut (.I0(GND_net), .I1(n22501[4]), .I2(n475_adj_4589), 
            .I3(n53008), .O(n22177[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4501));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n11135[8]), .I2(n731), 
            .I3(n53900), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_7 (.CI(n53008), .I0(n22501[4]), .I1(n475_adj_4589), 
            .CO(n53009));
    SB_LUT4 n71541_bdd_4_lut (.I0(n71541), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4749), .O(n71544));
    defparam n71541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5427_6_lut (.I0(GND_net), .I1(n22501[3]), .I2(n402_adj_4590), 
            .I3(n53007), .O(n22177[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_6 (.CI(n53007), .I0(n22501[3]), .I1(n402_adj_4590), 
            .CO(n53008));
    SB_CARRY mult_23_add_1221_11 (.CI(n53900), .I0(n11135[8]), .I1(n731), 
            .CO(n53901));
    SB_LUT4 add_5427_5_lut (.I0(GND_net), .I1(n22501[2]), .I2(n329_adj_4591), 
            .I3(n53006), .O(n22177[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5427_5 (.CI(n53006), .I0(n22501[2]), .I1(n329_adj_4591), 
            .CO(n53007));
    SB_LUT4 add_5427_4_lut (.I0(GND_net), .I1(n22501[1]), .I2(n256_adj_4592), 
            .I3(n53005), .O(n22177[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n11135[7]), .I2(n658), 
            .I3(n53899), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_10 (.CI(n53899), .I0(n11135[7]), .I1(n658), 
            .CO(n53900));
    SB_CARRY add_5427_4 (.CI(n53005), .I0(n22501[1]), .I1(n256_adj_4592), 
            .CO(n53006));
    SB_LUT4 add_5427_3_lut (.I0(GND_net), .I1(n22501[0]), .I2(n183_adj_4593), 
            .I3(n53004), .O(n22177[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n11135[6]), .I2(n585), 
            .I3(n53898), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_3 (.CI(n53004), .I0(n22501[0]), .I1(n183_adj_4593), 
            .CO(n53005));
    SB_LUT4 add_5427_2_lut (.I0(GND_net), .I1(n41_adj_4595), .I2(n110_adj_4596), 
            .I3(GND_net), .O(n22177[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5427_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5427_2 (.CI(GND_net), .I0(n41_adj_4595), .I1(n110_adj_4596), 
            .CO(n53004));
    SB_LUT4 add_5451_11_lut (.I0(GND_net), .I1(n22739[8]), .I2(n770), 
            .I3(n53003), .O(n22501[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n53898), .I0(n11135[6]), .I1(n585), 
            .CO(n53899));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n11135[5]), .I2(n512), 
            .I3(n53897), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5451_10_lut (.I0(GND_net), .I1(n22739[7]), .I2(n697), 
            .I3(n53002), .O(n22501[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_10 (.CI(n53002), .I0(n22739[7]), .I1(n697), .CO(n53003));
    SB_LUT4 add_5451_9_lut (.I0(GND_net), .I1(n22739[6]), .I2(n624), .I3(n53001), 
            .O(n22501[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_9 (.CI(n53001), .I0(n22739[6]), .I1(n624), .CO(n53002));
    SB_CARRY mult_23_add_1221_8 (.CI(n53897), .I0(n11135[5]), .I1(n512), 
            .CO(n53898));
    SB_LUT4 add_5451_8_lut (.I0(GND_net), .I1(n22739[5]), .I2(n551), .I3(n53000), 
            .O(n22501[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_8 (.CI(n53000), .I0(n22739[5]), .I1(n551), .CO(n53001));
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n11135[4]), .I2(n439), 
            .I3(n53896), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_7 (.CI(n53896), .I0(n11135[4]), .I1(n439), 
            .CO(n53897));
    SB_LUT4 add_5451_7_lut (.I0(GND_net), .I1(n22739[4]), .I2(n478_adj_4597), 
            .I3(n52999), .O(n22501[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_7 (.CI(n52999), .I0(n22739[4]), .I1(n478_adj_4597), 
            .CO(n53000));
    SB_LUT4 add_5451_6_lut (.I0(GND_net), .I1(n22739[3]), .I2(n405), .I3(n52998), 
            .O(n22501[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n11135[3]), .I2(n366), 
            .I3(n53895), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n53895), .I0(n11135[3]), .I1(n366), 
            .CO(n53896));
    SB_CARRY add_5451_6 (.CI(n52998), .I0(n22739[3]), .I1(n405), .CO(n52999));
    SB_LUT4 add_5451_5_lut (.I0(GND_net), .I1(n22739[2]), .I2(n332), .I3(n52997), 
            .O(n22501[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n11135[2]), .I2(n293_adj_4599), 
            .I3(n53894), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_5 (.CI(n52997), .I0(n22739[2]), .I1(n332), .CO(n52998));
    SB_CARRY mult_23_add_1221_5 (.CI(n53894), .I0(n11135[2]), .I1(n293_adj_4599), 
            .CO(n53895));
    SB_LUT4 add_5451_4_lut (.I0(GND_net), .I1(n22739[1]), .I2(n259), .I3(n52996), 
            .O(n22501[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_4 (.CI(n52996), .I0(n22739[1]), .I1(n259), .CO(n52997));
    SB_LUT4 add_5451_3_lut (.I0(GND_net), .I1(n22739[0]), .I2(n186), .I3(n52995), 
            .O(n22501[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_3 (.CI(n52995), .I0(n22739[0]), .I1(n186), .CO(n52996));
    SB_LUT4 add_5451_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n22501[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5451_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n11135[1]), .I2(n220), 
            .I3(n53893), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_4 (.CI(n53893), .I0(n11135[1]), .I1(n220), 
            .CO(n53894));
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4600));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n11135[0]), .I2(n147), 
            .I3(n53892), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5451_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n52995));
    SB_CARRY mult_23_add_1221_3 (.CI(n53892), .I0(n11135[0]), .I1(n147), 
            .CO(n53893));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5), .I2(n74_adj_4602), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5), .I1(n74_adj_4602), 
            .CO(n53892));
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n10676[0]), .I2(n10017[0]), 
            .I3(n52803), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4500));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n28[22]), 
            .I3(n52802), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n71550), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_25_24 (.CI(n52802), .I0(n360[22]), .I1(n28[22]), .CO(n52803));
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n28[21]), 
            .I3(n52801), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n52801), .I0(n360[21]), .I1(n28[21]), .CO(n52802));
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n71544), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n71532), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n71520), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n71514), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n71508), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n71502), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n71496), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n71490), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n71484), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n71478), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n71472), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n71466), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n71460), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n71454), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n71448), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n71442), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n71436), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n71430), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n71424), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n71418), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n71412), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n28[20]), 
            .I3(n52800), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n52800), .I0(n360[20]), .I1(n28[20]), .CO(n52801));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n28[19]), 
            .I3(n52799), .O(n455[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n52799), .I0(n360[19]), .I1(n28[19]), .CO(n52800));
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n28[18]), 
            .I3(n52798), .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n52798), .I0(n360[18]), .I1(n28[18]), .CO(n52799));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n28[17]), 
            .I3(n52797), .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n52797), .I0(n360[17]), .I1(n28[17]), .CO(n52798));
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n28[16]), 
            .I3(n52796), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n52796), .I0(n360[16]), .I1(n28[16]), .CO(n52797));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n28[15]), 
            .I3(n52795), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_17 (.CI(n52795), .I0(n360[15]), .I1(n28[15]), .CO(n52796));
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n28[14]), 
            .I3(n52794), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_16 (.CI(n52794), .I0(n360[14]), .I1(n28[14]), .CO(n52795));
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n28[13]), 
            .I3(n52793), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n52793), .I0(n360[13]), .I1(n28[13]), .CO(n52794));
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n28[12]), 
            .I3(n52792), .O(n455[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n52792), .I0(n360[12]), .I1(n28[12]), .CO(n52793));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n28[11]), 
            .I3(n52791), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n52791), .I0(n360[11]), .I1(n28[11]), .CO(n52792));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n28[10]), 
            .I3(n52790), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_12 (.CI(n52790), .I0(n360[10]), .I1(n28[10]), .CO(n52791));
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n335[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n28[9]), .I3(n52789), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_11 (.CI(n52789), .I0(n360[9]), .I1(n28[9]), .CO(n52790));
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4498));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51983 (.I0(n9977), .I1(n67734), .I2(setpoint[20]), 
            .I3(n4749), .O(n71529));
    defparam n9977_bdd_4_lut_51983.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71529_bdd_4_lut (.I0(n71529), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4749), .O(n71532));
    defparam n71529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4496));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4495));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51973 (.I0(n9977), .I1(n67733), .I2(setpoint[19]), 
            .I3(n4749), .O(n71517));
    defparam n9977_bdd_4_lut_51973.LUT_INIT = 16'he4aa;
    SB_LUT4 n71517_bdd_4_lut (.I0(n71517), .I1(n535[19]), .I2(n455[19]), 
            .I3(n4749), .O(n71520));
    defparam n71517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4609));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51964 (.I0(n9977), .I1(n67732), .I2(setpoint[18]), 
            .I3(n4749), .O(n71511));
    defparam n9977_bdd_4_lut_51964.LUT_INIT = 16'he4aa;
    SB_LUT4 n71511_bdd_4_lut (.I0(n71511), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4749), .O(n71514));
    defparam n71511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n233[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51959 (.I0(n9977), .I1(n67731), .I2(setpoint[17]), 
            .I3(n4749), .O(n71505));
    defparam n9977_bdd_4_lut_51959.LUT_INIT = 16'he4aa;
    SB_LUT4 n71505_bdd_4_lut (.I0(n71505), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4749), .O(n71508));
    defparam n71505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9977_bdd_4_lut_51954 (.I0(n9977), .I1(n67730), .I2(setpoint[16]), 
            .I3(n4749), .O(n71499));
    defparam n9977_bdd_4_lut_51954.LUT_INIT = 16'he4aa;
    SB_LUT4 n71499_bdd_4_lut (.I0(n71499), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4749), .O(n71502));
    defparam n71499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51949 (.I0(n9977), .I1(n67729), .I2(setpoint[15]), 
            .I3(n4749), .O(n71493));
    defparam n9977_bdd_4_lut_51949.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5459_11_lut (.I0(GND_net), .I1(n22816[8]), .I2(n770_adj_4612), 
            .I3(n53241), .O(n22597[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_23_lut (.I0(GND_net), .I1(n13103[20]), .I2(GND_net), 
            .I3(n53870), .O(n11135[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_22_lut (.I0(GND_net), .I1(n13103[19]), .I2(GND_net), 
            .I3(n53869), .O(n11135[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_22 (.CI(n53869), .I0(n13103[19]), .I1(GND_net), 
            .CO(n53870));
    SB_LUT4 add_5459_10_lut (.I0(GND_net), .I1(n22816[7]), .I2(n697_adj_4613), 
            .I3(n53240), .O(n22597[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_10 (.CI(n53240), .I0(n22816[7]), .I1(n697_adj_4613), 
            .CO(n53241));
    SB_LUT4 add_4659_21_lut (.I0(GND_net), .I1(n13103[18]), .I2(GND_net), 
            .I3(n53868), .O(n11135[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5459_9_lut (.I0(GND_net), .I1(n22816[6]), .I2(n624_adj_4614), 
            .I3(n53239), .O(n22597[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_9 (.CI(n53239), .I0(n22816[6]), .I1(n624_adj_4614), 
            .CO(n53240));
    SB_LUT4 add_5459_8_lut (.I0(GND_net), .I1(n22816[5]), .I2(n551_adj_4615), 
            .I3(n53238), .O(n22597[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_21 (.CI(n53868), .I0(n13103[18]), .I1(GND_net), 
            .CO(n53869));
    SB_CARRY add_5459_8 (.CI(n53238), .I0(n22816[5]), .I1(n551_adj_4615), 
            .CO(n53239));
    SB_LUT4 add_5459_7_lut (.I0(GND_net), .I1(n22816[4]), .I2(n478_adj_4616), 
            .I3(n53237), .O(n22597[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_20_lut (.I0(GND_net), .I1(n13103[17]), .I2(GND_net), 
            .I3(n53867), .O(n11135[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_7 (.CI(n53237), .I0(n22816[4]), .I1(n478_adj_4616), 
            .CO(n53238));
    SB_LUT4 add_5459_6_lut (.I0(GND_net), .I1(n22816[3]), .I2(n405_adj_4617), 
            .I3(n53236), .O(n22597[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_20 (.CI(n53867), .I0(n13103[17]), .I1(GND_net), 
            .CO(n53868));
    SB_CARRY add_5459_6 (.CI(n53236), .I0(n22816[3]), .I1(n405_adj_4617), 
            .CO(n53237));
    SB_LUT4 add_5459_5_lut (.I0(GND_net), .I1(n22816[2]), .I2(n332_adj_4618), 
            .I3(n53235), .O(n22597[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_19_lut (.I0(GND_net), .I1(n13103[16]), .I2(GND_net), 
            .I3(n53866), .O(n11135[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_5 (.CI(n53235), .I0(n22816[2]), .I1(n332_adj_4618), 
            .CO(n53236));
    SB_LUT4 add_5459_4_lut (.I0(GND_net), .I1(n22816[1]), .I2(n259_adj_4619), 
            .I3(n53234), .O(n22597[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_19 (.CI(n53866), .I0(n13103[16]), .I1(GND_net), 
            .CO(n53867));
    SB_CARRY add_5459_4 (.CI(n53234), .I0(n22816[1]), .I1(n259_adj_4619), 
            .CO(n53235));
    SB_LUT4 add_5459_3_lut (.I0(GND_net), .I1(n22816[0]), .I2(n186_adj_4620), 
            .I3(n53233), .O(n22597[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_18_lut (.I0(GND_net), .I1(n13103[15]), .I2(GND_net), 
            .I3(n53865), .O(n11135[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5459_3 (.CI(n53233), .I0(n22816[0]), .I1(n186_adj_4620), 
            .CO(n53234));
    SB_LUT4 add_5459_2_lut (.I0(GND_net), .I1(n44_adj_4621), .I2(n113_adj_4622), 
            .I3(GND_net), .O(n22597[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5459_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_18 (.CI(n53865), .I0(n13103[15]), .I1(GND_net), 
            .CO(n53866));
    SB_CARRY add_5459_2 (.CI(GND_net), .I0(n44_adj_4621), .I1(n113_adj_4622), 
            .CO(n53233));
    SB_LUT4 add_4659_17_lut (.I0(GND_net), .I1(n13103[14]), .I2(GND_net), 
            .I3(n53864), .O(n11135[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_17 (.CI(n53864), .I0(n13103[14]), .I1(GND_net), 
            .CO(n53865));
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4494));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4659_16_lut (.I0(GND_net), .I1(n13103[13]), .I2(n1099), 
            .I3(n53863), .O(n11135[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_16 (.CI(n53863), .I0(n13103[13]), .I1(n1099), .CO(n53864));
    SB_LUT4 add_4659_15_lut (.I0(GND_net), .I1(n13103[12]), .I2(n1026), 
            .I3(n53862), .O(n11135[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n335[23]), .I1(n10524[21]), .I2(GND_net), 
            .I3(n53232), .O(n10017[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n10524[20]), .I2(GND_net), 
            .I3(n53231), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_23 (.CI(n53231), .I0(n10524[20]), .I1(GND_net), 
            .CO(n53232));
    SB_CARRY add_4659_15 (.CI(n53862), .I0(n13103[12]), .I1(n1026), .CO(n53863));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n10524[19]), .I2(GND_net), 
            .I3(n53230), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_14_lut (.I0(GND_net), .I1(n13103[11]), .I2(n953), 
            .I3(n53861), .O(n11135[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_22 (.CI(n53230), .I0(n10524[19]), .I1(GND_net), 
            .CO(n53231));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n10524[18]), .I2(GND_net), 
            .I3(n53229), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_14 (.CI(n53861), .I0(n13103[11]), .I1(n953), .CO(n53862));
    SB_CARRY mult_24_add_1225_21 (.CI(n53229), .I0(n10524[18]), .I1(GND_net), 
            .CO(n53230));
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n10524[17]), .I2(GND_net), 
            .I3(n53228), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_13_lut (.I0(GND_net), .I1(n13103[10]), .I2(n880), 
            .I3(n53860), .O(n11135[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n53228), .I0(n10524[17]), .I1(GND_net), 
            .CO(n53229));
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n10524[16]), .I2(GND_net), 
            .I3(n53227), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_13 (.CI(n53860), .I0(n13103[10]), .I1(n880), .CO(n53861));
    SB_CARRY mult_24_add_1225_19 (.CI(n53227), .I0(n10524[16]), .I1(GND_net), 
            .CO(n53228));
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n10524[15]), .I2(GND_net), 
            .I3(n53226), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_12_lut (.I0(GND_net), .I1(n13103[9]), .I2(n807), 
            .I3(n53859), .O(n11135[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_18 (.CI(n53226), .I0(n10524[15]), .I1(GND_net), 
            .CO(n53227));
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n10524[14]), .I2(GND_net), 
            .I3(n53225), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_12 (.CI(n53859), .I0(n13103[9]), .I1(n807), .CO(n53860));
    SB_CARRY mult_24_add_1225_17 (.CI(n53225), .I0(n10524[14]), .I1(GND_net), 
            .CO(n53226));
    SB_LUT4 add_4659_11_lut (.I0(GND_net), .I1(n13103[8]), .I2(n734), 
            .I3(n53858), .O(n11135[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_11 (.CI(n53858), .I0(n13103[8]), .I1(n734), .CO(n53859));
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n10524[13]), .I2(n1096_adj_4623), 
            .I3(n53224), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_10_lut (.I0(GND_net), .I1(n13103[7]), .I2(n661), 
            .I3(n53857), .O(n11135[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_16 (.CI(n53224), .I0(n10524[13]), .I1(n1096_adj_4623), 
            .CO(n53225));
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n10524[12]), .I2(n1023_adj_4624), 
            .I3(n53223), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_10 (.CI(n53857), .I0(n13103[7]), .I1(n661), .CO(n53858));
    SB_CARRY mult_24_add_1225_15 (.CI(n53223), .I0(n10524[12]), .I1(n1023_adj_4624), 
            .CO(n53224));
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n10524[11]), .I2(n950_adj_4625), 
            .I3(n53222), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_9_lut (.I0(GND_net), .I1(n13103[6]), .I2(n588), .I3(n53856), 
            .O(n11135[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_14 (.CI(n53222), .I0(n10524[11]), .I1(n950_adj_4625), 
            .CO(n53223));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n10524[10]), .I2(n877_adj_4626), 
            .I3(n53221), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_9 (.CI(n53856), .I0(n13103[6]), .I1(n588), .CO(n53857));
    SB_CARRY mult_24_add_1225_13 (.CI(n53221), .I0(n10524[10]), .I1(n877_adj_4626), 
            .CO(n53222));
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n10524[9]), .I2(n804_adj_4627), 
            .I3(n53220), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71493_bdd_4_lut (.I0(n71493), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4749), .O(n71496));
    defparam n71493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_24_add_1225_12 (.CI(n53220), .I0(n10524[9]), .I1(n804_adj_4627), 
            .CO(n53221));
    SB_LUT4 add_4659_8_lut (.I0(GND_net), .I1(n13103[5]), .I2(n515), .I3(n53855), 
            .O(n11135[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4493));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4659_8 (.CI(n53855), .I0(n13103[5]), .I1(n515), .CO(n53856));
    SB_LUT4 add_4659_7_lut (.I0(GND_net), .I1(n13103[4]), .I2(n442_adj_4629), 
            .I3(n53854), .O(n11135[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n10524[8]), .I2(n731_adj_4630), 
            .I3(n53219), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_7 (.CI(n53854), .I0(n13103[4]), .I1(n442_adj_4629), 
            .CO(n53855));
    SB_CARRY mult_24_add_1225_11 (.CI(n53219), .I0(n10524[8]), .I1(n731_adj_4630), 
            .CO(n53220));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n10524[7]), .I2(n658_adj_4631), 
            .I3(n53218), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n28[8]), .I3(n52788), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n53218), .I0(n10524[7]), .I1(n658_adj_4631), 
            .CO(n53219));
    SB_LUT4 add_4659_6_lut (.I0(GND_net), .I1(n13103[3]), .I2(n369), .I3(n53853), 
            .O(n11135[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n10524[6]), .I2(n585_adj_4632), 
            .I3(n53217), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_9 (.CI(n53217), .I0(n10524[6]), .I1(n585_adj_4632), 
            .CO(n53218));
    SB_CARRY add_25_10 (.CI(n52788), .I0(n360[8]), .I1(n28[8]), .CO(n52789));
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4550));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4659_6 (.CI(n53853), .I0(n13103[3]), .I1(n369), .CO(n53854));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n10524[5]), .I2(n512_adj_4633), 
            .I3(n53216), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n53216), .I0(n10524[5]), .I1(n512_adj_4633), 
            .CO(n53217));
    SB_LUT4 add_4659_5_lut (.I0(GND_net), .I1(n13103[2]), .I2(n296), .I3(n53852), 
            .O(n11135[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n10524[4]), .I2(n439_adj_4634), 
            .I3(n53215), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n28[7]), .I3(n52787), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4636));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_24_add_1225_7 (.CI(n53215), .I0(n10524[4]), .I1(n439_adj_4634), 
            .CO(n53216));
    SB_CARRY add_25_9 (.CI(n52787), .I0(n360[7]), .I1(n28[7]), .CO(n52788));
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n28[6]), .I3(n52786), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i11_3_lut (.I0(n233[10]), .I1(n285[10]), .I2(n284), 
            .I3(GND_net), .O(n310[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i11_3_lut (.I0(n310[10]), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n335[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n10524[3]), .I2(n366_adj_4637), 
            .I3(n53214), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_5 (.CI(n53852), .I0(n13103[2]), .I1(n296), .CO(n53853));
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4549));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_6 (.CI(n53214), .I0(n10524[3]), .I1(n366_adj_4637), 
            .CO(n53215));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n10524[2]), .I2(n293_adj_4638), 
            .I3(n53213), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_4_lut (.I0(GND_net), .I1(n13103[1]), .I2(n223_adj_4639), 
            .I3(n53851), .O(n11135[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_5 (.CI(n53213), .I0(n10524[2]), .I1(n293_adj_4638), 
            .CO(n53214));
    SB_CARRY add_4659_4 (.CI(n53851), .I0(n13103[1]), .I1(n223_adj_4639), 
            .CO(n53852));
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4548));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n10524[1]), .I2(n220_adj_4640), 
            .I3(n53212), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_4 (.CI(n53212), .I0(n10524[1]), .I1(n220_adj_4640), 
            .CO(n53213));
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n10524[0]), .I2(n147_adj_4641), 
            .I3(n53211), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4547));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_25_8 (.CI(n52786), .I0(n360[6]), .I1(n28[6]), .CO(n52787));
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4659_3_lut (.I0(GND_net), .I1(n13103[0]), .I2(n150), .I3(n53850), 
            .O(n11135[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_3 (.CI(n53850), .I0(n13103[0]), .I1(n150), .CO(n53851));
    SB_CARRY mult_24_add_1225_3 (.CI(n53211), .I0(n10524[0]), .I1(n147_adj_4641), 
            .CO(n53212));
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4642), .I2(n74_adj_4643), 
            .I3(GND_net), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4659_2_lut (.I0(GND_net), .I1(n8_adj_4644), .I2(n77), 
            .I3(GND_net), .O(n11135[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4659_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5_adj_4642), .I1(n74_adj_4643), 
            .CO(n53211));
    SB_LUT4 add_4511_23_lut (.I0(GND_net), .I1(n12531[20]), .I2(GND_net), 
            .I3(n53210), .O(n10524[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4659_2 (.CI(GND_net), .I0(n8_adj_4644), .I1(n77), .CO(n53850));
    SB_LUT4 add_4511_22_lut (.I0(GND_net), .I1(n12531[19]), .I2(GND_net), 
            .I3(n53209), .O(n10524[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[23]), 
            .I3(n52949), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_22 (.CI(n53209), .I0(n12531[19]), .I1(GND_net), 
            .CO(n53210));
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[22]), 
            .I3(n52948), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n52948), .I0(GND_net), .I1(n1_adj_5019[22]), 
            .CO(n52949));
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n28[5]), .I3(n52785), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_22_lut (.I0(GND_net), .I1(n14630[19]), .I2(GND_net), 
            .I3(n53849), .O(n13103[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_21_lut (.I0(GND_net), .I1(n12531[18]), .I2(GND_net), 
            .I3(n53208), .O(n10524[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[21]), 
            .I3(n52947), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_23 (.CI(n52947), .I0(GND_net), .I1(n1_adj_5019[21]), 
            .CO(n52948));
    SB_CARRY add_4511_21 (.CI(n53208), .I0(n12531[18]), .I1(GND_net), 
            .CO(n53209));
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[20]), 
            .I3(n52946), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n52946), .I0(GND_net), .I1(n1_adj_5019[20]), 
            .CO(n52947));
    SB_CARRY add_25_7 (.CI(n52785), .I0(n360[5]), .I1(n28[5]), .CO(n52786));
    SB_LUT4 add_4982_21_lut (.I0(GND_net), .I1(n14630[18]), .I2(GND_net), 
            .I3(n53848), .O(n13103[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_20_lut (.I0(GND_net), .I1(n12531[17]), .I2(GND_net), 
            .I3(n53207), .O(n10524[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[19]), 
            .I3(n52945), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n52945), .I0(GND_net), .I1(n1_adj_5019[19]), 
            .CO(n52946));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n28[4]), .I3(n52784), 
            .O(n455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[18]), 
            .I3(n52944), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n52784), .I0(n360[4]), .I1(n28[4]), .CO(n52785));
    SB_CARRY add_4511_20 (.CI(n53207), .I0(n12531[17]), .I1(GND_net), 
            .CO(n53208));
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4492));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4511_19_lut (.I0(GND_net), .I1(n12531[16]), .I2(GND_net), 
            .I3(n53206), .O(n10524[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_20 (.CI(n52944), .I0(GND_net), .I1(n1_adj_5019[18]), 
            .CO(n52945));
    SB_CARRY add_4982_21 (.CI(n53848), .I0(n14630[18]), .I1(GND_net), 
            .CO(n53849));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[17]), 
            .I3(n52943), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n52943), .I0(GND_net), .I1(n1_adj_5019[17]), 
            .CO(n52944));
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n335[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n28[3]), .I3(n52783), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4491));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[16]), 
            .I3(n52942), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4489));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4982_20_lut (.I0(GND_net), .I1(n14630[17]), .I2(GND_net), 
            .I3(n53847), .O(n13103[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4488));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_25_5 (.CI(n52783), .I0(n360[3]), .I1(n28[3]), .CO(n52784));
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4544));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4982_20 (.CI(n53847), .I0(n14630[17]), .I1(GND_net), 
            .CO(n53848));
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4543));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4982_19_lut (.I0(GND_net), .I1(n14630[16]), .I2(GND_net), 
            .I3(n53846), .O(n13103[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_19 (.CI(n53206), .I0(n12531[16]), .I1(GND_net), 
            .CO(n53207));
    SB_CARRY unary_minus_33_add_3_18 (.CI(n52942), .I0(GND_net), .I1(n1_adj_5019[16]), 
            .CO(n52943));
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[15]), 
            .I3(n52941), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n28[2]), .I3(n52782), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_4 (.CI(n52782), .I0(n360[2]), .I1(n28[2]), .CO(n52783));
    SB_LUT4 add_4511_18_lut (.I0(GND_net), .I1(n12531[15]), .I2(GND_net), 
            .I3(n53205), .O(n10524[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_17 (.CI(n52941), .I0(GND_net), .I1(n1_adj_5019[15]), 
            .CO(n52942));
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[14]), 
            .I3(n52940), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n28[1]), .I3(n52781), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_3 (.CI(n52781), .I0(n360[1]), .I1(n28[1]), .CO(n52782));
    SB_CARRY add_4982_19 (.CI(n53846), .I0(n14630[16]), .I1(GND_net), 
            .CO(n53847));
    SB_LUT4 add_4982_18_lut (.I0(GND_net), .I1(n14630[15]), .I2(GND_net), 
            .I3(n53845), .O(n13103[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_18 (.CI(n53205), .I0(n12531[15]), .I1(GND_net), 
            .CO(n53206));
    SB_CARRY unary_minus_33_add_3_16 (.CI(n52940), .I0(GND_net), .I1(n1_adj_5019[14]), 
            .CO(n52941));
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4541));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n207[23]), .I1(\Kp[2] ), .I2(n52458), 
            .I3(n207[22]), .O(n64059));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[13]), 
            .I3(n52939), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n28[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n28[0]), .CO(n52781));
    SB_CARRY add_4982_18 (.CI(n53845), .I0(n14630[15]), .I1(GND_net), 
            .CO(n53846));
    SB_LUT4 add_4982_17_lut (.I0(GND_net), .I1(n14630[14]), .I2(GND_net), 
            .I3(n53844), .O(n13103[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_17_lut (.I0(GND_net), .I1(n12531[14]), .I2(GND_net), 
            .I3(n53204), .O(n10524[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_15 (.CI(n52939), .I0(GND_net), .I1(n1_adj_5019[13]), 
            .CO(n52940));
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[12]), 
            .I3(n52938), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n52780), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n52779), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4540));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4486));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4982_17 (.CI(n53844), .I0(n14630[14]), .I1(GND_net), 
            .CO(n53845));
    SB_LUT4 i1_4_lut_adj_951 (.I0(n207[22]), .I1(n23335[1]), .I2(n4_adj_4652), 
            .I3(\Kp[3] ), .O(n23287[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4485));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_952 (.I0(n23335[1]), .I1(n6_adj_4653), .I2(n347), 
            .I3(n60165), .O(n23287[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4539));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34557_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n52458));   // verilog/motorControl.v(61[20:26])
    defparam i34557_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(n64055), .I1(n207[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4652));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4538));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34626_4_lut (.I0(n23335[1]), .I1(\Kp[3] ), .I2(n4_adj_4652), 
            .I3(n207[22]), .O(n6_adj_4653));   // verilog/motorControl.v(61[20:26])
    defparam i34626_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_23_i46_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_4654));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i46_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4511_17 (.CI(n53204), .I0(n12531[14]), .I1(GND_net), 
            .CO(n53205));
    SB_CARRY unary_minus_33_add_3_14 (.CI(n52938), .I0(GND_net), .I1(n1_adj_5019[12]), 
            .CO(n52939));
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[11]), 
            .I3(n52937), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_24 (.CI(n52779), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n52780));
    SB_LUT4 add_4511_16_lut (.I0(GND_net), .I1(n12531[13]), .I2(n1099_adj_4656), 
            .I3(n53203), .O(n10524[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_16 (.CI(n53203), .I0(n12531[13]), .I1(n1099_adj_4656), 
            .CO(n53204));
    SB_LUT4 add_4511_15_lut (.I0(GND_net), .I1(n12531[12]), .I2(n1026_adj_4657), 
            .I3(n53202), .O(n10524[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n52937), .I0(GND_net), .I1(n1_adj_5019[11]), 
            .CO(n52938));
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n32594), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n52778), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_16_lut (.I0(GND_net), .I1(n14630[13]), .I2(n1102), 
            .I3(n53843), .O(n13103[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n32593), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n32592), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n32591), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n32590), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n32589), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n32588), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n32587), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n32586), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n32585), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n32584), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n32583), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n32582), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n32581), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n32580), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n32579), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n32578), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n32577), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n32576), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n32575), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n32574), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n32573), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n32570), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n9977_bdd_4_lut_51944 (.I0(n9977), .I1(n67728), .I2(setpoint[14]), 
            .I3(n4749), .O(n71487));
    defparam n9977_bdd_4_lut_51944.LUT_INIT = 16'he4aa;
    SB_CARRY add_4511_15 (.CI(n53202), .I0(n12531[12]), .I1(n1026_adj_4657), 
            .CO(n53203));
    SB_LUT4 add_4511_14_lut (.I0(GND_net), .I1(n12531[11]), .I2(n953_adj_4658), 
            .I3(n53201), .O(n10524[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_23 (.CI(n52778), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n52779));
    SB_CARRY add_4511_14 (.CI(n53201), .I0(n12531[11]), .I1(n953_adj_4658), 
            .CO(n53202));
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[10]), 
            .I3(n52936), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_12 (.CI(n52936), .I0(GND_net), .I1(n1_adj_5019[10]), 
            .CO(n52937));
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[9]), 
            .I3(n52935), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n52777), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_16 (.CI(n53843), .I0(n14630[13]), .I1(n1102), .CO(n53844));
    SB_LUT4 add_4511_13_lut (.I0(GND_net), .I1(n12531[10]), .I2(n880_adj_4659), 
            .I3(n53200), .O(n10524[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_11 (.CI(n52935), .I0(GND_net), .I1(n1_adj_5019[9]), 
            .CO(n52936));
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[8]), 
            .I3(n52934), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_22 (.CI(n52777), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n52778));
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n52776), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_15_lut (.I0(GND_net), .I1(n14630[12]), .I2(n1029), 
            .I3(n53842), .O(n13103[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_13 (.CI(n53200), .I0(n12531[10]), .I1(n880_adj_4659), 
            .CO(n53201));
    SB_CARRY unary_minus_33_add_3_10 (.CI(n52934), .I0(GND_net), .I1(n1_adj_5019[8]), 
            .CO(n52935));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[7]), 
            .I3(n52933), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n52776), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n52777));
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n52775), .O(n233[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_12_lut (.I0(GND_net), .I1(n12531[9]), .I2(n807_adj_4662), 
            .I3(n53199), .O(n10524[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n52933), .I0(GND_net), .I1(n1_adj_5019[7]), 
            .CO(n52934));
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[6]), 
            .I3(n52932), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_20 (.CI(n52775), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n52776));
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n52774), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_15 (.CI(n53842), .I0(n14630[12]), .I1(n1029), .CO(n53843));
    SB_CARRY add_16_19 (.CI(n52774), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n52775));
    SB_LUT4 add_4982_14_lut (.I0(GND_net), .I1(n14630[11]), .I2(n956), 
            .I3(n53841), .O(n13103[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_14 (.CI(n53841), .I0(n14630[11]), .I1(n956), .CO(n53842));
    SB_CARRY add_4511_12 (.CI(n53199), .I0(n12531[9]), .I1(n807_adj_4662), 
            .CO(n53200));
    SB_CARRY unary_minus_33_add_3_8 (.CI(n52932), .I0(GND_net), .I1(n1_adj_5019[6]), 
            .CO(n52933));
    SB_LUT4 add_4511_11_lut (.I0(GND_net), .I1(n12531[8]), .I2(n734_adj_4664), 
            .I3(n53198), .O(n10524[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[5]), 
            .I3(n52931), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n52773), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n52931), .I0(GND_net), .I1(n1_adj_5019[5]), 
            .CO(n52932));
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4537));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_18 (.CI(n52773), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n52774));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n52772), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_13_lut (.I0(GND_net), .I1(n14630[10]), .I2(n883), 
            .I3(n53840), .O(n13103[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_11 (.CI(n53198), .I0(n12531[8]), .I1(n734_adj_4664), 
            .CO(n53199));
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4536));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n64055));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i44888_3_lut (.I0(n207[23]), .I1(n64055), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n60165));   // verilog/motorControl.v(61[20:26])
    defparam i44888_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[4]), 
            .I3(n52930), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34566_3_lut (.I0(n207[23]), .I1(n52453), .I2(n54083), .I3(GND_net), 
            .O(n23335[1]));   // verilog/motorControl.v(61[20:26])
    defparam i34566_3_lut.LUT_INIT = 16'h6c6c;
    SB_CARRY add_4982_13 (.CI(n53840), .I0(n14630[10]), .I1(n883), .CO(n53841));
    SB_CARRY add_16_17 (.CI(n52772), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n52773));
    SB_LUT4 add_4982_12_lut (.I0(GND_net), .I1(n14630[9]), .I2(n810), 
            .I3(n53839), .O(n13103[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_10_lut (.I0(GND_net), .I1(n12531[7]), .I2(n661_adj_4668), 
            .I3(n53197), .O(n10524[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_6 (.CI(n52930), .I0(GND_net), .I1(n1_adj_5019[4]), 
            .CO(n52931));
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[3]), 
            .I3(n52929), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n52771), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_16 (.CI(n52771), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n52772));
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4535));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4982_12 (.CI(n53839), .I0(n14630[9]), .I1(n810), .CO(n53840));
    SB_CARRY add_4511_10 (.CI(n53197), .I0(n12531[7]), .I1(n661_adj_4668), 
            .CO(n53198));
    SB_CARRY unary_minus_33_add_3_5 (.CI(n52929), .I0(GND_net), .I1(n1_adj_5019[3]), 
            .CO(n52930));
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[2]), 
            .I3(n52928), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_9_lut (.I0(GND_net), .I1(n12531[6]), .I2(n588_adj_4670), 
            .I3(n53196), .O(n10524[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_4 (.CI(n52928), .I0(GND_net), .I1(n1_adj_5019[2]), 
            .CO(n52929));
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[1]), 
            .I3(n52927), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4534));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4982_11_lut (.I0(GND_net), .I1(n14630[8]), .I2(n737), 
            .I3(n53838), .O(n13103[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_9 (.CI(n53196), .I0(n12531[6]), .I1(n588_adj_4670), 
            .CO(n53197));
    SB_CARRY unary_minus_33_add_3_3 (.CI(n52927), .I0(GND_net), .I1(n1_adj_5019[1]), 
            .CO(n52928));
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5019[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_8_lut (.I0(GND_net), .I1(n12531[5]), .I2(n515_adj_4672), 
            .I3(n53195), .O(n10524[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_11 (.CI(n53838), .I0(n14630[8]), .I1(n737), .CO(n53839));
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5019[0]), 
            .CO(n52927));
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_5020[23]), 
            .I3(n52926), .O(n47_adj_4673)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_953 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n54083), 
            .I3(n207[22]), .O(n64045));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'hc60a;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4511_8 (.CI(n53195), .I0(n12531[5]), .I1(n515_adj_4672), 
            .CO(n53196));
    SB_LUT4 add_4982_10_lut (.I0(GND_net), .I1(n14630[7]), .I2(n664), 
            .I3(n53837), .O(n13103[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_rep_239_2_lut (.I0(n23335[1]), .I1(n60165), .I2(GND_net), 
            .I3(GND_net), .O(n71973));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_239_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_954 (.I0(n52453), .I1(n64045), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n64049));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_954.LUT_INIT = 16'h9666;
    SB_CARRY add_4982_10 (.CI(n53837), .I0(n14630[7]), .I1(n664), .CO(n53838));
    SB_LUT4 i34634_4_lut (.I0(n71973), .I1(\Kp[4] ), .I2(n6_adj_4653), 
            .I3(n207[22]), .O(n8_adj_4675));   // verilog/motorControl.v(61[20:26])
    defparam i34634_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4511_7_lut (.I0(GND_net), .I1(n12531[4]), .I2(n442_adj_4676), 
            .I3(n53194), .O(n10524[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n335[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4532));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[22]), 
            .I3(n52925), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34580_4_lut (.I0(n23335[1]), .I1(\Kp[3] ), .I2(n64055), .I3(n207[23]), 
            .O(n6_adj_4678));   // verilog/motorControl.v(61[20:26])
    defparam i34580_4_lut.LUT_INIT = 16'he800;
    SB_DFFSR counter_2045_2046__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 i1_4_lut_adj_955 (.I0(n6_adj_4678), .I1(n8_adj_4675), .I2(n64049), 
            .I3(n60165), .O(n62834));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_DFFSR counter_2045_2046__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY unary_minus_27_add_3_24 (.CI(n52925), .I0(GND_net), .I1(n1_adj_5020[22]), 
            .CO(n52926));
    SB_CARRY add_4511_7 (.CI(n53194), .I0(n12531[4]), .I1(n442_adj_4676), 
            .CO(n53195));
    SB_LUT4 add_4982_9_lut (.I0(GND_net), .I1(n14630[6]), .I2(n591), .I3(n53836), 
            .O(n13103[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_9 (.CI(n53836), .I0(n14630[6]), .I1(n591), .CO(n53837));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[21]), 
            .I3(n52924), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n52924), .I0(GND_net), .I1(n1_adj_5020[21]), 
            .CO(n52925));
    SB_LUT4 add_4511_6_lut (.I0(GND_net), .I1(n12531[3]), .I2(n369_adj_4681), 
            .I3(n53193), .O(n10524[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n52770), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[20]), 
            .I3(n52923), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_15 (.CI(n52770), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n52771));
    SB_LUT4 add_4982_8_lut (.I0(GND_net), .I1(n14630[5]), .I2(n518), .I3(n53835), 
            .O(n13103[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_6 (.CI(n53193), .I0(n12531[3]), .I1(n369_adj_4681), 
            .CO(n53194));
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n31682), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_27_add_3_22 (.CI(n52923), .I0(GND_net), .I1(n1_adj_5020[20]), 
            .CO(n52924));
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[19]), 
            .I3(n52922), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_8 (.CI(n53835), .I0(n14630[5]), .I1(n518), .CO(n53836));
    SB_LUT4 add_4982_7_lut (.I0(GND_net), .I1(n14630[4]), .I2(n445_adj_4684), 
            .I3(n53834), .O(n13103[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_5_lut (.I0(GND_net), .I1(n12531[2]), .I2(n296_adj_4685), 
            .I3(n53192), .O(n10524[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_21 (.CI(n52922), .I0(GND_net), .I1(n1_adj_5020[19]), 
            .CO(n52923));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[18]), 
            .I3(n52921), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n52769), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_7 (.CI(n53834), .I0(n14630[4]), .I1(n445_adj_4684), 
            .CO(n53835));
    SB_LUT4 add_4982_6_lut (.I0(GND_net), .I1(n14630[3]), .I2(n372), .I3(n53833), 
            .O(n13103[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_6 (.CI(n53833), .I0(n14630[3]), .I1(n372), .CO(n53834));
    SB_CARRY add_4511_5 (.CI(n53192), .I0(n12531[2]), .I1(n296_adj_4685), 
            .CO(n53193));
    SB_CARRY unary_minus_27_add_3_20 (.CI(n52921), .I0(GND_net), .I1(n1_adj_5020[18]), 
            .CO(n52922));
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[17]), 
            .I3(n52920), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_4_lut (.I0(GND_net), .I1(n12531[1]), .I2(n223_adj_4689), 
            .I3(n53191), .O(n10524[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n52920), .I0(GND_net), .I1(n1_adj_5020[17]), 
            .CO(n52921));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[16]), 
            .I3(n52919), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_5_lut (.I0(GND_net), .I1(n14630[2]), .I2(n299_adj_4691), 
            .I3(n53832), .O(n13103[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4511_4 (.CI(n53191), .I0(n12531[1]), .I1(n223_adj_4689), 
            .CO(n53192));
    SB_CARRY unary_minus_27_add_3_18 (.CI(n52919), .I0(GND_net), .I1(n1_adj_5020[16]), 
            .CO(n52920));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[15]), 
            .I3(n52918), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4511_3_lut (.I0(GND_net), .I1(n12531[0]), .I2(n150_adj_4694), 
            .I3(n53190), .O(n10524[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_5 (.CI(n53832), .I0(n14630[2]), .I1(n299_adj_4691), 
            .CO(n53833));
    SB_CARRY add_4511_3 (.CI(n53190), .I0(n12531[0]), .I1(n150_adj_4694), 
            .CO(n53191));
    SB_CARRY unary_minus_27_add_3_17 (.CI(n52918), .I0(GND_net), .I1(n1_adj_5020[15]), 
            .CO(n52919));
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[14]), 
            .I3(n52917), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_4_lut (.I0(GND_net), .I1(n14630[1]), .I2(n226_adj_4696), 
            .I3(n53831), .O(n13103[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n52917), .I0(GND_net), .I1(n1_adj_5020[14]), 
            .CO(n52918));
    SB_LUT4 add_4511_2_lut (.I0(GND_net), .I1(n8_adj_4697), .I2(n77_adj_4698), 
            .I3(GND_net), .O(n10524[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4511_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_14 (.CI(n52769), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n52770));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[13]), 
            .I3(n52916), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_15 (.CI(n52916), .I0(GND_net), .I1(n1_adj_5020[13]), 
            .CO(n52917));
    SB_CARRY add_4511_2 (.CI(GND_net), .I0(n8_adj_4697), .I1(n77_adj_4698), 
            .CO(n53190));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[12]), 
            .I3(n52915), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n52915), .I0(GND_net), .I1(n1_adj_5020[12]), 
            .CO(n52916));
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n52768), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_4 (.CI(n53831), .I0(n14630[1]), .I1(n226_adj_4696), 
            .CO(n53832));
    SB_LUT4 add_4982_3_lut (.I0(GND_net), .I1(n14630[0]), .I2(n153), .I3(n53830), 
            .O(n13103[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_22_lut (.I0(GND_net), .I1(n14124[19]), .I2(GND_net), 
            .I3(n53189), .O(n12531[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[11]), 
            .I3(n52914), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_13 (.CI(n52914), .I0(GND_net), .I1(n1_adj_5020[11]), 
            .CO(n52915));
    SB_LUT4 add_4957_21_lut (.I0(GND_net), .I1(n14124[18]), .I2(GND_net), 
            .I3(n53188), .O(n12531[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[10]), 
            .I3(n52913), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n52913), .I0(GND_net), .I1(n1_adj_5020[10]), 
            .CO(n52914));
    SB_CARRY add_16_13 (.CI(n52768), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n52769));
    SB_CARRY add_4982_3 (.CI(n53830), .I0(n14630[0]), .I1(n153), .CO(n53831));
    SB_CARRY add_4957_21 (.CI(n53188), .I0(n14124[18]), .I1(GND_net), 
            .CO(n53189));
    SB_LUT4 add_4957_20_lut (.I0(GND_net), .I1(n14124[17]), .I2(GND_net), 
            .I3(n53187), .O(n12531[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[9]), 
            .I3(n52912), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n52767), .O(n233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4982_2_lut (.I0(GND_net), .I1(n11_adj_4704), .I2(n80), 
            .I3(GND_net), .O(n13103[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4982_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_20 (.CI(n53187), .I0(n14124[17]), .I1(GND_net), 
            .CO(n53188));
    SB_CARRY unary_minus_27_add_3_11 (.CI(n52912), .I0(GND_net), .I1(n1_adj_5020[9]), 
            .CO(n52913));
    SB_CARRY add_16_12 (.CI(n52767), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n52768));
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n52766), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[8]), 
            .I3(n52911), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n52911), .I0(GND_net), .I1(n1_adj_5020[8]), 
            .CO(n52912));
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[7]), 
            .I3(n52910), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n52766), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n52767));
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n52765), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_19_lut (.I0(GND_net), .I1(n14124[16]), .I2(GND_net), 
            .I3(n53186), .O(n12531[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n52910), .I0(GND_net), .I1(n1_adj_5020[7]), 
            .CO(n52911));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[6]), 
            .I3(n52909), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_10 (.CI(n52765), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n52766));
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n52764), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4982_2 (.CI(GND_net), .I0(n11_adj_4704), .I1(n80), .CO(n53830));
    SB_CARRY add_4957_19 (.CI(n53186), .I0(n14124[16]), .I1(GND_net), 
            .CO(n53187));
    SB_CARRY unary_minus_27_add_3_8 (.CI(n52909), .I0(GND_net), .I1(n1_adj_5020[6]), 
            .CO(n52910));
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[5]), 
            .I3(n52908), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_18_lut (.I0(GND_net), .I1(n14124[15]), .I2(GND_net), 
            .I3(n53185), .O(n12531[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n52908), .I0(GND_net), .I1(n1_adj_5020[5]), 
            .CO(n52909));
    SB_CARRY add_16_9 (.CI(n52764), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n52765));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n52763), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_18 (.CI(n53185), .I0(n14124[15]), .I1(GND_net), 
            .CO(n53186));
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[4]), 
            .I3(n52907), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_21_lut (.I0(GND_net), .I1(n16003[18]), .I2(GND_net), 
            .I3(n53829), .O(n14630[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_20_lut (.I0(GND_net), .I1(n16003[17]), .I2(GND_net), 
            .I3(n53828), .O(n14630[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_6 (.CI(n52907), .I0(GND_net), .I1(n1_adj_5020[4]), 
            .CO(n52908));
    SB_CARRY add_16_8 (.CI(n52763), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n52764));
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n52762), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_20 (.CI(n53828), .I0(n16003[17]), .I1(GND_net), 
            .CO(n53829));
    SB_LUT4 add_5045_19_lut (.I0(GND_net), .I1(n16003[16]), .I2(GND_net), 
            .I3(n53827), .O(n14630[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_17_lut (.I0(GND_net), .I1(n14124[14]), .I2(GND_net), 
            .I3(n53184), .O(n12531[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[3]), 
            .I3(n52906), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n52906), .I0(GND_net), .I1(n1_adj_5020[3]), 
            .CO(n52907));
    SB_CARRY add_16_7 (.CI(n52762), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n52763));
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4531));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n52761), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_19 (.CI(n53827), .I0(n16003[16]), .I1(GND_net), 
            .CO(n53828));
    SB_LUT4 add_5045_18_lut (.I0(GND_net), .I1(n16003[15]), .I2(GND_net), 
            .I3(n53826), .O(n14630[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_17 (.CI(n53184), .I0(n14124[14]), .I1(GND_net), 
            .CO(n53185));
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[2]), 
            .I3(n52905), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_4 (.CI(n52905), .I0(GND_net), .I1(n1_adj_5020[2]), 
            .CO(n52906));
    SB_CARRY add_16_6 (.CI(n52761), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n52762));
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n52760), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_18 (.CI(n53826), .I0(n16003[15]), .I1(GND_net), 
            .CO(n53827));
    SB_LUT4 add_4957_16_lut (.I0(GND_net), .I1(n14124[13]), .I2(n1102_adj_4715), 
            .I3(n53183), .O(n12531[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5020[1]), 
            .I3(n52904), .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n52904), .I0(GND_net), .I1(n1_adj_5020[1]), 
            .CO(n52905));
    SB_CARRY add_16_5 (.CI(n52760), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n52761));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n52759), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_16 (.CI(n53183), .I0(n14124[13]), .I1(n1102_adj_4715), 
            .CO(n53184));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n41203), .I1(GND_net), .I2(n1_adj_5020[0]), 
            .I3(VCC_net), .O(n67585)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5020[0]), 
            .CO(n52904));
    SB_CARRY add_16_4 (.CI(n52759), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n52760));
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n52758), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_17_lut (.I0(GND_net), .I1(n16003[14]), .I2(GND_net), 
            .I3(n53825), .O(n14630[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_15_lut (.I0(GND_net), .I1(n14124[12]), .I2(n1029_adj_4719), 
            .I3(n53182), .O(n12531[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[23]), 
            .I3(n52903), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[22]), 
            .I3(n52902), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_17 (.CI(n53825), .I0(n16003[14]), .I1(GND_net), 
            .CO(n53826));
    SB_CARRY add_16_3 (.CI(n52758), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n52759));
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n52758));
    SB_CARRY add_4957_15 (.CI(n53182), .I0(n14124[12]), .I1(n1029_adj_4719), 
            .CO(n53183));
    SB_CARRY unary_minus_20_add_3_24 (.CI(n52902), .I0(GND_net), .I1(n1_adj_5021[22]), 
            .CO(n52903));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[21]), 
            .I3(n52901), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n52757), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n52756), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_16_lut (.I0(GND_net), .I1(n16003[13]), .I2(n1105), 
            .I3(n53824), .O(n14630[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_16 (.CI(n53824), .I0(n16003[13]), .I1(n1105), .CO(n53825));
    SB_LUT4 add_4957_14_lut (.I0(GND_net), .I1(n14124[11]), .I2(n956_adj_4723), 
            .I3(n53181), .O(n12531[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n52901), .I0(GND_net), .I1(n1_adj_5021[21]), 
            .CO(n52902));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[20]), 
            .I3(n52900), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_24 (.CI(n52756), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n52757));
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n52755), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51495_4_lut (.I0(\encoder1_position_scaled[0] ), .I1(n15), 
            .I2(n67541), .I3(n15_adj_1), .O(motor_state_c[0]));   // verilog/motorControl.v(53[17:33])
    defparam i51495_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 add_5045_15_lut (.I0(GND_net), .I1(n16003[12]), .I2(n1032), 
            .I3(n53823), .O(n14630[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_15 (.CI(n53823), .I0(n16003[12]), .I1(n1032), .CO(n53824));
    SB_CARRY add_4957_14 (.CI(n53181), .I0(n14124[11]), .I1(n956_adj_4723), 
            .CO(n53182));
    SB_CARRY unary_minus_20_add_3_22 (.CI(n52900), .I0(GND_net), .I1(n1_adj_5021[20]), 
            .CO(n52901));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[19]), 
            .I3(n52899), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_23 (.CI(n52755), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n52756));
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n52754), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_14_lut (.I0(GND_net), .I1(n16003[11]), .I2(n959), 
            .I3(n53822), .O(n14630[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_13_lut (.I0(GND_net), .I1(n14124[10]), .I2(n883_adj_4728), 
            .I3(n53180), .O(n12531[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_13 (.CI(n53180), .I0(n14124[10]), .I1(n883_adj_4728), 
            .CO(n53181));
    SB_CARRY add_5045_14 (.CI(n53822), .I0(n16003[11]), .I1(n959), .CO(n53823));
    SB_LUT4 add_4957_12_lut (.I0(GND_net), .I1(n14124[9]), .I2(n810_adj_4729), 
            .I3(n53179), .O(n12531[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_12 (.CI(n53179), .I0(n14124[9]), .I1(n810_adj_4729), 
            .CO(n53180));
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5045_13_lut (.I0(GND_net), .I1(n16003[10]), .I2(n886), 
            .I3(n53821), .O(n14630[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_11_lut (.I0(GND_net), .I1(n14124[8]), .I2(n737_adj_4730), 
            .I3(n53178), .O(n12531[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_11 (.CI(n53178), .I0(n14124[8]), .I1(n737_adj_4730), 
            .CO(n53179));
    SB_CARRY add_5045_13 (.CI(n53821), .I0(n16003[10]), .I1(n886), .CO(n53822));
    SB_LUT4 add_4957_10_lut (.I0(GND_net), .I1(n14124[7]), .I2(n664_adj_4731), 
            .I3(n53177), .O(n12531[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_10 (.CI(n53177), .I0(n14124[7]), .I1(n664_adj_4731), 
            .CO(n53178));
    SB_LUT4 add_5045_12_lut (.I0(GND_net), .I1(n16003[9]), .I2(n813), 
            .I3(n53820), .O(n14630[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_9_lut (.I0(GND_net), .I1(n14124[6]), .I2(n591_adj_4732), 
            .I3(n53176), .O(n12531[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_9 (.CI(n53176), .I0(n14124[6]), .I1(n591_adj_4732), 
            .CO(n53177));
    SB_CARRY add_5045_12 (.CI(n53820), .I0(n16003[9]), .I1(n813), .CO(n53821));
    SB_LUT4 add_4957_8_lut (.I0(GND_net), .I1(n14124[5]), .I2(n518_adj_4733), 
            .I3(n53175), .O(n12531[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_22 (.CI(n52754), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n52755));
    SB_CARRY unary_minus_20_add_3_21 (.CI(n52899), .I0(GND_net), .I1(n1_adj_5021[19]), 
            .CO(n52900));
    SB_LUT4 add_5045_11_lut (.I0(GND_net), .I1(n16003[8]), .I2(n740), 
            .I3(n53819), .O(n14630[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_8 (.CI(n53175), .I0(n14124[5]), .I1(n518_adj_4733), 
            .CO(n53176));
    SB_LUT4 add_4957_7_lut (.I0(GND_net), .I1(n14124[4]), .I2(n445_adj_4734), 
            .I3(n53174), .O(n12531[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_11 (.CI(n53819), .I0(n16003[8]), .I1(n740), .CO(n53820));
    SB_LUT4 add_5045_10_lut (.I0(GND_net), .I1(n16003[7]), .I2(n667), 
            .I3(n53818), .O(n14630[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_7 (.CI(n53174), .I0(n14124[4]), .I1(n445_adj_4734), 
            .CO(n53175));
    SB_CARRY add_5045_10 (.CI(n53818), .I0(n16003[7]), .I1(n667), .CO(n53819));
    SB_LUT4 add_5045_9_lut (.I0(GND_net), .I1(n16003[6]), .I2(n594), .I3(n53817), 
            .O(n14630[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4957_6_lut (.I0(GND_net), .I1(n14124[3]), .I2(n372_adj_4735), 
            .I3(n53173), .O(n12531[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[18]), 
            .I3(n52898), .O(n285[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_9 (.CI(n53817), .I0(n16003[6]), .I1(n594), .CO(n53818));
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n52753), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n52898), .I0(GND_net), .I1(n1_adj_5021[18]), 
            .CO(n52899));
    SB_LUT4 add_5045_8_lut (.I0(GND_net), .I1(n16003[5]), .I2(n521), .I3(n53816), 
            .O(n14630[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_8 (.CI(n53816), .I0(n16003[5]), .I1(n521), .CO(n53817));
    SB_CARRY add_4957_6 (.CI(n53173), .I0(n14124[3]), .I1(n372_adj_4735), 
            .CO(n53174));
    SB_LUT4 add_4957_5_lut (.I0(GND_net), .I1(n14124[2]), .I2(n299_adj_4737), 
            .I3(n53172), .O(n12531[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_7_lut (.I0(GND_net), .I1(n16003[4]), .I2(n448_adj_4738), 
            .I3(n53815), .O(n14630[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_5 (.CI(n53172), .I0(n14124[2]), .I1(n299_adj_4737), 
            .CO(n53173));
    SB_LUT4 add_4957_4_lut (.I0(GND_net), .I1(n14124[1]), .I2(n226_adj_4739), 
            .I3(n53171), .O(n12531[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_7 (.CI(n53815), .I0(n16003[4]), .I1(n448_adj_4738), 
            .CO(n53816));
    SB_CARRY add_4957_4 (.CI(n53171), .I0(n14124[1]), .I1(n226_adj_4739), 
            .CO(n53172));
    SB_LUT4 add_4957_3_lut (.I0(GND_net), .I1(n14124[0]), .I2(n153_adj_4740), 
            .I3(n53170), .O(n12531[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_6_lut (.I0(GND_net), .I1(n16003[3]), .I2(n375), .I3(n53814), 
            .O(n14630[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4957_3 (.CI(n53170), .I0(n14124[0]), .I1(n153_adj_4740), 
            .CO(n53171));
    SB_LUT4 add_4957_2_lut (.I0(GND_net), .I1(n11_adj_4741), .I2(n80_adj_4742), 
            .I3(GND_net), .O(n12531[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4957_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_6 (.CI(n53814), .I0(n16003[3]), .I1(n375), .CO(n53815));
    SB_CARRY add_4957_2 (.CI(GND_net), .I0(n11_adj_4741), .I1(n80_adj_4742), 
            .CO(n53170));
    SB_LUT4 add_5045_5_lut (.I0(GND_net), .I1(n16003[2]), .I2(n302), .I3(n53813), 
            .O(n14630[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_5 (.CI(n53813), .I0(n16003[2]), .I1(n302), .CO(n53814));
    SB_LUT4 add_5022_21_lut (.I0(GND_net), .I1(n15560[18]), .I2(GND_net), 
            .I3(n53169), .O(n14124[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[17]), 
            .I3(n52897), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_4_lut (.I0(GND_net), .I1(n16003[1]), .I2(n229), .I3(n53812), 
            .O(n14630[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_20_lut (.I0(GND_net), .I1(n15560[17]), .I2(GND_net), 
            .I3(n53168), .O(n14124[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_20 (.CI(n53168), .I0(n15560[17]), .I1(GND_net), 
            .CO(n53169));
    SB_CARRY unary_minus_20_add_3_19 (.CI(n52897), .I0(GND_net), .I1(n1_adj_5021[17]), 
            .CO(n52898));
    SB_CARRY add_5045_4 (.CI(n53812), .I0(n16003[1]), .I1(n229), .CO(n53813));
    SB_LUT4 add_5022_19_lut (.I0(GND_net), .I1(n15560[16]), .I2(GND_net), 
            .I3(n53167), .O(n14124[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_19 (.CI(n53167), .I0(n15560[16]), .I1(GND_net), 
            .CO(n53168));
    SB_LUT4 add_5045_3_lut (.I0(GND_net), .I1(n16003[0]), .I2(n156), .I3(n53811), 
            .O(n14630[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_18_lut (.I0(GND_net), .I1(n15560[15]), .I2(GND_net), 
            .I3(n53166), .O(n14124[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_18 (.CI(n53166), .I0(n15560[15]), .I1(GND_net), 
            .CO(n53167));
    SB_CARRY add_5045_3 (.CI(n53811), .I0(n16003[0]), .I1(n156), .CO(n53812));
    SB_LUT4 add_5022_17_lut (.I0(GND_net), .I1(n15560[14]), .I2(GND_net), 
            .I3(n53165), .O(n14124[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_17 (.CI(n53165), .I0(n15560[14]), .I1(GND_net), 
            .CO(n53166));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[16]), 
            .I3(n52896), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5045_2_lut (.I0(GND_net), .I1(n14_adj_4745), .I2(n83), 
            .I3(GND_net), .O(n14630[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_16_lut (.I0(GND_net), .I1(n15560[13]), .I2(n1105_adj_4746), 
            .I3(n53164), .O(n14124[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_16 (.CI(n53164), .I0(n15560[13]), .I1(n1105_adj_4746), 
            .CO(n53165));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n52896), .I0(GND_net), .I1(n1_adj_5021[16]), 
            .CO(n52897));
    SB_CARRY add_5045_2 (.CI(GND_net), .I0(n14_adj_4745), .I1(n83), .CO(n53811));
    SB_LUT4 add_5022_15_lut (.I0(GND_net), .I1(n15560[12]), .I2(n1032_adj_4747), 
            .I3(n53163), .O(n14124[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_15 (.CI(n53163), .I0(n15560[12]), .I1(n1032_adj_4747), 
            .CO(n53164));
    SB_LUT4 add_5104_20_lut (.I0(GND_net), .I1(n17230[17]), .I2(GND_net), 
            .I3(n53810), .O(n16003[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_14_lut (.I0(GND_net), .I1(n15560[11]), .I2(n959_adj_4748), 
            .I3(n53162), .O(n14124[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_14 (.CI(n53162), .I0(n15560[11]), .I1(n959_adj_4748), 
            .CO(n53163));
    SB_LUT4 add_5104_19_lut (.I0(GND_net), .I1(n17230[16]), .I2(GND_net), 
            .I3(n53809), .O(n16003[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_13_lut (.I0(GND_net), .I1(n15560[10]), .I2(n886_adj_4749), 
            .I3(n53161), .O(n14124[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_13 (.CI(n53161), .I0(n15560[10]), .I1(n886_adj_4749), 
            .CO(n53162));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[15]), 
            .I3(n52895), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_19 (.CI(n53809), .I0(n17230[16]), .I1(GND_net), 
            .CO(n53810));
    SB_LUT4 add_5104_18_lut (.I0(GND_net), .I1(n17230[15]), .I2(GND_net), 
            .I3(n53808), .O(n16003[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_12_lut (.I0(GND_net), .I1(n15560[9]), .I2(n813_adj_4751), 
            .I3(n53160), .O(n14124[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_12 (.CI(n53160), .I0(n15560[9]), .I1(n813_adj_4751), 
            .CO(n53161));
    SB_CARRY add_5104_18 (.CI(n53808), .I0(n17230[15]), .I1(GND_net), 
            .CO(n53809));
    SB_LUT4 add_5022_11_lut (.I0(GND_net), .I1(n15560[8]), .I2(n740_adj_4752), 
            .I3(n53159), .O(n14124[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_11 (.CI(n53159), .I0(n15560[8]), .I1(n740_adj_4752), 
            .CO(n53160));
    SB_LUT4 add_5104_17_lut (.I0(GND_net), .I1(n17230[14]), .I2(GND_net), 
            .I3(n53807), .O(n16003[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_10_lut (.I0(GND_net), .I1(n15560[7]), .I2(n667_adj_4753), 
            .I3(n53158), .O(n14124[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_10 (.CI(n53158), .I0(n15560[7]), .I1(n667_adj_4753), 
            .CO(n53159));
    SB_CARRY add_5104_17 (.CI(n53807), .I0(n17230[14]), .I1(GND_net), 
            .CO(n53808));
    SB_LUT4 add_5022_9_lut (.I0(GND_net), .I1(n15560[6]), .I2(n594_adj_4754), 
            .I3(n53157), .O(n14124[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_9 (.CI(n53157), .I0(n15560[6]), .I1(n594_adj_4754), 
            .CO(n53158));
    SB_LUT4 add_5104_16_lut (.I0(GND_net), .I1(n17230[13]), .I2(n1108), 
            .I3(n53806), .O(n16003[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_8_lut (.I0(GND_net), .I1(n15560[5]), .I2(n521_adj_4755), 
            .I3(n53156), .O(n14124[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_16 (.CI(n53806), .I0(n17230[13]), .I1(n1108), .CO(n53807));
    SB_CARRY add_5022_8 (.CI(n53156), .I0(n15560[5]), .I1(n521_adj_4755), 
            .CO(n53157));
    SB_LUT4 add_5104_15_lut (.I0(GND_net), .I1(n17230[12]), .I2(n1035), 
            .I3(n53805), .O(n16003[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_7_lut (.I0(GND_net), .I1(n15560[4]), .I2(n448_adj_4756), 
            .I3(n53155), .O(n14124[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_7 (.CI(n53155), .I0(n15560[4]), .I1(n448_adj_4756), 
            .CO(n53156));
    SB_CARRY add_5104_15 (.CI(n53805), .I0(n17230[12]), .I1(n1035), .CO(n53806));
    SB_LUT4 add_5022_6_lut (.I0(GND_net), .I1(n15560[3]), .I2(n375_adj_4757), 
            .I3(n53154), .O(n14124[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_6 (.CI(n53154), .I0(n15560[3]), .I1(n375_adj_4757), 
            .CO(n53155));
    SB_LUT4 add_5104_14_lut (.I0(GND_net), .I1(n17230[11]), .I2(n962), 
            .I3(n53804), .O(n16003[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_5_lut (.I0(GND_net), .I1(n15560[2]), .I2(n302_adj_4758), 
            .I3(n53153), .O(n14124[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_5 (.CI(n53153), .I0(n15560[2]), .I1(n302_adj_4758), 
            .CO(n53154));
    SB_CARRY add_5104_14 (.CI(n53804), .I0(n17230[11]), .I1(n962), .CO(n53805));
    SB_LUT4 add_5022_4_lut (.I0(GND_net), .I1(n15560[1]), .I2(n229_adj_4759), 
            .I3(n53152), .O(n14124[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_4 (.CI(n53152), .I0(n15560[1]), .I1(n229_adj_4759), 
            .CO(n53153));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n52895), .I0(GND_net), .I1(n1_adj_5021[15]), 
            .CO(n52896));
    SB_LUT4 add_5104_13_lut (.I0(GND_net), .I1(n17230[10]), .I2(n889), 
            .I3(n53803), .O(n16003[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_13 (.CI(n53803), .I0(n17230[10]), .I1(n889), .CO(n53804));
    SB_LUT4 add_5022_3_lut (.I0(GND_net), .I1(n15560[0]), .I2(n156_adj_4760), 
            .I3(n53151), .O(n14124[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_3 (.CI(n53151), .I0(n15560[0]), .I1(n156_adj_4760), 
            .CO(n53152));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[14]), 
            .I3(n52894), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5104_12_lut (.I0(GND_net), .I1(n17230[9]), .I2(n816), 
            .I3(n53802), .O(n16003[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_2_lut (.I0(GND_net), .I1(n14_adj_4762), .I2(n83_adj_4763), 
            .I3(GND_net), .O(n14124[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_2 (.CI(GND_net), .I0(n14_adj_4762), .I1(n83_adj_4763), 
            .CO(n53151));
    SB_CARRY add_5104_12 (.CI(n53802), .I0(n17230[9]), .I1(n816), .CO(n53803));
    SB_LUT4 add_5083_20_lut (.I0(GND_net), .I1(n16847[17]), .I2(GND_net), 
            .I3(n53150), .O(n15560[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_19_lut (.I0(GND_net), .I1(n16847[16]), .I2(GND_net), 
            .I3(n53149), .O(n15560[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5104_11_lut (.I0(GND_net), .I1(n17230[8]), .I2(n743), 
            .I3(n53801), .O(n16003[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_11 (.CI(n53801), .I0(n17230[8]), .I1(n743), .CO(n53802));
    SB_CARRY add_5083_19 (.CI(n53149), .I0(n16847[16]), .I1(GND_net), 
            .CO(n53150));
    SB_LUT4 add_5083_18_lut (.I0(GND_net), .I1(n16847[15]), .I2(GND_net), 
            .I3(n53148), .O(n15560[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n52894), .I0(GND_net), .I1(n1_adj_5021[14]), 
            .CO(n52895));
    SB_LUT4 add_5104_10_lut (.I0(GND_net), .I1(n17230[7]), .I2(n670), 
            .I3(n53800), .O(n16003[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_18 (.CI(n53148), .I0(n16847[15]), .I1(GND_net), 
            .CO(n53149));
    SB_LUT4 add_5083_17_lut (.I0(GND_net), .I1(n16847[14]), .I2(GND_net), 
            .I3(n53147), .O(n15560[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_10 (.CI(n53800), .I0(n17230[7]), .I1(n670), .CO(n53801));
    SB_CARRY add_5083_17 (.CI(n53147), .I0(n16847[14]), .I1(GND_net), 
            .CO(n53148));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[13]), 
            .I3(n52893), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n52893), .I0(GND_net), .I1(n1_adj_5021[13]), 
            .CO(n52894));
    SB_LUT4 add_5083_16_lut (.I0(GND_net), .I1(n16847[13]), .I2(n1108_adj_4766), 
            .I3(n53146), .O(n15560[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[12]), 
            .I3(n52892), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n52892), .I0(GND_net), .I1(n1_adj_5021[12]), 
            .CO(n52893));
    SB_LUT4 add_5104_9_lut (.I0(GND_net), .I1(n17230[6]), .I2(n597), .I3(n53799), 
            .O(n16003[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_16 (.CI(n53146), .I0(n16847[13]), .I1(n1108_adj_4766), 
            .CO(n53147));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[11]), 
            .I3(n52891), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_15_lut (.I0(GND_net), .I1(n16847[12]), .I2(n1035_adj_4769), 
            .I3(n53145), .O(n15560[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_9 (.CI(n53799), .I0(n17230[6]), .I1(n597), .CO(n53800));
    SB_LUT4 add_5104_8_lut (.I0(GND_net), .I1(n17230[5]), .I2(n524), .I3(n53798), 
            .O(n16003[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n52891), .I0(GND_net), .I1(n1_adj_5021[11]), 
            .CO(n52892));
    SB_CARRY add_5083_15 (.CI(n53145), .I0(n16847[12]), .I1(n1035_adj_4769), 
            .CO(n53146));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[10]), 
            .I3(n52890), .O(n285[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n52890), .I0(GND_net), .I1(n1_adj_5021[10]), 
            .CO(n52891));
    SB_CARRY add_5104_8 (.CI(n53798), .I0(n17230[5]), .I1(n524), .CO(n53799));
    SB_LUT4 add_5083_14_lut (.I0(GND_net), .I1(n16847[11]), .I2(n962_adj_4771), 
            .I3(n53144), .O(n15560[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[9]), 
            .I3(n52889), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n52889), .I0(GND_net), .I1(n1_adj_5021[9]), 
            .CO(n52890));
    SB_CARRY add_5083_14 (.CI(n53144), .I0(n16847[11]), .I1(n962_adj_4771), 
            .CO(n53145));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[8]), 
            .I3(n52888), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n52888), .I0(GND_net), .I1(n1_adj_5021[8]), 
            .CO(n52889));
    SB_CARRY sub_15_add_2_21 (.CI(n52753), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n52754));
    SB_LUT4 add_5104_7_lut (.I0(GND_net), .I1(n17230[4]), .I2(n451_adj_4774), 
            .I3(n53797), .O(n16003[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_13_lut (.I0(GND_net), .I1(n16847[10]), .I2(n889_adj_4775), 
            .I3(n53143), .O(n15560[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[7]), 
            .I3(n52887), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n52887), .I0(GND_net), .I1(n1_adj_5021[7]), 
            .CO(n52888));
    SB_CARRY add_5083_13 (.CI(n53143), .I0(n16847[10]), .I1(n889_adj_4775), 
            .CO(n53144));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[6]), 
            .I3(n52886), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n52886), .I0(GND_net), .I1(n1_adj_5021[6]), 
            .CO(n52887));
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n52752), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_7 (.CI(n53797), .I0(n17230[4]), .I1(n451_adj_4774), 
            .CO(n53798));
    SB_LUT4 add_5083_12_lut (.I0(GND_net), .I1(n16847[9]), .I2(n816_adj_4779), 
            .I3(n53142), .O(n15560[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[5]), 
            .I3(n52885), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n52885), .I0(GND_net), .I1(n1_adj_5021[5]), 
            .CO(n52886));
    SB_CARRY add_5083_12 (.CI(n53142), .I0(n16847[9]), .I1(n816_adj_4779), 
            .CO(n53143));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[4]), 
            .I3(n52884), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n52884), .I0(GND_net), .I1(n1_adj_5021[4]), 
            .CO(n52885));
    SB_LUT4 add_5104_6_lut (.I0(GND_net), .I1(n17230[3]), .I2(n378), .I3(n53796), 
            .O(n16003[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_11_lut (.I0(GND_net), .I1(n16847[8]), .I2(n743_adj_4782), 
            .I3(n53141), .O(n15560[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[3]), 
            .I3(n52883), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n52883), .I0(GND_net), .I1(n1_adj_5021[3]), 
            .CO(n52884));
    SB_CARRY add_5104_6 (.CI(n53796), .I0(n17230[3]), .I1(n378), .CO(n53797));
    SB_LUT4 add_5104_5_lut (.I0(GND_net), .I1(n17230[2]), .I2(n305_adj_4784), 
            .I3(n53795), .O(n16003[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_5 (.CI(n53795), .I0(n17230[2]), .I1(n305_adj_4784), 
            .CO(n53796));
    SB_LUT4 add_5104_4_lut (.I0(GND_net), .I1(n17230[1]), .I2(n232), .I3(n53794), 
            .O(n16003[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_11 (.CI(n53141), .I0(n16847[8]), .I1(n743_adj_4782), 
            .CO(n53142));
    SB_CARRY add_5104_4 (.CI(n53794), .I0(n17230[1]), .I1(n232), .CO(n53795));
    SB_LUT4 add_5083_10_lut (.I0(GND_net), .I1(n16847[7]), .I2(n670_adj_4785), 
            .I3(n53140), .O(n15560[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5104_3_lut (.I0(GND_net), .I1(n17230[0]), .I2(n159), .I3(n53793), 
            .O(n16003[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_3 (.CI(n53793), .I0(n17230[0]), .I1(n159), .CO(n53794));
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[2]), 
            .I3(n52882), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_10 (.CI(n53140), .I0(n16847[7]), .I1(n670_adj_4785), 
            .CO(n53141));
    SB_CARRY unary_minus_20_add_3_4 (.CI(n52882), .I0(GND_net), .I1(n1_adj_5021[2]), 
            .CO(n52883));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[1]), 
            .I3(n52881), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_9_lut (.I0(GND_net), .I1(n16847[6]), .I2(n597_adj_4789), 
            .I3(n53139), .O(n15560[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n52881), .I0(GND_net), .I1(n1_adj_5021[1]), 
            .CO(n52882));
    SB_LUT4 add_5104_2_lut (.I0(GND_net), .I1(n17_adj_4790), .I2(n86), 
            .I3(GND_net), .O(n16003[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5104_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5104_2 (.CI(GND_net), .I0(n17_adj_4790), .I1(n86), .CO(n53793));
    SB_CARRY add_5083_9 (.CI(n53139), .I0(n16847[6]), .I1(n597_adj_4789), 
            .CO(n53140));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5021[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5021[0]), 
            .CO(n52881));
    SB_LUT4 add_5083_8_lut (.I0(GND_net), .I1(n16847[5]), .I2(n524_adj_4792), 
            .I3(n53138), .O(n15560[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n52752), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n52753));
    SB_CARRY add_5083_8 (.CI(n53138), .I0(n16847[5]), .I1(n524_adj_4792), 
            .CO(n53139));
    SB_LUT4 add_5083_7_lut (.I0(GND_net), .I1(n16847[4]), .I2(n451_adj_4793), 
            .I3(n53137), .O(n15560[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n52751), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_7 (.CI(n53137), .I0(n16847[4]), .I1(n451_adj_4793), 
            .CO(n53138));
    SB_LUT4 add_5083_6_lut (.I0(GND_net), .I1(n16847[3]), .I2(n378_adj_4794), 
            .I3(n53136), .O(n15560[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_19 (.CI(n52751), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n52752));
    SB_CARRY add_5083_6 (.CI(n53136), .I0(n16847[3]), .I1(n378_adj_4794), 
            .CO(n53137));
    SB_LUT4 add_5083_5_lut (.I0(GND_net), .I1(n16847[2]), .I2(n305_adj_4795), 
            .I3(n53135), .O(n15560[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n52750), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n52750), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n52751));
    SB_CARRY add_5083_5 (.CI(n53135), .I0(n16847[2]), .I1(n305_adj_4795), 
            .CO(n53136));
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n52749), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n52749), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n52750));
    SB_LUT4 add_5083_4_lut (.I0(GND_net), .I1(n16847[1]), .I2(n232_adj_4796), 
            .I3(n53134), .O(n15560[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_4 (.CI(n53134), .I0(n16847[1]), .I1(n232_adj_4796), 
            .CO(n53135));
    SB_LUT4 add_5083_3_lut (.I0(GND_net), .I1(n16847[0]), .I2(n159_adj_4797), 
            .I3(n53133), .O(n15560[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n52748), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_16 (.CI(n52748), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n52749));
    SB_CARRY add_5083_3 (.CI(n53133), .I0(n16847[0]), .I1(n159_adj_4797), 
            .CO(n53134));
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n52747), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n52747), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n52748));
    SB_LUT4 add_5083_2_lut (.I0(GND_net), .I1(n17_adj_4798), .I2(n86_adj_4799), 
            .I3(GND_net), .O(n15560[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n52746), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n52746), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n52747));
    SB_CARRY add_5083_2 (.CI(GND_net), .I0(n17_adj_4798), .I1(n86_adj_4799), 
            .CO(n53133));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n52745), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n52745), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n52746));
    SB_LUT4 add_5140_19_lut (.I0(GND_net), .I1(n17992[16]), .I2(GND_net), 
            .I3(n53132), .O(n16847[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_18_lut (.I0(GND_net), .I1(n17992[15]), .I2(GND_net), 
            .I3(n53131), .O(n16847[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_18 (.CI(n53131), .I0(n17992[15]), .I1(GND_net), 
            .CO(n53132));
    SB_LUT4 add_5140_17_lut (.I0(GND_net), .I1(n17992[14]), .I2(GND_net), 
            .I3(n53130), .O(n16847[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4800));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5140_17 (.CI(n53130), .I0(n17992[14]), .I1(GND_net), 
            .CO(n53131));
    SB_LUT4 add_5140_16_lut (.I0(GND_net), .I1(n17992[13]), .I2(n1111_adj_4801), 
            .I3(n53129), .O(n16847[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_16 (.CI(n53129), .I0(n17992[13]), .I1(n1111_adj_4801), 
            .CO(n53130));
    SB_LUT4 add_5140_15_lut (.I0(GND_net), .I1(n17992[12]), .I2(n1038_adj_4802), 
            .I3(n53128), .O(n16847[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_15 (.CI(n53128), .I0(n17992[12]), .I1(n1038_adj_4802), 
            .CO(n53129));
    SB_LUT4 add_5140_14_lut (.I0(GND_net), .I1(n17992[11]), .I2(n965_adj_4803), 
            .I3(n53127), .O(n16847[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_14 (.CI(n53127), .I0(n17992[11]), .I1(n965_adj_4803), 
            .CO(n53128));
    SB_LUT4 add_5140_13_lut (.I0(GND_net), .I1(n17992[10]), .I2(n892_adj_4804), 
            .I3(n53126), .O(n16847[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_13 (.CI(n53126), .I0(n17992[10]), .I1(n892_adj_4804), 
            .CO(n53127));
    SB_LUT4 add_5140_12_lut (.I0(GND_net), .I1(n17992[9]), .I2(n819_adj_4805), 
            .I3(n53125), .O(n16847[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_12 (.CI(n53125), .I0(n17992[9]), .I1(n819_adj_4805), 
            .CO(n53126));
    SB_LUT4 add_5140_11_lut (.I0(GND_net), .I1(n17992[8]), .I2(n746_adj_4806), 
            .I3(n53124), .O(n16847[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n335[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4453));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4452));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44827_2_lut (.I0(counter[13]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n64310));
    defparam i44827_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(counter[5]), .I1(counter[4]), .I2(counter[3]), 
            .I3(counter[8]), .O(n23_adj_4807));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5140_11 (.CI(n53124), .I0(n17992[8]), .I1(n746_adj_4806), 
            .CO(n53125));
    SB_LUT4 add_5159_19_lut (.I0(GND_net), .I1(n18318[16]), .I2(GND_net), 
            .I3(n53772), .O(n17230[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_18_lut (.I0(GND_net), .I1(n18318[15]), .I2(GND_net), 
            .I3(n53771), .O(n17230[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_18 (.CI(n53771), .I0(n18318[15]), .I1(GND_net), 
            .CO(n53772));
    SB_LUT4 i8_4_lut (.I0(counter[1]), .I1(counter[6]), .I2(counter[10]), 
            .I3(counter[0]), .O(n22_adj_4808));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i12_4_lut (.I0(n23_adj_4807), .I1(counter[2]), .I2(n64310), 
            .I3(counter[9]), .O(n26_adj_4809));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 add_5159_17_lut (.I0(GND_net), .I1(n18318[14]), .I2(GND_net), 
            .I3(n53770), .O(n17230[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51514_4_lut (.I0(counter[12]), .I1(n26_adj_4809), .I2(n22_adj_4808), 
            .I3(counter[7]), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i51514_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 add_5140_10_lut (.I0(GND_net), .I1(n17992[7]), .I2(n673), 
            .I3(n53123), .O(n16847[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5159_17 (.CI(n53770), .I0(n18318[14]), .I1(GND_net), 
            .CO(n53771));
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4451));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4450));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4529));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71487_bdd_4_lut (.I0(n71487), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4749), .O(n71490));
    defparam n71487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n233[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51939 (.I0(n9977), .I1(n67727), .I2(setpoint[13]), 
            .I3(n4749), .O(n71481));
    defparam n9977_bdd_4_lut_51939.LUT_INIT = 16'he4aa;
    SB_LUT4 i49015_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9_adj_4810), 
            .O(n68510));
    defparam i49015_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48994_4_lut (.I0(n27), .I1(n15_adj_4811), .I2(n13_adj_4812), 
            .I3(n11_adj_4813), .O(n68489));
    defparam i48994_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4814));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4528));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4810));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4813));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4812));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4811));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4815));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4816));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4817));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n335[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4477));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4818));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4476));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4475));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4526));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4472));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4469));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5159_16_lut (.I0(GND_net), .I1(n18318[13]), .I2(n1111), 
            .I3(n53769), .O(n17230[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4464));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4806));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4805));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4804));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4803));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4802));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4801));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4799));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4798));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4462));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4797));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4796));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4795));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4794));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4793));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4461));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4460));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4792));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4790));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4789));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4459));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4458));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4785));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4784));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4782));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4457));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4456));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4779));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4775));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4774));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4771));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4769));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4766));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4763));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4762));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4760));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4759));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4758));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4757));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4756));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4755));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4754));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4753));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4752));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4751));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4748));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4747));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4746));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4745));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4742));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4741));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4739));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4738));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4735));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4734));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4733));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4732));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4730));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4729));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4728));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4723));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5021[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4719));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23108_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41203));   // verilog/motorControl.v(61[20:40])
    defparam i23108_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4715));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4704));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4698));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4696));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4694));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4689));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4685));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4684));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4681));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4525));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_4812), 
            .I3(GND_net), .O(n10_adj_4819));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_4814), .I1(n233[17]), .I2(n35_adj_4800), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5020[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4672));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4523));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4668));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50019_4_lut (.I0(n13_adj_4812), .I1(n11_adj_4813), .I2(n9_adj_4810), 
            .I3(n68528), .O(n69514));
    defparam i50019_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4820));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4821));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4822));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4522));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4662));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4659));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4823));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50013_4_lut (.I0(n19), .I1(n17), .I2(n15_adj_4811), .I3(n69514), 
            .O(n69508));
    defparam i50013_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4824));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4825));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4826));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4827));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4828));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4829));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4830));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4831));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4832));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4833));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4834));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4835));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4836));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4837));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4838));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49093_4_lut (.I0(n21_adj_4838), .I1(n19_adj_4837), .I2(n17_adj_4836), 
            .I3(n9_adj_4835), .O(n68588));
    defparam i49093_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49081_4_lut (.I0(n27_adj_4834), .I1(n15_adj_4833), .I2(n13_adj_4832), 
            .I3(n11_adj_4831), .O(n68576));
    defparam i49081_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4830), 
            .I3(GND_net), .O(n12_adj_4839));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4832), 
            .I3(GND_net), .O(n10_adj_4840));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4839), .I1(n535[17]), .I2(n35_adj_4829), 
            .I3(GND_net), .O(n30_adj_4841));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50085_4_lut (.I0(n13_adj_4832), .I1(n11_adj_4831), .I2(n9_adj_4835), 
            .I3(n68608), .O(n69580));
    defparam i50085_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50077_4_lut (.I0(n19_adj_4837), .I1(n17_adj_4836), .I2(n15_adj_4833), 
            .I3(n69580), .O(n69572));
    defparam i50077_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51109_4_lut (.I0(n25_adj_4828), .I1(n23_adj_4827), .I2(n21_adj_4838), 
            .I3(n69572), .O(n70604));
    defparam i51109_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50537_4_lut (.I0(n31_adj_4825), .I1(n29_adj_4824), .I2(n27_adj_4834), 
            .I3(n70604), .O(n70032));
    defparam i50537_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51242_4_lut (.I0(n37_adj_4826), .I1(n35_adj_4829), .I2(n33_adj_4830), 
            .I3(n70032), .O(n70737));
    defparam i51242_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4823), 
            .I3(GND_net), .O(n16_adj_4842));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50799_3_lut (.I0(n6_adj_4843), .I1(n535[10]), .I2(n21_adj_4838), 
            .I3(GND_net), .O(n70294));   // verilog/motorControl.v(47[25:43])
    defparam i50799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50800_3_lut (.I0(n70294), .I1(n535[11]), .I2(n23_adj_4827), 
            .I3(GND_net), .O(n70295));   // verilog/motorControl.v(47[25:43])
    defparam i50800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51101_4_lut (.I0(n25), .I1(n23_adj_4609), .I2(n21), .I3(n69508), 
            .O(n70596));
    defparam i51101_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4836), 
            .I3(GND_net), .O(n8_adj_4844));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4842), .I1(n535[22]), .I2(n45_adj_4822), 
            .I3(GND_net), .O(n24_adj_4845));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49042_4_lut (.I0(n43_adj_4823), .I1(n25_adj_4828), .I2(n23_adj_4827), 
            .I3(n68588), .O(n68537));
    defparam i49042_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50299_4_lut (.I0(n24_adj_4845), .I1(n8_adj_4844), .I2(n45_adj_4822), 
            .I3(n68530), .O(n69794));   // verilog/motorControl.v(47[25:43])
    defparam i50299_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50505_4_lut (.I0(n31), .I1(n29_adj_4636), .I2(n27), .I3(n70596), 
            .O(n70000));
    defparam i50505_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49504_3_lut (.I0(n70295), .I1(n535[12]), .I2(n25_adj_4828), 
            .I3(GND_net), .O(n68999));   // verilog/motorControl.v(47[25:43])
    defparam i49504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4846));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50795_3_lut (.I0(n4_adj_4846), .I1(n535[13]), .I2(n27_adj_4834), 
            .I3(GND_net), .O(n70290));   // verilog/motorControl.v(47[25:43])
    defparam i50795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50796_3_lut (.I0(n70290), .I1(n535[14]), .I2(n29_adj_4824), 
            .I3(GND_net), .O(n70291));   // verilog/motorControl.v(47[25:43])
    defparam i50796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49058_4_lut (.I0(n33_adj_4830), .I1(n31_adj_4825), .I2(n29_adj_4824), 
            .I3(n68576), .O(n68553));
    defparam i49058_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51115_4_lut (.I0(n30_adj_4841), .I1(n10_adj_4840), .I2(n35_adj_4829), 
            .I3(n68551), .O(n70610));   // verilog/motorControl.v(47[25:43])
    defparam i51115_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 n71481_bdd_4_lut (.I0(n71481), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4749), .O(n71484));
    defparam n71481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49506_3_lut (.I0(n70291), .I1(n535[15]), .I2(n31_adj_4825), 
            .I3(GND_net), .O(n69001));   // verilog/motorControl.v(47[25:43])
    defparam i49506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51323_4_lut (.I0(n69001), .I1(n70610), .I2(n35_adj_4829), 
            .I3(n68553), .O(n70818));   // verilog/motorControl.v(47[25:43])
    defparam i51323_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48874_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n68369));
    defparam i48874_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51324_3_lut (.I0(n70818), .I1(n535[18]), .I2(n37_adj_4826), 
            .I3(GND_net), .O(n70819));   // verilog/motorControl.v(47[25:43])
    defparam i51324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51310_3_lut (.I0(n70819), .I1(n535[19]), .I2(n39_adj_4821), 
            .I3(GND_net), .O(n70805));   // verilog/motorControl.v(47[25:43])
    defparam i51310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49044_4_lut (.I0(n43_adj_4823), .I1(n41_adj_4820), .I2(n39_adj_4821), 
            .I3(n70737), .O(n68539));
    defparam i49044_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50951_4_lut (.I0(n68999), .I1(n69794), .I2(n45_adj_4822), 
            .I3(n68537), .O(n70446));   // verilog/motorControl.v(47[25:43])
    defparam i50951_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49512_3_lut (.I0(n70805), .I1(n535[20]), .I2(n41_adj_4820), 
            .I3(GND_net), .O(n69007));   // verilog/motorControl.v(47[25:43])
    defparam i49512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51193_4_lut (.I0(n69007), .I1(n70446), .I2(n45_adj_4822), 
            .I3(n68539), .O(n70688));   // verilog/motorControl.v(47[25:43])
    defparam i51193_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48892_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n68387));
    defparam i48892_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51194_3_lut (.I0(n70688), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(GND_net), .O(n131_adj_4847));   // verilog/motorControl.v(47[25:43])
    defparam i51194_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4848));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n455[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4849));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4850));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4851));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4852));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4853));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n455[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4854));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4855));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4856));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n455[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4857));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4858));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n335[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4859));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4860));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4861));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n335[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n335[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4863));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4864));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4865));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4866));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4867));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i39_2_lut (.I0(deadband[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4868));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4869));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i45_2_lut (.I0(deadband[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4870));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(deadband[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4871));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(deadband[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4872));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48383_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n67878));
    defparam i48383_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i43_2_lut (.I0(deadband[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4873));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i37_2_lut (.I0(deadband[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4874));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4875));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4520));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(deadband[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4876));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(deadband[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4877));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i33_2_lut (.I0(deadband[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4878));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(deadband[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4879));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4880));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48447_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n67942));
    defparam i48447_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4881));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4882));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(deadband[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4883));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4884));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4885));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(deadband[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4886));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i41_2_lut (.I0(n455[20]), .I1(n34[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4887));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i39_2_lut (.I0(n455[19]), .I1(n34[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4888));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i45_2_lut (.I0(n455[22]), .I1(n34[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4889));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i37_2_lut (.I0(n455[18]), .I1(n34[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4890));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i43_2_lut (.I0(n455[21]), .I1(n34[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4891));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51234_4_lut (.I0(n37), .I1(n35_adj_4800), .I2(n33), .I3(n70000), 
            .O(n70729));
    defparam i51234_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_28_i23_2_lut (.I0(n455[11]), .I1(n34[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4892));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i25_2_lut (.I0(n455[12]), .I1(n34[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4893));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i29_2_lut (.I0(n455[14]), .I1(n34[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4894));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51934 (.I0(n9977), .I1(n67726), .I2(setpoint[12]), 
            .I3(n4749), .O(n71475));
    defparam n9977_bdd_4_lut_51934.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_28_i31_2_lut (.I0(n455[15]), .I1(n34[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4895));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i35_2_lut (.I0(n455[17]), .I1(n34[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4896));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i33_2_lut (.I0(n455[16]), .I1(n34[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4897));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i9_2_lut (.I0(n455[4]), .I1(n34[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4898));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i17_2_lut (.I0(n455[8]), .I1(n34[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4899));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i19_2_lut (.I0(n455[9]), .I1(n34[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4900));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i21_2_lut (.I0(n455[10]), .I1(n34[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4901));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i11_2_lut (.I0(n455[5]), .I1(n34[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4902));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i13_2_lut (.I0(n455[6]), .I1(n34[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4903));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i15_2_lut (.I0(n455[7]), .I1(n34[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4904));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i27_2_lut (.I0(n455[13]), .I1(n34[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4905));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48761_4_lut (.I0(n21_adj_4901), .I1(n19_adj_4900), .I2(n17_adj_4899), 
            .I3(n9_adj_4898), .O(n68256));
    defparam i48761_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48740_4_lut (.I0(n27_adj_4905), .I1(n15_adj_4904), .I2(n13_adj_4903), 
            .I3(n11_adj_4902), .O(n68235));
    defparam i48740_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n34[7]), .I1(n34[16]), .I2(n33_adj_4897), 
            .I3(GND_net), .O(n12_adj_4906));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n34[5]), .I1(n34[6]), .I2(n13_adj_4903), 
            .I3(GND_net), .O(n10_adj_4907));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_4906), .I1(n34[17]), .I2(n35_adj_4896), 
            .I3(GND_net), .O(n30_adj_4908));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49791_4_lut (.I0(n13_adj_4903), .I1(n11_adj_4902), .I2(n9_adj_4898), 
            .I3(n68277), .O(n69286));
    defparam i49791_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 n71475_bdd_4_lut (.I0(n71475), .I1(n535[12]), .I2(n455[12]), 
            .I3(n4749), .O(n71478));
    defparam n71475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49783_4_lut (.I0(n19_adj_4900), .I1(n17_adj_4899), .I2(n15_adj_4904), 
            .I3(n69286), .O(n69278));
    defparam i49783_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_9_i8_3_lut_3_lut (.I0(setpoint[4]), .I1(setpoint[8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_4909));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51051_4_lut (.I0(n25_adj_4893), .I1(n23_adj_4892), .I2(n21_adj_4901), 
            .I3(n69278), .O(n70546));
    defparam i51051_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49115_2_lut_4_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), .I2(PWMLimit[9]), 
            .I3(setpoint[9]), .O(n68610));
    defparam i49115_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50389_4_lut (.I0(n31_adj_4895), .I1(n29_adj_4894), .I2(n27_adj_4905), 
            .I3(n70546), .O(n69884));
    defparam i50389_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51216_4_lut (.I0(n37_adj_4890), .I1(n35_adj_4896), .I2(n33_adj_4897), 
            .I3(n69884), .O(n70711));
    defparam i51216_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n34[9]), .I1(n34[21]), .I2(n43_adj_4891), 
            .I3(GND_net), .O(n16_adj_4910));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50767_3_lut (.I0(n6_adj_4911), .I1(n34[10]), .I2(n21_adj_4901), 
            .I3(GND_net), .O(n70262));   // verilog/motorControl.v(62[35:55])
    defparam i50767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4657));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4656));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50768_3_lut (.I0(n70262), .I1(n34[11]), .I2(n23_adj_4892), 
            .I3(GND_net), .O(n70263));   // verilog/motorControl.v(62[35:55])
    defparam i50768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n34[4]), .I1(n34[8]), .I2(n17_adj_4899), 
            .I3(GND_net), .O(n8_adj_4912));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i24_3_lut (.I0(n16_adj_4910), .I1(n34[22]), .I2(n45_adj_4889), 
            .I3(GND_net), .O(n24_adj_4913));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48659_4_lut (.I0(n43_adj_4891), .I1(n25_adj_4893), .I2(n23_adj_4892), 
            .I3(n68256), .O(n68154));
    defparam i48659_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50307_4_lut (.I0(n24_adj_4913), .I1(n8_adj_4912), .I2(n45_adj_4889), 
            .I3(n68148), .O(n69802));   // verilog/motorControl.v(62[35:55])
    defparam i50307_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43_c), 
            .I3(GND_net), .O(n16_adj_4914));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49544_3_lut (.I0(n70263), .I1(n34[12]), .I2(n25_adj_4893), 
            .I3(GND_net), .O(n69039));   // verilog/motorControl.v(62[35:55])
    defparam i49544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n67585), .I1(n34[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_4915));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_9_i16_3_lut_3_lut (.I0(setpoint[9]), .I1(setpoint[21]), 
            .I2(PWMLimit[21]), .I3(GND_net), .O(n16_adj_4916));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50385_3_lut (.I0(n4_adj_4915), .I1(n34[13]), .I2(n27_adj_4905), 
            .I3(GND_net), .O(n69880));   // verilog/motorControl.v(62[35:55])
    defparam i50385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50386_3_lut (.I0(n69880), .I1(n34[14]), .I2(n29_adj_4894), 
            .I3(GND_net), .O(n69881));   // verilog/motorControl.v(62[35:55])
    defparam i50386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48730_4_lut (.I0(n33_adj_4897), .I1(n31_adj_4895), .I2(n29_adj_4894), 
            .I3(n68235), .O(n68225));
    defparam i48730_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9977_bdd_4_lut_51929 (.I0(n9977), .I1(n67725), .I2(setpoint[11]), 
            .I3(n4749), .O(n71469));
    defparam n9977_bdd_4_lut_51929.LUT_INIT = 16'he4aa;
    SB_LUT4 i51043_4_lut (.I0(n30_adj_4908), .I1(n10_adj_4907), .I2(n35_adj_4896), 
            .I3(n68220), .O(n70538));   // verilog/motorControl.v(62[35:55])
    defparam i51043_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49546_3_lut (.I0(n69881), .I1(n34[15]), .I2(n31_adj_4895), 
            .I3(GND_net), .O(n69041));   // verilog/motorControl.v(62[35:55])
    defparam i49546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51291_4_lut (.I0(n69041), .I1(n70538), .I2(n35_adj_4896), 
            .I3(n68225), .O(n70786));   // verilog/motorControl.v(62[35:55])
    defparam i51291_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51292_3_lut (.I0(n70786), .I1(n34[18]), .I2(n37_adj_4890), 
            .I3(GND_net), .O(n70787));   // verilog/motorControl.v(62[35:55])
    defparam i51292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51219_3_lut (.I0(n70787), .I1(n34[19]), .I2(n39_adj_4888), 
            .I3(GND_net), .O(n70714));   // verilog/motorControl.v(62[35:55])
    defparam i51219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i10_3_lut_3_lut (.I0(setpoint[5]), .I1(setpoint[6]), 
            .I2(PWMLimit[6]), .I3(GND_net), .O(n10_adj_4917));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48663_4_lut (.I0(n43_adj_4891), .I1(n41_adj_4887), .I2(n39_adj_4888), 
            .I3(n70711), .O(n68158));
    defparam i48663_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49168_2_lut_4_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), .I2(PWMLimit[7]), 
            .I3(setpoint[7]), .O(n68663));
    defparam i49168_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50959_4_lut (.I0(n69039), .I1(n69802), .I2(n45_adj_4889), 
            .I3(n68154), .O(n70454));   // verilog/motorControl.v(62[35:55])
    defparam i50959_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n71469_bdd_4_lut (.I0(n71469), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4749), .O(n71472));
    defparam n71469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49552_3_lut (.I0(n70714), .I1(n34[20]), .I2(n41_adj_4887), 
            .I3(GND_net), .O(n69047));   // verilog/motorControl.v(62[35:55])
    defparam i49552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51201_4_lut (.I0(n69047), .I1(n70454), .I2(n45_adj_4889), 
            .I3(n68158), .O(n70696));   // verilog/motorControl.v(62[35:55])
    defparam i51201_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51202_3_lut (.I0(n70696), .I1(n455[23]), .I2(n47_adj_4673), 
            .I3(GND_net), .O(n506));   // verilog/motorControl.v(62[35:55])
    defparam i51202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34367_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n23381[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34367_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i34369_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n52398));   // verilog/motorControl.v(61[29:40])
    defparam i34369_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_9_i12_3_lut_3_lut (.I0(setpoint[7]), .I1(setpoint[16]), 
            .I2(PWMLimit[16]), .I3(GND_net), .O(n12_adj_4918));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48848_4_lut (.I0(n21_adj_4882), .I1(n19_adj_4881), .I2(n17_adj_4880), 
            .I3(n9_adj_4879), .O(n68343));
    defparam i48848_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48834_4_lut (.I0(n27_adj_4886), .I1(n15_adj_4885), .I2(n13_adj_4884), 
            .I3(n11_adj_4883), .O(n68329));
    defparam i48834_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4878), 
            .I3(GND_net), .O(n12_adj_4919));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4884), 
            .I3(GND_net), .O(n10_adj_4920));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i30_3_lut (.I0(n12_adj_4919), .I1(n455[17]), .I2(n35_adj_4877), 
            .I3(GND_net), .O(n30_adj_4921));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48946_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n68441));
    defparam i48946_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i49871_4_lut (.I0(n13_adj_4884), .I1(n11_adj_4883), .I2(n9_adj_4879), 
            .I3(n68365), .O(n69366));
    defparam i49871_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i49861_4_lut (.I0(n19_adj_4881), .I1(n17_adj_4880), .I2(n15_adj_4885), 
            .I3(n69366), .O(n69356));
    defparam i49861_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51075_4_lut (.I0(n25_adj_4876), .I1(n23_adj_4875), .I2(n21_adj_4882), 
            .I3(n69356), .O(n70570));
    defparam i51075_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34396_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n23360[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34396_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i34398_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n52428));   // verilog/motorControl.v(61[29:40])
    defparam i34398_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i50437_4_lut (.I0(n31_adj_4872), .I1(n29_adj_4871), .I2(n27_adj_4886), 
            .I3(n70570), .O(n69932));
    defparam i50437_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51224_4_lut (.I0(n37_adj_4874), .I1(n35_adj_4877), .I2(n33_adj_4878), 
            .I3(n69932), .O(n70719));
    defparam i51224_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4873), 
            .I3(GND_net), .O(n16_adj_4922));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50773_3_lut (.I0(n6_adj_4923), .I1(n455[10]), .I2(n21_adj_4882), 
            .I3(GND_net), .O(n70268));   // verilog/motorControl.v(62[14:31])
    defparam i50773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50774_3_lut (.I0(n70268), .I1(n455[11]), .I2(n23_adj_4875), 
            .I3(GND_net), .O(n70269));   // verilog/motorControl.v(62[14:31])
    defparam i50774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4880), 
            .I3(GND_net), .O(n8_adj_4924));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i24_3_lut (.I0(n16_adj_4922), .I1(n455[22]), .I2(n45_adj_4870), 
            .I3(GND_net), .O(n24_adj_4925));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48789_4_lut (.I0(n43_adj_4873), .I1(n25_adj_4876), .I2(n23_adj_4875), 
            .I3(n68343), .O(n68284));
    defparam i48789_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50305_4_lut (.I0(n24_adj_4925), .I1(n8_adj_4924), .I2(n45_adj_4870), 
            .I3(n68279), .O(n69800));   // verilog/motorControl.v(62[14:31])
    defparam i50305_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49534_3_lut (.I0(n70269), .I1(n455[12]), .I2(n25_adj_4876), 
            .I3(GND_net), .O(n69029));   // verilog/motorControl.v(62[14:31])
    defparam i49534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_4926));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50771_3_lut (.I0(n4_adj_4926), .I1(n455[13]), .I2(n27_adj_4886), 
            .I3(GND_net), .O(n70266));   // verilog/motorControl.v(62[14:31])
    defparam i50771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48516_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(PWMLimit[9]), 
            .I3(n455[9]), .O(n68011));
    defparam i48516_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50772_3_lut (.I0(n70266), .I1(n455[14]), .I2(n29_adj_4871), 
            .I3(GND_net), .O(n70267));   // verilog/motorControl.v(62[14:31])
    defparam i50772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48825_4_lut (.I0(n33_adj_4878), .I1(n31_adj_4872), .I2(n29_adj_4871), 
            .I3(n68329), .O(n68320));
    defparam i48825_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51121_4_lut (.I0(n30_adj_4921), .I1(n10_adj_4920), .I2(n35_adj_4877), 
            .I3(n68314), .O(n70616));   // verilog/motorControl.v(62[14:31])
    defparam i51121_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49536_3_lut (.I0(n70267), .I1(n455[15]), .I2(n31_adj_4872), 
            .I3(GND_net), .O(n69031));   // verilog/motorControl.v(62[14:31])
    defparam i49536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51331_4_lut (.I0(n69031), .I1(n70616), .I2(n35_adj_4877), 
            .I3(n68320), .O(n70826));   // verilog/motorControl.v(62[14:31])
    defparam i51331_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51332_3_lut (.I0(n70826), .I1(n455[18]), .I2(n37_adj_4874), 
            .I3(GND_net), .O(n70827));   // verilog/motorControl.v(62[14:31])
    defparam i51332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48545_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(PWMLimit[7]), 
            .I3(n455[7]), .O(n68040));
    defparam i48545_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51302_3_lut (.I0(n70827), .I1(n455[19]), .I2(n39_adj_4868), 
            .I3(GND_net), .O(n70797));   // verilog/motorControl.v(62[14:31])
    defparam i51302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48797_4_lut (.I0(n43_adj_4873), .I1(n41_adj_4869), .I2(n39_adj_4868), 
            .I3(n70719), .O(n68292));
    defparam i48797_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50957_4_lut (.I0(n69029), .I1(n69800), .I2(n45_adj_4870), 
            .I3(n68284), .O(n70452));   // verilog/motorControl.v(62[14:31])
    defparam i50957_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49542_3_lut (.I0(n70797), .I1(n455[20]), .I2(n41_adj_4869), 
            .I3(GND_net), .O(n69037));   // verilog/motorControl.v(62[14:31])
    defparam i49542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51199_4_lut (.I0(n69037), .I1(n70452), .I2(n45_adj_4870), 
            .I3(n68292), .O(n70694));   // verilog/motorControl.v(62[14:31])
    defparam i51199_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51200_3_lut (.I0(n70694), .I1(deadband[23]), .I2(n455[23]), 
            .I3(GND_net), .O(n480));   // verilog/motorControl.v(62[14:31])
    defparam i51200_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4927));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4928));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i45_2_lut (.I0(PWMLimit[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4929));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4930));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4931));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i43_2_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4932));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4933));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48940_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n68435));   // verilog/motorControl.v(58[23:46])
    defparam i48940_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4934));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4519));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i23_2_lut (.I0(PWMLimit[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4935));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i25_2_lut (.I0(PWMLimit[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4936));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4937));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48784_2_lut_4_lut (.I0(deadband[21]), .I1(n455[21]), .I2(deadband[9]), 
            .I3(n455[9]), .O(n68279));
    defparam i48784_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4938));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4939));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4940));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n28[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4941));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50791_3_lut (.I0(n6), .I1(n233[10]), .I2(n21), .I3(GND_net), 
            .O(n70286));   // verilog/motorControl.v(56[14:36])
    defparam i50791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4942));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34539_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4943), 
            .I3(n23323[1]), .O(n6_adj_4483));   // verilog/motorControl.v(61[29:40])
    defparam i34539_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_30_i9_2_lut (.I0(PWMLimit[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4944));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4945));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4946));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5019[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i21_2_lut (.I0(PWMLimit[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4947));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23101_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41195));   // verilog/motorControl.v(42[14] 73[8])
    defparam i23101_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4644));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n335[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48615_4_lut (.I0(n21_adj_4947), .I1(n19_adj_4946), .I2(n17_adj_4945), 
            .I3(n9_adj_4944), .O(n68110));
    defparam i48615_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48593_4_lut (.I0(n27_adj_4942), .I1(n15_adj_4941), .I2(n13_adj_4940), 
            .I3(n11_adj_4939), .O(n68088));
    defparam i48593_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4643));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4642));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4938), 
            .I3(GND_net), .O(n12_adj_4949));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n335[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4517));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4940), 
            .I3(GND_net), .O(n10_adj_4950));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4641));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4640));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n12_adj_4949), .I1(n455[17]), .I2(n35_adj_4937), 
            .I3(GND_net), .O(n30_adj_4951));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4639));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4516));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49613_4_lut (.I0(n13_adj_4940), .I1(n11_adj_4939), .I2(n9_adj_4944), 
            .I3(n68146), .O(n69108));
    defparam i49613_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4638));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4637));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4634));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49607_4_lut (.I0(n19_adj_4946), .I1(n17_adj_4945), .I2(n15_adj_4941), 
            .I3(n69108), .O(n69102));
    defparam i49607_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4633));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50995_4_lut (.I0(n25_adj_4936), .I1(n23_adj_4935), .I2(n21_adj_4947), 
            .I3(n69102), .O(n70490));
    defparam i50995_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4632));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4631));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4630));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4629));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50327_4_lut (.I0(n31_adj_4931), .I1(n29_adj_4930), .I2(n27_adj_4942), 
            .I3(n70490), .O(n69822));
    defparam i50327_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51207_4_lut (.I0(n37_adj_4933), .I1(n35_adj_4937), .I2(n33_adj_4938), 
            .I3(n69822), .O(n70702));
    defparam i51207_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4932), 
            .I3(GND_net), .O(n16_adj_4952));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4626));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4625));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n335[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4623));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4622));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50377_3_lut (.I0(n6_adj_4953), .I1(n455[10]), .I2(n21_adj_4947), 
            .I3(GND_net), .O(n69872));   // verilog/motorControl.v(63[16:31])
    defparam i50377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4620));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4619));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50378_3_lut (.I0(n69872), .I1(n455[11]), .I2(n23_adj_4935), 
            .I3(GND_net), .O(n69873));   // verilog/motorControl.v(63[16:31])
    defparam i50378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4617));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4943), 
            .I3(n23323[1]), .O(n23266[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4945), 
            .I3(GND_net), .O(n8_adj_4954));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9977_bdd_4_lut_51924 (.I0(n9977), .I1(n67724), .I2(setpoint[10]), 
            .I3(n4749), .O(n71463));
    defparam n9977_bdd_4_lut_51924.LUT_INIT = 16'he4aa;
    SB_LUT4 n71463_bdd_4_lut (.I0(n71463), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4749), .O(n71466));
    defparam n71463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4616));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i24_3_lut (.I0(n16_adj_4952), .I1(n455[22]), .I2(n45_adj_4929), 
            .I3(GND_net), .O(n24_adj_4955));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4614));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4613));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48518_4_lut (.I0(n43_adj_4932), .I1(n25_adj_4936), .I2(n23_adj_4935), 
            .I3(n68110), .O(n68013));
    defparam i48518_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50309_4_lut (.I0(n24_adj_4955), .I1(n8_adj_4954), .I2(n45_adj_4929), 
            .I3(n68011), .O(n69804));   // verilog/motorControl.v(63[16:31])
    defparam i50309_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48819_2_lut_4_lut (.I0(deadband[16]), .I1(n455[16]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n68314));
    defparam i48819_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i49554_3_lut (.I0(n69873), .I1(n455[12]), .I2(n25_adj_4936), 
            .I3(GND_net), .O(n69049));   // verilog/motorControl.v(63[16:31])
    defparam i49554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4956));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i50375_3_lut (.I0(n4_adj_4956), .I1(n455[13]), .I2(n27_adj_4942), 
            .I3(GND_net), .O(n69870));   // verilog/motorControl.v(63[16:31])
    defparam i50375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50792_3_lut (.I0(n70286), .I1(n233[11]), .I2(n23_adj_4609), 
            .I3(GND_net), .O(n70287));   // verilog/motorControl.v(56[14:36])
    defparam i50792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50376_3_lut (.I0(n69870), .I1(n455[14]), .I2(n29_adj_4930), 
            .I3(GND_net), .O(n69871));   // verilog/motorControl.v(63[16:31])
    defparam i50376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48551_4_lut (.I0(n33_adj_4938), .I1(n31_adj_4931), .I2(n29_adj_4930), 
            .I3(n68088), .O(n68046));
    defparam i48551_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_3_lut_4_lut_adj_956 (.I0(\Ki[2] ), .I1(n335[18]), .I2(n52562), 
            .I3(n23323[0]), .O(n23266[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_956.LUT_INIT = 16'h8778;
    SB_LUT4 i51353_4_lut (.I0(n30_adj_4951), .I1(n10_adj_4950), .I2(n35_adj_4937), 
            .I3(n68040), .O(n70848));   // verilog/motorControl.v(63[16:31])
    defparam i51353_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49556_3_lut (.I0(n69871), .I1(n455[15]), .I2(n31_adj_4931), 
            .I3(GND_net), .O(n69051));   // verilog/motorControl.v(63[16:31])
    defparam i49556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51408_4_lut (.I0(n69051), .I1(n70848), .I2(n35_adj_4937), 
            .I3(n68046), .O(n70903));   // verilog/motorControl.v(63[16:31])
    defparam i51408_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51409_3_lut (.I0(n70903), .I1(n455[18]), .I2(n37_adj_4933), 
            .I3(GND_net), .O(n70904));   // verilog/motorControl.v(63[16:31])
    defparam i51409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34531_3_lut_4_lut (.I0(\Ki[2] ), .I1(n335[18]), .I2(n52562), 
            .I3(n23323[0]), .O(n4_adj_4943));   // verilog/motorControl.v(61[29:40])
    defparam i34531_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i48653_2_lut_4_lut (.I0(n455[21]), .I1(n34[21]), .I2(n455[9]), 
            .I3(n34[9]), .O(n68148));
    defparam i48653_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51391_3_lut (.I0(n70904), .I1(n455[19]), .I2(n39_adj_4928), 
            .I3(GND_net), .O(n70886));   // verilog/motorControl.v(63[16:31])
    defparam i51391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48522_4_lut (.I0(n43_adj_4932), .I1(n41_adj_4927), .I2(n39_adj_4928), 
            .I3(n70702), .O(n68017));
    defparam i48522_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50961_4_lut (.I0(n69049), .I1(n69804), .I2(n45_adj_4929), 
            .I3(n68013), .O(n70456));   // verilog/motorControl.v(63[16:31])
    defparam i50961_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51371_3_lut (.I0(n70886), .I1(n455[20]), .I2(n41_adj_4927), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(63[16:31])
    defparam i51371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50963_4_lut (.I0(n40), .I1(n70456), .I2(n45_adj_4929), .I3(n68017), 
            .O(n70458));   // verilog/motorControl.v(63[16:31])
    defparam i50963_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34518_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n23266[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34518_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i48725_2_lut_4_lut (.I0(n455[16]), .I1(n34[16]), .I2(n455[7]), 
            .I3(n34[7]), .O(n68220));
    defparam i48725_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i41_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4957));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4958));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i45_2_lut (.I0(PWMLimit[22]), .I1(setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4959));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4960));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34520_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n52562));   // verilog/motorControl.v(61[29:40])
    defparam i34520_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_9_i31_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4961));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4962));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i25_2_lut (.I0(PWMLimit[12]), .I1(setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4963));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i37_2_lut (.I0(PWMLimit[18]), .I1(setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4964));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i35_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4965));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i11_2_lut (.I0(PWMLimit[5]), .I1(setpoint[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4966));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4602));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i13_2_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4967));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i15_2_lut (.I0(PWMLimit[7]), .I1(setpoint[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4968));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17), 
            .I3(GND_net), .O(n8_adj_4969));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4599));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4970));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i33_2_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4971));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(\control_mode[0] ), .I1(\control_mode[7] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4972));
    defparam i2_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut (.I0(\control_mode[6] ), .I1(n62692), .I2(n10_adj_4972), 
            .I3(\control_mode[1] ), .O(n59791));
    defparam i7_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 n9977_bdd_4_lut_51919 (.I0(n9977), .I1(n67723), .I2(setpoint[9]), 
            .I3(n4749), .O(n71457));
    defparam n9977_bdd_4_lut_51919.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4914), .I1(n233[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4973));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i9_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4974));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48949_4_lut (.I0(n43_c), .I1(n25), .I2(n23_adj_4609), .I3(n68510), 
            .O(n68444));
    defparam i48949_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n71457_bdd_4_lut (.I0(n71457), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4749), .O(n71460));
    defparam n71457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50301_4_lut (.I0(n24_adj_4973), .I1(n8_adj_4969), .I2(n45), 
            .I3(n68441), .O(n69796));   // verilog/motorControl.v(56[14:36])
    defparam i50301_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 LessThan_9_i17_2_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4975));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49514_3_lut (.I0(n70287), .I1(n233[12]), .I2(n25), .I3(GND_net), 
            .O(n69009));   // verilog/motorControl.v(56[14:36])
    defparam i49514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i19_2_lut (.I0(PWMLimit[9]), .I1(setpoint[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4976));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4977));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i21_2_lut (.I0(PWMLimit[10]), .I1(setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4978));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n335[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i75_2_lut (.I0(\Ki[1] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4596));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4595));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49217_4_lut (.I0(n21_adj_4978), .I1(n19_adj_4976), .I2(n17_adj_4975), 
            .I3(n9_adj_4974), .O(n68712));
    defparam i49217_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50789_3_lut (.I0(n4_adj_4977), .I1(n233[13]), .I2(n27), .I3(GND_net), 
            .O(n70284));   // verilog/motorControl.v(56[14:36])
    defparam i50789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49192_4_lut (.I0(n27_adj_4970), .I1(n15_adj_4968), .I2(n13_adj_4967), 
            .I3(n11_adj_4966), .O(n68687));
    defparam i49192_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i30_3_lut (.I0(n12_adj_4918), .I1(setpoint[17]), 
            .I2(n35_adj_4965), .I3(GND_net), .O(n30_adj_4980));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4592));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50790_3_lut (.I0(n70284), .I1(n233[14]), .I2(n29_adj_4636), 
            .I3(GND_net), .O(n70285));   // verilog/motorControl.v(56[14:36])
    defparam i50790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4590));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50205_4_lut (.I0(n13_adj_4967), .I1(n11_adj_4966), .I2(n9_adj_4974), 
            .I3(n68829), .O(n69700));
    defparam i50205_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4589));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4587));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9977_bdd_4_lut_51914 (.I0(n9977), .I1(n67722), .I2(setpoint[8]), 
            .I3(n4749), .O(n71451));
    defparam n9977_bdd_4_lut_51914.LUT_INIT = 16'he4aa;
    SB_LUT4 i50169_4_lut (.I0(n19_adj_4976), .I1(n17_adj_4975), .I2(n15_adj_4968), 
            .I3(n69700), .O(n69664));
    defparam i50169_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48980_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4636), .I3(n68489), 
            .O(n68475));
    defparam i48980_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51167_4_lut (.I0(n25_adj_4963), .I1(n23_adj_4962), .I2(n21_adj_4978), 
            .I3(n69664), .O(n70662));
    defparam i51167_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51117_4_lut (.I0(n30), .I1(n10_adj_4819), .I2(n35_adj_4800), 
            .I3(n68467), .O(n70612));   // verilog/motorControl.v(56[14:36])
    defparam i51117_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49516_3_lut (.I0(n70285), .I1(n233[15]), .I2(n31), .I3(GND_net), 
            .O(n69011));   // verilog/motorControl.v(56[14:36])
    defparam i49516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51325_4_lut (.I0(n69011), .I1(n70612), .I2(n35_adj_4800), 
            .I3(n68475), .O(n70820));   // verilog/motorControl.v(56[14:36])
    defparam i51325_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51326_3_lut (.I0(n70820), .I1(n233[18]), .I2(n37), .I3(GND_net), 
            .O(n70821));   // verilog/motorControl.v(56[14:36])
    defparam i51326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51308_3_lut (.I0(n70821), .I1(n233[19]), .I2(n39), .I3(GND_net), 
            .O(n70803));   // verilog/motorControl.v(56[14:36])
    defparam i51308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50579_4_lut (.I0(n31_adj_4961), .I1(n29_adj_4960), .I2(n27_adj_4970), 
            .I3(n70662), .O(n70074));
    defparam i50579_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4584));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51254_4_lut (.I0(n37_adj_4964), .I1(n35_adj_4965), .I2(n33_adj_4971), 
            .I3(n70074), .O(n70749));
    defparam i51254_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4583));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4582));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4581));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50807_3_lut (.I0(n6_adj_4981), .I1(setpoint[10]), .I2(n21_adj_4978), 
            .I3(GND_net), .O(n70302));   // verilog/motorControl.v(45[16:33])
    defparam i50807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50808_3_lut (.I0(n70302), .I1(setpoint[11]), .I2(n23_adj_4962), 
            .I3(GND_net), .O(n70303));   // verilog/motorControl.v(45[16:33])
    defparam i50808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i24_3_lut (.I0(n16_adj_4916), .I1(setpoint[22]), 
            .I2(n45_adj_4959), .I3(GND_net), .O(n24_adj_4982));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49125_4_lut (.I0(n43), .I1(n25_adj_4963), .I2(n23_adj_4962), 
            .I3(n68712), .O(n68620));
    defparam i49125_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50297_4_lut (.I0(n24_adj_4982), .I1(n8_adj_4909), .I2(n45_adj_4959), 
            .I3(n68610), .O(n69792));   // verilog/motorControl.v(45[16:33])
    defparam i50297_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49494_3_lut (.I0(n70303), .I1(setpoint[12]), .I2(n25_adj_4963), 
            .I3(GND_net), .O(n68989));   // verilog/motorControl.v(45[16:33])
    defparam i49494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48953_4_lut (.I0(n43_c), .I1(n41_adj_4600), .I2(n39), .I3(n70729), 
            .O(n68448));
    defparam i48953_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_4984));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50803_3_lut (.I0(n4_adj_4984), .I1(setpoint[13]), .I2(n27_adj_4970), 
            .I3(GND_net), .O(n70298));   // verilog/motorControl.v(45[16:33])
    defparam i50803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50804_3_lut (.I0(n70298), .I1(setpoint[14]), .I2(n29_adj_4960), 
            .I3(GND_net), .O(n70299));   // verilog/motorControl.v(45[16:33])
    defparam i50804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49181_4_lut (.I0(n33_adj_4971), .I1(n31_adj_4961), .I2(n29_adj_4960), 
            .I3(n68687), .O(n68676));
    defparam i49181_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4580));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4579));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50953_4_lut (.I0(n69009), .I1(n69796), .I2(n45), .I3(n68444), 
            .O(n70448));   // verilog/motorControl.v(56[14:36])
    defparam i50953_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4577));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4576));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49522_3_lut (.I0(n70803), .I1(n233[20]), .I2(n41_adj_4600), 
            .I3(GND_net), .O(n69017));   // verilog/motorControl.v(56[14:36])
    defparam i49522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51113_4_lut (.I0(n30_adj_4980), .I1(n10_adj_4917), .I2(n35_adj_4965), 
            .I3(n68663), .O(n70608));   // verilog/motorControl.v(45[16:33])
    defparam i51113_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4575));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49496_3_lut (.I0(n70299), .I1(setpoint[15]), .I2(n31_adj_4961), 
            .I3(GND_net), .O(n68991));   // verilog/motorControl.v(45[16:33])
    defparam i49496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51321_4_lut (.I0(n68991), .I1(n70608), .I2(n35_adj_4965), 
            .I3(n68676), .O(n70816));   // verilog/motorControl.v(45[16:33])
    defparam i51321_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51322_3_lut (.I0(n70816), .I1(setpoint[18]), .I2(n37_adj_4964), 
            .I3(GND_net), .O(n70817));   // verilog/motorControl.v(45[16:33])
    defparam i51322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51312_3_lut (.I0(n70817), .I1(setpoint[19]), .I2(n39_adj_4958), 
            .I3(GND_net), .O(n70807));   // verilog/motorControl.v(45[16:33])
    defparam i51312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51195_4_lut (.I0(n69017), .I1(n70448), .I2(n45), .I3(n68448), 
            .O(n70690));   // verilog/motorControl.v(56[14:36])
    defparam i51195_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49129_4_lut (.I0(n43), .I1(n41_adj_4957), .I2(n39_adj_4958), 
            .I3(n70749), .O(n68624));
    defparam i49129_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50949_4_lut (.I0(n68989), .I1(n69792), .I2(n45_adj_4959), 
            .I3(n68620), .O(n70444));   // verilog/motorControl.v(45[16:33])
    defparam i50949_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51196_3_lut (.I0(n70690), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i51196_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49502_3_lut (.I0(n70807), .I1(setpoint[20]), .I2(n41_adj_4957), 
            .I3(GND_net), .O(n68997));   // verilog/motorControl.v(45[16:33])
    defparam i49502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51191_4_lut (.I0(n68997), .I1(n70444), .I2(n45_adj_4959), 
            .I3(n68624), .O(n70686));   // verilog/motorControl.v(45[16:33])
    defparam i51191_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51192_3_lut (.I0(n70686), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i51192_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49035_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n68530));
    defparam i49035_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i49056_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n68551));
    defparam i49056_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i3_4_lut (.I0(n7067), .I1(n7069), .I2(n27766), .I3(n62775), 
            .O(n4749));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i48473_4_lut (.I0(n27_adj_4865), .I1(n15_adj_4866), .I2(n13_adj_4864), 
            .I3(n11_adj_4863), .O(n67968));
    defparam i48473_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4867), 
            .I3(GND_net), .O(n12_adj_4985));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4864), 
            .I3(GND_net), .O(n10_adj_4986));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_4985), .I1(n535[17]), .I2(n35_adj_4858), 
            .I3(GND_net), .O(n30_adj_4987));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4574));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49477_4_lut (.I0(n13_adj_4864), .I1(n11_adj_4863), .I2(n9_adj_4857), 
            .I3(n68003), .O(n68972));
    defparam i49477_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_update), .I1(n59791), .I2(n105), 
            .I3(GND_net), .O(n7069));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i49471_4_lut (.I0(n19_adj_4856), .I1(n17_adj_4855), .I2(n15_adj_4866), 
            .I3(n68972), .O(n68966));
    defparam i49471_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50943_4_lut (.I0(n25_adj_4854), .I1(n23_adj_4853), .I2(n21_adj_4852), 
            .I3(n68966), .O(n70438));
    defparam i50943_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(control_update), .I1(n59791), .I2(n131_adj_4847), 
            .I3(n105), .O(n7067));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_957 (.I0(control_update), .I1(n59791), 
            .I2(n131_adj_4847), .I3(n105), .O(n27800));
    defparam i1_2_lut_3_lut_4_lut_adj_957.LUT_INIT = 16'h0080;
    SB_LUT4 i1_3_lut_4_lut_adj_958 (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4988), 
            .I3(n23360[1]), .O(n23323[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_958.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), 
            .I2(setpoint[2]), .I3(GND_net), .O(n6_adj_4981));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50271_4_lut (.I0(n31_adj_4861), .I1(n29_adj_4860), .I2(n27_adj_4865), 
            .I3(n70438), .O(n69766));
    defparam i50271_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49334_3_lut_4_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(setpoint[2]), 
            .I3(PWMLimit[2]), .O(n68829));   // verilog/motorControl.v(45[16:33])
    defparam i49334_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51187_4_lut (.I0(n37_adj_4851), .I1(n35_adj_4858), .I2(n33_adj_4867), 
            .I3(n69766), .O(n70682));
    defparam i51187_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34464_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4988), 
            .I3(n23360[1]), .O(n6_adj_4552));   // verilog/motorControl.v(61[29:40])
    defparam i34464_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i50915_3_lut (.I0(n6_adj_4989), .I1(n535[10]), .I2(n21_adj_4852), 
            .I3(GND_net), .O(n70410));   // verilog/motorControl.v(65[25:41])
    defparam i50915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50916_3_lut (.I0(n70410), .I1(n535[11]), .I2(n23_adj_4853), 
            .I3(GND_net), .O(n70411));   // verilog/motorControl.v(65[25:41])
    defparam i50916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4859), 
            .I3(GND_net), .O(n16_adj_4990));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n70458), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n27764), .O(n27766));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff71;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4855), 
            .I3(GND_net), .O(n8_adj_4991));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_4990), .I1(n535[22]), .I2(n45_adj_4850), 
            .I3(GND_net), .O(n24_adj_4992));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_959 (.I0(n70458), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n27764), .O(n4_adj_4993));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_959.LUT_INIT = 16'hff8e;
    SB_LUT4 i48491_4_lut (.I0(n21_adj_4852), .I1(n19_adj_4856), .I2(n17_adj_4855), 
            .I3(n9_adj_4857), .O(n67986));
    defparam i48491_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48393_4_lut (.I0(n43_adj_4859), .I1(n25_adj_4854), .I2(n23_adj_4853), 
            .I3(n67986), .O(n67888));
    defparam i48393_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50311_4_lut (.I0(n24_adj_4992), .I1(n8_adj_4991), .I2(n45_adj_4850), 
            .I3(n67878), .O(n69806));   // verilog/motorControl.v(65[25:41])
    defparam i50311_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50645_3_lut (.I0(n70411), .I1(n535[12]), .I2(n25_adj_4854), 
            .I3(GND_net), .O(n70140));   // verilog/motorControl.v(65[25:41])
    defparam i50645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_4994));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50881_3_lut (.I0(n4_adj_4994), .I1(n535[13]), .I2(n27_adj_4865), 
            .I3(GND_net), .O(n70376));   // verilog/motorControl.v(65[25:41])
    defparam i50881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48972_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n68467));
    defparam i48972_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50882_3_lut (.I0(n70376), .I1(n535[14]), .I2(n29_adj_4860), 
            .I3(GND_net), .O(n70377));   // verilog/motorControl.v(65[25:41])
    defparam i50882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48453_4_lut (.I0(n33_adj_4867), .I1(n31_adj_4861), .I2(n29_adj_4860), 
            .I3(n67968), .O(n67948));
    defparam i48453_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51240_4_lut (.I0(n30_adj_4987), .I1(n10_adj_4986), .I2(n35_adj_4858), 
            .I3(n67942), .O(n70735));   // verilog/motorControl.v(65[25:41])
    defparam i51240_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50647_3_lut (.I0(n70377), .I1(n535[15]), .I2(n31_adj_4861), 
            .I3(GND_net), .O(n70142));   // verilog/motorControl.v(65[25:41])
    defparam i50647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51394_4_lut (.I0(n70142), .I1(n70735), .I2(n35_adj_4858), 
            .I3(n67948), .O(n70889));   // verilog/motorControl.v(65[25:41])
    defparam i51394_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4995));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51395_3_lut (.I0(n70889), .I1(n535[18]), .I2(n37_adj_4851), 
            .I3(GND_net), .O(n70890));   // verilog/motorControl.v(65[25:41])
    defparam i51395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51348_3_lut (.I0(n70890), .I1(n535[19]), .I2(n39_adj_4849), 
            .I3(GND_net), .O(n70843));   // verilog/motorControl.v(65[25:41])
    defparam i51348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48397_4_lut (.I0(n43_adj_4859), .I1(n41_adj_4848), .I2(n39_adj_4849), 
            .I3(n70682), .O(n67892));
    defparam i48397_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50650_4_lut (.I0(n70140), .I1(n69806), .I2(n45_adj_4850), 
            .I3(n67888), .O(n70145));   // verilog/motorControl.v(65[25:41])
    defparam i50650_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51271_3_lut (.I0(n70843), .I1(n535[20]), .I2(n41_adj_4848), 
            .I3(GND_net), .O(n40_adj_4996));   // verilog/motorControl.v(65[25:41])
    defparam i51271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50967_4_lut (.I0(n40_adj_4996), .I1(n70145), .I2(n45_adj_4850), 
            .I3(n67892), .O(n70462));   // verilog/motorControl.v(65[25:41])
    defparam i50967_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_4_lut (.I0(n70462), .I1(n4_adj_4993), .I2(n455[23]), .I3(n535[23]), 
            .O(n62767));
    defparam i2_4_lut.LUT_INIT = 16'hdfcd;
    SB_LUT4 i4428_4_lut (.I0(n7067), .I1(n4749), .I2(n62767), .I3(n27800), 
            .O(n9977));
    defparam i4428_4_lut.LUT_INIT = 16'hbbab;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4446));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4445));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34456_3_lut_4_lut (.I0(n62_adj_4506), .I1(n131), .I2(n204), 
            .I3(n23360[0]), .O(n4_adj_4988));   // verilog/motorControl.v(61[29:40])
    defparam i34456_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4997));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48651_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(PWMLimit[2]), .O(n68146));   // verilog/motorControl.v(63[16:31])
    defparam i48651_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4444));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4953));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_3_lut_4_lut_adj_960 (.I0(n62_adj_4506), .I1(n131), .I2(n204), 
            .I3(n23360[0]), .O(n23323[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_960.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_961 (.I0(n59791), .I1(control_update), .I2(n506), 
            .I3(n480), .O(n27764));
    defparam i1_3_lut_4_lut_adj_961.LUT_INIT = 16'hbbbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(n59791), .I1(control_update), .I2(n506), 
            .I3(n480), .O(n62775));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4443));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4998));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4442));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4441));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n310[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i13_3_lut (.I0(n310[12]), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n335[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4573));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i26_2_lut (.I0(\Ki[0] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4572));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4571));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4569));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4567));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4999));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4566));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4565));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4564));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5000));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4562));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4561));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5001));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4559));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71451_bdd_4_lut (.I0(n71451), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4749), .O(n71454));
    defparam n71451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5002));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5003));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5004));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5005));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5006));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5007));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9977_bdd_4_lut_51909 (.I0(n9977), .I1(n67721), .I2(setpoint[7]), 
            .I3(n4749), .O(n71445));
    defparam n9977_bdd_4_lut_51909.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5008));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(n233[18]), .I1(n285[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5009));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34427_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n54083));   // verilog/motorControl.v(61[20:26])
    defparam i34427_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i34421_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n52453));   // verilog/motorControl.v(61[20:26])
    defparam i34421_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(n233[10]), .I1(n285[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5010));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48912_4_lut (.I0(n21_adj_5010), .I1(n19_adj_5004), .I2(n17_adj_5002), 
            .I3(n9_adj_4815), .O(n68407));
    defparam i48912_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4440));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48782_3_lut_4_lut (.I0(n455[3]), .I1(n34[3]), .I2(n34[2]), 
            .I3(n455[2]), .O(n68277));   // verilog/motorControl.v(62[35:55])
    defparam i48782_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_28_i6_3_lut_3_lut (.I0(n455[3]), .I1(n34[3]), .I2(n34[2]), 
            .I3(GND_net), .O(n6_adj_4911));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48870_3_lut_4_lut (.I0(deadband[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(deadband[2]), .O(n68365));   // verilog/motorControl.v(62[14:31])
    defparam i48870_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4923));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i48900_4_lut (.I0(n27_adj_5000), .I1(n15_adj_4818), .I2(n13_adj_4817), 
            .I3(n11_adj_4816), .O(n68395));
    defparam i48900_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_5007), 
            .I3(GND_net), .O(n12_adj_5011));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48585_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[4]), 
            .I3(GND_net), .O(n67718));
    defparam i48585_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48584_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n67719));
    defparam i48584_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4439));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4817), 
            .I3(GND_net), .O(n10_adj_5012));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_5011), .I1(n285[17]), .I2(n35_adj_5008), 
            .I3(GND_net), .O(n30_adj_5013));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48583_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n67720));
    defparam i48583_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48582_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n67721));
    defparam i48582_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48581_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n67722));
    defparam i48581_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48580_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n67723));
    defparam i48580_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48579_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n67724));
    defparam i48579_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48578_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n67725));
    defparam i48578_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48577_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n67726));
    defparam i48577_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48576_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n67727));
    defparam i48576_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48575_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n67728));
    defparam i48575_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48574_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[15]), 
            .I3(GND_net), .O(n67729));
    defparam i48574_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48573_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n67730));
    defparam i48573_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48586_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n67717));
    defparam i48586_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48399_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n67715));
    defparam i48399_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i49937_4_lut (.I0(n13_adj_4817), .I1(n11_adj_4816), .I2(n9_adj_4815), 
            .I3(n68435), .O(n69432));
    defparam i49937_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4438));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48587_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n67716));
    defparam i48587_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49929_4_lut (.I0(n19_adj_5004), .I1(n17_adj_5002), .I2(n15_adj_4818), 
            .I3(n69432), .O(n69424));
    defparam i49929_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48431_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n67737));
    defparam i48431_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48564_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n67735));
    defparam i48564_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48565_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[20]), 
            .I3(GND_net), .O(n67734));
    defparam i48565_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48566_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n67733));
    defparam i48566_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48572_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n67731));
    defparam i48572_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4437));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48567_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n67732));
    defparam i48567_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4436));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4435));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48403_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[23]), 
            .I3(GND_net), .O(n67775));
    defparam i48403_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48328_2_lut_3_lut (.I0(n7069), .I1(n27766), .I2(PWMLimit[0]), 
            .I3(GND_net), .O(n67714));
    defparam i48328_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i51085_4_lut (.I0(n25_adj_5001), .I1(n23_adj_5006), .I2(n21_adj_5010), 
            .I3(n69424), .O(n70580));
    defparam i51085_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50469_4_lut (.I0(n31_adj_4999), .I1(n29_adj_4998), .I2(n27_adj_5000), 
            .I3(n70580), .O(n69964));
    defparam i50469_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51230_4_lut (.I0(n37_adj_5009), .I1(n35_adj_5008), .I2(n33_adj_5007), 
            .I3(n69964), .O(n70725));
    defparam i51230_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48508_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n68003));   // verilog/motorControl.v(65[25:41])
    defparam i48508_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4989));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_5005), 
            .I3(GND_net), .O(n16_adj_5014));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34443_2_lut_4_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(\Ki[1] ), 
            .I3(n335[19]), .O(n23323[0]));   // verilog/motorControl.v(61[29:40])
    defparam i34443_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i50785_3_lut (.I0(n6_adj_4934), .I1(n285[10]), .I2(n21_adj_5010), 
            .I3(GND_net), .O(n70280));   // verilog/motorControl.v(58[23:46])
    defparam i50785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50786_3_lut (.I0(n70280), .I1(n285[11]), .I2(n23_adj_5006), 
            .I3(GND_net), .O(n70281));   // verilog/motorControl.v(58[23:46])
    defparam i50786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_5002), 
            .I3(GND_net), .O(n8_adj_5015));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_5014), .I1(n285[22]), .I2(n45_adj_5003), 
            .I3(GND_net), .O(n24_adj_5016));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48878_4_lut (.I0(n43_adj_5005), .I1(n25_adj_5001), .I2(n23_adj_5006), 
            .I3(n68407), .O(n68373));
    defparam i48878_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50303_4_lut (.I0(n24_adj_5016), .I1(n8_adj_5015), .I2(n45_adj_5003), 
            .I3(n68369), .O(n69798));   // verilog/motorControl.v(58[23:46])
    defparam i50303_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49524_3_lut (.I0(n70281), .I1(n285[12]), .I2(n25_adj_5001), 
            .I3(GND_net), .O(n69019));   // verilog/motorControl.v(58[23:46])
    defparam i49524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_5017));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i50783_3_lut (.I0(n4_adj_5017), .I1(n285[13]), .I2(n27_adj_5000), 
            .I3(GND_net), .O(n70278));   // verilog/motorControl.v(58[23:46])
    defparam i50783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49113_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n68608));   // verilog/motorControl.v(47[25:43])
    defparam i49113_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_4843));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50784_3_lut (.I0(n70278), .I1(n285[14]), .I2(n29_adj_4998), 
            .I3(GND_net), .O(n70279));   // verilog/motorControl.v(58[23:46])
    defparam i50784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48896_4_lut (.I0(n33_adj_5007), .I1(n31_adj_4999), .I2(n29_adj_4998), 
            .I3(n68395), .O(n68391));
    defparam i48896_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n71445_bdd_4_lut (.I0(n71445), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4749), .O(n71448));
    defparam n71445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51119_4_lut (.I0(n30_adj_5013), .I1(n10_adj_5012), .I2(n35_adj_5008), 
            .I3(n68387), .O(n70614));   // verilog/motorControl.v(58[23:46])
    defparam i51119_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 n9977_bdd_4_lut_51904 (.I0(n9977), .I1(n67720), .I2(setpoint[6]), 
            .I3(n4749), .O(n71439));
    defparam n9977_bdd_4_lut_51904.LUT_INIT = 16'he4aa;
    SB_LUT4 i49526_3_lut (.I0(n70279), .I1(n285[15]), .I2(n31_adj_4999), 
            .I3(GND_net), .O(n69021));   // verilog/motorControl.v(58[23:46])
    defparam i49526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51329_4_lut (.I0(n69021), .I1(n70614), .I2(n35_adj_5008), 
            .I3(n68391), .O(n70824));   // verilog/motorControl.v(58[23:46])
    defparam i51329_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51330_3_lut (.I0(n70824), .I1(n285[18]), .I2(n37_adj_5009), 
            .I3(GND_net), .O(n70825));   // verilog/motorControl.v(58[23:46])
    defparam i51330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51304_3_lut (.I0(n70825), .I1(n285[19]), .I2(n39_adj_4997), 
            .I3(GND_net), .O(n70799));   // verilog/motorControl.v(58[23:46])
    defparam i51304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4434));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4433));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4432));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4431));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4430));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71439_bdd_4_lut (.I0(n71439), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4749), .O(n71442));
    defparam n71439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48882_4_lut (.I0(n43_adj_5005), .I1(n41_adj_4995), .I2(n39_adj_4997), 
            .I3(n70725), .O(n68377));
    defparam i48882_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50955_4_lut (.I0(n69019), .I1(n69798), .I2(n45_adj_5003), 
            .I3(n68373), .O(n70450));   // verilog/motorControl.v(58[23:46])
    defparam i50955_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49532_3_lut (.I0(n70799), .I1(n285[20]), .I2(n41_adj_4995), 
            .I3(GND_net), .O(n69027));   // verilog/motorControl.v(58[23:46])
    defparam i49532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51197_4_lut (.I0(n69027), .I1(n70450), .I2(n45_adj_5003), 
            .I3(n68377), .O(n70692));   // verilog/motorControl.v(58[23:46])
    defparam i51197_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51198_3_lut (.I0(n70692), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i51198_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n335[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9977_bdd_4_lut_51899 (.I0(n9977), .I1(n67719), .I2(setpoint[5]), 
            .I3(n4749), .O(n71433));
    defparam n9977_bdd_4_lut_51899.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71433_bdd_4_lut (.I0(n71433), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4749), .O(n71436));
    defparam n71433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9977_bdd_4_lut_51894 (.I0(n9977), .I1(n67718), .I2(setpoint[4]), 
            .I3(n4749), .O(n71427));
    defparam n9977_bdd_4_lut_51894.LUT_INIT = 16'he4aa;
    SB_LUT4 n71427_bdd_4_lut (.I0(n71427), .I1(n535[4]), .I2(n455[4]), 
            .I3(n4749), .O(n71430));
    defparam n71427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i34605_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4654), 
            .I3(GND_net), .O(n23287[0]));   // verilog/motorControl.v(61[20:26])
    defparam i34605_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_3_lut_4_lut_adj_962 (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4654), 
            .I3(n64059), .O(n23287[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut_adj_962.LUT_INIT = 16'h7f80;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4513));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    
endmodule
